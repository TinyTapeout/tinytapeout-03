VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO dwisehart_top
  CLASS BLOCK ;
  FOREIGN dwisehart_top ;
  ORIGIN 0.000 0.000 ;
  SIZE 150.000 BY 170.000 ;
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 8.200 2.000 8.800 ;
    END
  END io_in[0]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 18.400 2.000 19.000 ;
    END
  END io_in[1]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 28.600 2.000 29.200 ;
    END
  END io_in[2]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 38.800 2.000 39.400 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 49.000 2.000 49.600 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 59.200 2.000 59.800 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 69.400 2.000 70.000 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 79.600 2.000 80.200 ;
    END
  END io_in[7]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 89.800 2.000 90.400 ;
    END
  END io_out[0]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 100.000 2.000 100.600 ;
    END
  END io_out[1]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 110.200 2.000 110.800 ;
    END
  END io_out[2]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 120.400 2.000 121.000 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 130.600 2.000 131.200 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 140.800 2.000 141.400 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 151.000 2.000 151.600 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 161.200 2.000 161.800 ;
    END
  END io_out[7]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 22.085 5.200 23.685 163.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 56.815 5.200 58.415 163.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 91.545 5.200 93.145 163.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 126.275 5.200 127.875 163.440 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 39.450 5.200 41.050 163.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 74.180 5.200 75.780 163.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 108.910 5.200 110.510 163.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 143.640 5.200 145.240 163.440 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 5.355 144.440 163.285 ;
      LAYER met1 ;
        RECT 1.450 2.420 145.240 163.440 ;
      LAYER met2 ;
        RECT 1.010 2.195 145.210 163.385 ;
      LAYER met3 ;
        RECT 0.985 162.200 145.230 163.365 ;
        RECT 2.400 160.800 145.230 162.200 ;
        RECT 0.985 152.000 145.230 160.800 ;
        RECT 2.400 150.600 145.230 152.000 ;
        RECT 0.985 141.800 145.230 150.600 ;
        RECT 2.400 140.400 145.230 141.800 ;
        RECT 0.985 131.600 145.230 140.400 ;
        RECT 2.400 130.200 145.230 131.600 ;
        RECT 0.985 121.400 145.230 130.200 ;
        RECT 2.400 120.000 145.230 121.400 ;
        RECT 0.985 111.200 145.230 120.000 ;
        RECT 2.400 109.800 145.230 111.200 ;
        RECT 0.985 101.000 145.230 109.800 ;
        RECT 2.400 99.600 145.230 101.000 ;
        RECT 0.985 90.800 145.230 99.600 ;
        RECT 2.400 89.400 145.230 90.800 ;
        RECT 0.985 80.600 145.230 89.400 ;
        RECT 2.400 79.200 145.230 80.600 ;
        RECT 0.985 70.400 145.230 79.200 ;
        RECT 2.400 69.000 145.230 70.400 ;
        RECT 0.985 60.200 145.230 69.000 ;
        RECT 2.400 58.800 145.230 60.200 ;
        RECT 0.985 50.000 145.230 58.800 ;
        RECT 2.400 48.600 145.230 50.000 ;
        RECT 0.985 39.800 145.230 48.600 ;
        RECT 2.400 38.400 145.230 39.800 ;
        RECT 0.985 29.600 145.230 38.400 ;
        RECT 2.400 28.200 145.230 29.600 ;
        RECT 0.985 19.400 145.230 28.200 ;
        RECT 2.400 18.000 145.230 19.400 ;
        RECT 0.985 9.200 145.230 18.000 ;
        RECT 2.400 7.800 145.230 9.200 ;
        RECT 0.985 2.215 145.230 7.800 ;
      LAYER met4 ;
        RECT 3.055 4.800 21.685 161.665 ;
        RECT 24.085 4.800 39.050 161.665 ;
        RECT 41.450 4.800 56.415 161.665 ;
        RECT 58.815 4.800 73.780 161.665 ;
        RECT 76.180 4.800 91.145 161.665 ;
        RECT 93.545 4.800 108.510 161.665 ;
        RECT 110.910 4.800 124.825 161.665 ;
        RECT 3.055 2.215 124.825 4.800 ;
  END
END dwisehart_top
END LIBRARY

