/* Automatically generated from https://wokwi.com/projects/361684719151591425 */

`default_nettype none

module user_module_361684719151591425(
  input [7:0] io_in,
  output [7:0] io_out
);
  wire net1 = io_in[0];
  wire net2 = io_in[1];
  wire net3 = io_in[2];
  wire net4 = io_in[3];
  wire net5 = io_in[6];
  wire net6 = io_in[7];
  wire net7;
  wire net8;
  wire net9;
  wire net10;
  wire net11;
  wire net12;
  wire net13;
  wire net14;
  wire net15 = 1'b0;
  wire net16 = 1'b1;
  wire net17;
  wire net18;
  wire net19;
  wire net20;
  wire net21;
  wire net22;
  wire net23;
  wire net24;
  wire net25;
  wire net26;
  wire net27;
  wire net28;
  wire net29;
  wire net30;
  wire net31;
  wire net32;
  wire net33;
  wire net34;
  wire net35;
  wire net36;
  wire net37;
  wire net38;
  wire net39;
  wire net40;
  wire net41;
  wire net42;
  wire net43;
  wire net44;
  wire net45;
  wire net46;
  wire net47;
  wire net48;
  wire net49;
  wire net50;
  wire net51;
  wire net52;
  wire net53;
  wire net54;
  wire net55;
  wire net56;
  wire net57;
  wire net58;
  wire net59;
  wire net60;
  wire net61;
  wire net62;
  wire net63;
  wire net64;
  wire net65;
  wire net66;
  wire net67;
  wire net68;
  wire net69;
  wire net70;
  wire net71;
  wire net72;
  wire net73;
  wire net74;
  wire net75;
  wire net76;
  wire net77;
  wire net78;
  wire net79;
  wire net80;
  wire net81;
  wire net82;
  wire net83;
  wire net84;
  wire net85;
  wire net86;
  wire net87;
  wire net88;
  wire net89;
  wire net90;
  wire net91;
  wire net92;
  wire net93;
  wire net94;
  wire net95;
  wire net96;
  wire net97;
  wire net98;
  wire net99;
  wire net100;
  wire net101;
  wire net102;
  wire net103;
  wire net104;
  wire net105;
  wire net106;
  wire net107;
  wire net108;
  wire net109;
  wire net110;
  wire net111;
  wire net112;
  wire net113;
  wire net114;
  wire net115;
  wire net116;
  wire net117;
  wire net118;
  wire net119;
  wire net120;
  wire net121;
  wire net122;
  wire net123;
  wire net124;
  wire net125;
  wire net126;
  wire net127;
  wire net128;
  wire net129;
  wire net130;
  wire net131;
  wire net132;
  wire net133;
  wire net134;
  wire net135;
  wire net136;
  wire net137;
  wire net138;
  wire net139;
  wire net140;
  wire net141;
  wire net142;
  wire net143;
  wire net144;
  wire net145;
  wire net146;
  wire net147;
  wire net148;
  wire net149;
  wire net150;
  wire net151;
  wire net152;
  wire net153;
  wire net154;
  wire net155;
  wire net156;
  wire net157;
  wire net158;
  wire net159;
  wire net160;
  wire net161;
  wire net162;
  wire net163;
  wire net164;
  wire net165;
  wire net166;
  wire net167;
  wire net168;
  wire net169;
  wire net170;
  wire net171;
  wire net172;
  wire net173;
  wire net174;
  wire net175;
  wire net176;
  wire net177;
  wire net178;
  wire net179;
  wire net180;
  wire net181;
  wire net182;
  wire net183;
  wire net184;
  wire net185;
  wire net186;
  wire net187;
  wire net188;
  wire net189;
  wire net190;
  wire net191;
  wire net192;
  wire net193;
  wire net194;
  wire net195;
  wire net196;
  wire net197;
  wire net198;
  wire net199;
  wire net200;
  wire net201;
  wire net202;
  wire net203;
  wire net204;
  wire net205;
  wire net206;
  wire net207;
  wire net208;
  wire net209;
  wire net210;
  wire net211;
  wire net212;
  wire net213;
  wire net214;
  wire net215;
  wire net216;
  wire net217;
  wire net218;
  wire net219;
  wire net220;
  wire net221;
  wire net222;
  wire net223;
  wire net224;
  wire net225;
  wire net226;
  wire net227;
  wire net228;
  wire net229;
  wire net230;
  wire net231;
  wire net232;
  wire net233;
  wire net234;
  wire net235;
  wire net236;
  wire net237;
  wire net238;
  wire net239;
  wire net240;
  wire net241;
  wire net242;
  wire net243;
  wire net244;
  wire net245;
  wire net246;
  wire net247;
  wire net248;
  wire net249;
  wire net250;
  wire net251;
  wire net252;
  wire net253;
  wire net254;
  wire net255;
  wire net256;
  wire net257;
  wire net258;
  wire net259;
  wire net260;
  wire net261;
  wire net262;
  wire net263;
  wire net264;
  wire net265;
  wire net266;
  wire net267;
  wire net268;
  wire net269;
  wire net270;
  wire net271;
  wire net272;
  wire net273;
  wire net274;
  wire net275;
  wire net276;
  wire net277;
  wire net278;
  wire net279;
  wire net280;
  wire net281;
  wire net282;
  wire net283;
  wire net284;

  assign io_out[0] = net7;
  assign io_out[1] = net8;
  assign io_out[2] = net9;
  assign io_out[3] = net10;
  assign io_out[4] = net11;
  assign io_out[5] = net12;
  assign io_out[6] = net13;
  assign io_out[7] = net14;

  not_cell not1 (
    .in (net1),
    .out (net17)
  );
  not_cell not2 (
    .in (net2),
    .out (net18)
  );
  not_cell not3 (
    .in (net3),
    .out (net19)
  );
  not_cell not4 (
    .in (net4),
    .out (net20)
  );
  not_cell not5 (
    .in (net5),
    .out (net21)
  );
  not_cell not6 (
    .in (net6),
    .out (net22)
  );
  and_cell and1 (
    .a (net22),
    .b (net5),
    .out (net23)
  );
  and_cell and2 (
    .a (net20),
    .b (net2),
    .out (net24)
  );
  and_cell and3 (
    .a (net23),
    .b (net24),
    .out (net25)
  );
  and_cell and4 (
    .a (net6),
    .b (net21),
    .out (net26)
  );
  and_cell and5 (
    .a (net19),
    .b (net17),
    .out (net27)
  );
  and_cell and6 (
    .a (net26),
    .b (net27),
    .out (net28)
  );
  or_cell or1 (
    .a (net25),
    .b (net28),
    .out (net29)
  );
  and_cell and7 (
    .a (net6),
    .b (net21),
    .out (net30)
  );
  and_cell and8 (
    .a (net20),
    .b (net2),
    .out (net31)
  );
  and_cell and9 (
    .a (net30),
    .b (net31),
    .out (net32)
  );
  and_cell and10 (
    .a (net6),
    .b (net21),
    .out (net33)
  );
  and_cell and11 (
    .a (net3),
    .b (net2),
    .out (net34)
  );
  and_cell and12 (
    .a (net33),
    .b (net34),
    .out (net35)
  );
  or_cell or2 (
    .a (net32),
    .b (net35),
    .out (net36)
  );
  and_cell and13 (
    .a (net6),
    .b (net21),
    .out (net37)
  );
  and_cell and14 (
    .a (net4),
    .b (net17),
    .out (net38)
  );
  and_cell and15 (
    .a (net37),
    .b (net38),
    .out (net39)
  );
  and_cell and16 (
    .a (net22),
    .b (net5),
    .out (net40)
  );
  and_cell and17 (
    .a (net20),
    .b (net19),
    .out (net41)
  );
  and_cell and18 (
    .a (net40),
    .b (net41),
    .out (net42)
  );
  and_cell and19 (
    .a (net42),
    .b (net17),
    .out (net43)
  );
  or_cell or3 (
    .a (net39),
    .b (net43),
    .out (net44)
  );
  or_cell or4 (
    .a (net29),
    .b (net36),
    .out (net45)
  );
  and_cell and20 (
    .a (net22),
    .b (net5),
    .out (net46)
  );
  and_cell and21 (
    .a (net20),
    .b (net3),
    .out (net47)
  );
  and_cell and22 (
    .a (net46),
    .b (net47),
    .out (net48)
  );
  and_cell and23 (
    .a (net48),
    .b (net1),
    .out (net49)
  );
  and_cell and24 (
    .a (net22),
    .b (net5),
    .out (net50)
  );
  and_cell and25 (
    .a (net4),
    .b (net19),
    .out (net51)
  );
  and_cell and26 (
    .a (net50),
    .b (net51),
    .out (net52)
  );
  and_cell and27 (
    .a (net52),
    .b (net18),
    .out (net53)
  );
  or_cell or5 (
    .a (net49),
    .b (net53),
    .out (net54)
  );
  and_cell and28 (
    .a (net6),
    .b (net21),
    .out (net55)
  );
  and_cell and29 (
    .a (net20),
    .b (net3),
    .out (net56)
  );
  and_cell and30 (
    .a (net55),
    .b (net56),
    .out (net57)
  );
  and_cell and31 (
    .a (net57),
    .b (net1),
    .out (net58)
  );
  and_cell and32 (
    .a (net6),
    .b (net21),
    .out (net59)
  );
  and_cell and33 (
    .a (net4),
    .b (net19),
    .out (net60)
  );
  and_cell and34 (
    .a (net59),
    .b (net60),
    .out (net61)
  );
  and_cell and35 (
    .a (net61),
    .b (net18),
    .out (net62)
  );
  or_cell or6 (
    .a (net58),
    .b (net62),
    .out (net63)
  );
  or_cell or7 (
    .a (net44),
    .b (net54),
    .out (net64)
  );
  or_cell or8 (
    .a (net64),
    .b (net63),
    .out (net65)
  );
  or_cell or9 (
    .a (net45),
    .b (net65),
    .out (net7)
  );
  and_cell and36 (
    .a (net22),
    .b (net5),
    .out (net66)
  );
  and_cell and37 (
    .a (net20),
    .b (net19),
    .out (net67)
  );
  and_cell and38 (
    .a (net66),
    .b (net67),
    .out (net68)
  );
  and_cell and39 (
    .a (net22),
    .b (net5),
    .out (net69)
  );
  and_cell and40 (
    .a (net19),
    .b (net18),
    .out (net70)
  );
  and_cell and41 (
    .a (net69),
    .b (net70),
    .out (net71)
  );
  or_cell or10 (
    .a (net68),
    .b (net71),
    .out (net72)
  );
  and_cell and42 (
    .a (net6),
    .b (net21),
    .out (net73)
  );
  and_cell and43 (
    .a (net20),
    .b (net19),
    .out (net74)
  );
  and_cell and44 (
    .a (net73),
    .b (net74),
    .out (net75)
  );
  and_cell and45 (
    .a (net6),
    .b (net21),
    .out (net76)
  );
  and_cell and46 (
    .a (net19),
    .b (net17),
    .out (net77)
  );
  and_cell and47 (
    .a (net76),
    .b (net77),
    .out (net78)
  );
  or_cell or11 (
    .a (net75),
    .b (net78),
    .out (net79)
  );
  or_cell or12 (
    .a (net72),
    .b (net79),
    .out (net80)
  );
  and_cell and48 (
    .a (net22),
    .b (net5),
    .out (net81)
  );
  and_cell and49 (
    .a (net20),
    .b (net18),
    .out (net82)
  );
  and_cell and50 (
    .a (net81),
    .b (net82),
    .out (net83)
  );
  and_cell and51 (
    .a (net83),
    .b (net17),
    .out (net84)
  );
  and_cell and52 (
    .a (net22),
    .b (net5),
    .out (net85)
  );
  and_cell and53 (
    .a (net20),
    .b (net2),
    .out (net86)
  );
  and_cell and54 (
    .a (net85),
    .b (net86),
    .out (net87)
  );
  and_cell and55 (
    .a (net87),
    .b (net1),
    .out (net88)
  );
  or_cell or13 (
    .a (net84),
    .b (net88),
    .out (net89)
  );
  and_cell and56 (
    .a (net6),
    .b (net21),
    .out (net90)
  );
  and_cell and57 (
    .a (net20),
    .b (net18),
    .out (net91)
  );
  and_cell and58 (
    .a (net90),
    .b (net91),
    .out (net92)
  );
  and_cell and59 (
    .a (net92),
    .b (net17),
    .out (net93)
  );
  and_cell and60 (
    .a (net6),
    .b (net21),
    .out (net94)
  );
  and_cell and61 (
    .a (net20),
    .b (net2),
    .out (net95)
  );
  and_cell and62 (
    .a (net94),
    .b (net95),
    .out (net96)
  );
  and_cell and63 (
    .a (net96),
    .b (net1),
    .out (net97)
  );
  or_cell or14 (
    .a (net93),
    .b (net97),
    .out (net98)
  );
  or_cell or15 (
    .a (net89),
    .b (net98),
    .out (net99)
  );
  and_cell and64 (
    .a (net6),
    .b (net21),
    .out (net100)
  );
  and_cell and65 (
    .a (net4),
    .b (net18),
    .out (net101)
  );
  and_cell and66 (
    .a (net100),
    .b (net101),
    .out (net102)
  );
  and_cell and67 (
    .a (net102),
    .b (net1),
    .out (net103)
  );
  or_cell or16 (
    .a (net104),
    .b (net103),
    .out (net8)
  );
  or_cell or17 (
    .a (net80),
    .b (net99),
    .out (net104)
  );
  and_cell and68 (
    .a (net22),
    .b (net5),
    .out (net105)
  );
  and_cell and69 (
    .a (net19),
    .b (net18),
    .out (net106)
  );
  and_cell and70 (
    .a (net105),
    .b (net106),
    .out (net107)
  );
  and_cell and71 (
    .a (net22),
    .b (net5),
    .out (net108)
  );
  and_cell and72 (
    .a (net20),
    .b (net1),
    .out (net109)
  );
  and_cell and73 (
    .a (net108),
    .b (net109),
    .out (net110)
  );
  or_cell or18 (
    .a (net107),
    .b (net110),
    .out (net111)
  );
  and_cell and74 (
    .a (net22),
    .b (net5),
    .out (net112)
  );
  and_cell and75 (
    .a (net20),
    .b (net3),
    .out (net113)
  );
  and_cell and76 (
    .a (net112),
    .b (net113),
    .out (net114)
  );
  and_cell and77 (
    .a (net6),
    .b (net21),
    .out (net115)
  );
  and_cell and78 (
    .a (net20),
    .b (net18),
    .out (net116)
  );
  and_cell and79 (
    .a (net115),
    .b (net116),
    .out (net117)
  );
  or_cell or19 (
    .a (net114),
    .b (net117),
    .out (net118)
  );
  or_cell or20 (
    .a (net111),
    .b (net118),
    .out (net119)
  );
  and_cell and80 (
    .a (net6),
    .b (net21),
    .out (net120)
  );
  and_cell and81 (
    .a (net20),
    .b (net1),
    .out (net121)
  );
  and_cell and82 (
    .a (net120),
    .b (net121),
    .out (net122)
  );
  and_cell and83 (
    .a (net6),
    .b (net21),
    .out (net123)
  );
  and_cell and84 (
    .a (net18),
    .b (net1),
    .out (net124)
  );
  and_cell and85 (
    .a (net123),
    .b (net124),
    .out (net125)
  );
  or_cell or21 (
    .a (net122),
    .b (net125),
    .out (net126)
  );
  and_cell and86 (
    .a (net6),
    .b (net21),
    .out (net127)
  );
  and_cell and87 (
    .a (net20),
    .b (net3),
    .out (net128)
  );
  and_cell and88 (
    .a (net127),
    .b (net128),
    .out (net129)
  );
  and_cell and89 (
    .a (net6),
    .b (net21),
    .out (net130)
  );
  and_cell and90 (
    .a (net4),
    .b (net19),
    .out (net131)
  );
  and_cell and91 (
    .a (net130),
    .b (net131),
    .out (net132)
  );
  or_cell or22 (
    .a (net129),
    .b (net132),
    .out (net133)
  );
  or_cell or23 (
    .a (net126),
    .b (net133),
    .out (net134)
  );
  or_cell or24 (
    .a (net119),
    .b (net134),
    .out (net9)
  );
  and_cell and92 (
    .a (net6),
    .b (net21),
    .out (net135)
  );
  and_cell and93 (
    .a (net4),
    .b (net18),
    .out (net136)
  );
  and_cell and94 (
    .a (net135),
    .b (net136),
    .out (net137)
  );
  or_cell or25 (
    .a (net137),
    .b (net138),
    .out (net139)
  );
  and_cell and95 (
    .a (net22),
    .b (net5),
    .out (net140)
  );
  and_cell and96 (
    .a (net20),
    .b (net19),
    .out (net141)
  );
  and_cell and97 (
    .a (net140),
    .b (net141),
    .out (net142)
  );
  and_cell and98 (
    .a (net142),
    .b (net17),
    .out (net138)
  );
  and_cell and99 (
    .a (net22),
    .b (net5),
    .out (net143)
  );
  and_cell and100 (
    .a (net20),
    .b (net19),
    .out (net144)
  );
  and_cell and101 (
    .a (net143),
    .b (net144),
    .out (net145)
  );
  and_cell and102 (
    .a (net145),
    .b (net2),
    .out (net146)
  );
  and_cell and103 (
    .a (net22),
    .b (net5),
    .out (net147)
  );
  and_cell and104 (
    .a (net20),
    .b (net2),
    .out (net148)
  );
  and_cell and105 (
    .a (net147),
    .b (net148),
    .out (net149)
  );
  and_cell and106 (
    .a (net149),
    .b (net17),
    .out (net150)
  );
  or_cell or26 (
    .a (net146),
    .b (net150),
    .out (net151)
  );
  and_cell and107 (
    .a (net22),
    .b (net5),
    .out (net152)
  );
  and_cell and108 (
    .a (net4),
    .b (net19),
    .out (net153)
  );
  and_cell and109 (
    .a (net152),
    .b (net153),
    .out (net154)
  );
  and_cell and110 (
    .a (net154),
    .b (net18),
    .out (net155)
  );
  and_cell and111 (
    .a (net6),
    .b (net21),
    .out (net156)
  );
  and_cell and112 (
    .a (net20),
    .b (net19),
    .out (net157)
  );
  and_cell and113 (
    .a (net156),
    .b (net157),
    .out (net158)
  );
  and_cell and114 (
    .a (net158),
    .b (net17),
    .out (net159)
  );
  or_cell or27 (
    .a (net155),
    .b (net159),
    .out (net160)
  );
  and_cell and115 (
    .a (net6),
    .b (net21),
    .out (net161)
  );
  and_cell and116 (
    .a (net19),
    .b (net2),
    .out (net162)
  );
  and_cell and117 (
    .a (net161),
    .b (net162),
    .out (net163)
  );
  and_cell and118 (
    .a (net163),
    .b (net1),
    .out (net164)
  );
  and_cell and119 (
    .a (net6),
    .b (net21),
    .out (net165)
  );
  and_cell and120 (
    .a (net3),
    .b (net18),
    .out (net166)
  );
  and_cell and121 (
    .a (net165),
    .b (net166),
    .out (net167)
  );
  and_cell and122 (
    .a (net167),
    .b (net1),
    .out (net168)
  );
  or_cell or28 (
    .a (net164),
    .b (net168),
    .out (net169)
  );
  and_cell and123 (
    .a (net6),
    .b (net21),
    .out (net170)
  );
  and_cell and124 (
    .a (net3),
    .b (net2),
    .out (net171)
  );
  and_cell and125 (
    .a (net170),
    .b (net171),
    .out (net172)
  );
  and_cell and126 (
    .a (net172),
    .b (net17),
    .out (net173)
  );
  and_cell and127 (
    .a (net22),
    .b (net5),
    .out (net174)
  );
  and_cell and128 (
    .a (net20),
    .b (net3),
    .out (net175)
  );
  and_cell and129 (
    .a (net174),
    .b (net175),
    .out (net176)
  );
  and_cell and130 (
    .a (net176),
    .b (net177),
    .out (net178)
  );
  or_cell or29 (
    .a (net173),
    .b (net178),
    .out (net179)
  );
  and_cell and131 (
    .a (net18),
    .b (net1),
    .out (net177)
  );
  or_cell or30 (
    .a (net169),
    .b (net179),
    .out (net180)
  );
  or_cell or31 (
    .a (net151),
    .b (net160),
    .out (net181)
  );
  or_cell or32 (
    .a (net181),
    .b (net180),
    .out (net182)
  );
  or_cell or33 (
    .a (net139),
    .b (net182),
    .out (net10)
  );
  and_cell and132 (
    .a (net6),
    .b (net21),
    .out (net183)
  );
  and_cell and133 (
    .a (net19),
    .b (net17),
    .out (net184)
  );
  and_cell and134 (
    .a (net183),
    .b (net184),
    .out (net185)
  );
  or_cell or34 (
    .a (net185),
    .b (net186),
    .out (net187)
  );
  and_cell and135 (
    .a (net22),
    .b (net5),
    .out (net188)
  );
  and_cell and136 (
    .a (net19),
    .b (net18),
    .out (net189)
  );
  and_cell and137 (
    .a (net188),
    .b (net189),
    .out (net190)
  );
  and_cell and138 (
    .a (net190),
    .b (net17),
    .out (net191)
  );
  and_cell and139 (
    .a (net22),
    .b (net5),
    .out (net192)
  );
  and_cell and140 (
    .a (net20),
    .b (net2),
    .out (net193)
  );
  and_cell and141 (
    .a (net192),
    .b (net193),
    .out (net194)
  );
  and_cell and142 (
    .a (net194),
    .b (net17),
    .out (net195)
  );
  or_cell or35 (
    .a (net191),
    .b (net195),
    .out (net196)
  );
  and_cell and143 (
    .a (net6),
    .b (net21),
    .out (net197)
  );
  and_cell and144 (
    .a (net2),
    .b (net17),
    .out (net198)
  );
  and_cell and145 (
    .a (net197),
    .b (net198),
    .out (net186)
  );
  and_cell and146 (
    .a (net6),
    .b (net21),
    .out (net199)
  );
  and_cell and147 (
    .a (net4),
    .b (net2),
    .out (net200)
  );
  and_cell and148 (
    .a (net199),
    .b (net200),
    .out (net201)
  );
  or_cell or36 (
    .a (net201),
    .b (net202),
    .out (net203)
  );
  and_cell and149 (
    .a (net6),
    .b (net21),
    .out (net204)
  );
  and_cell and150 (
    .a (net4),
    .b (net3),
    .out (net205)
  );
  and_cell and151 (
    .a (net204),
    .b (net205),
    .out (net202)
  );
  or_cell or37 (
    .a (net203),
    .b (net196),
    .out (net206)
  );
  or_cell or38 (
    .a (net187),
    .b (net206),
    .out (net11)
  );
  and_cell and152 (
    .a (net6),
    .b (net21),
    .out (net207)
  );
  and_cell and153 (
    .a (net18),
    .b (net17),
    .out (net208)
  );
  and_cell and154 (
    .a (net207),
    .b (net208),
    .out (net209)
  );
  or_cell or39 (
    .a (net209),
    .b (net210),
    .out (net211)
  );
  and_cell and155 (
    .a (net6),
    .b (net21),
    .out (net212)
  );
  and_cell and156 (
    .a (net3),
    .b (net17),
    .out (net213)
  );
  and_cell and157 (
    .a (net212),
    .b (net213),
    .out (net210)
  );
  and_cell and158 (
    .a (net6),
    .b (net21),
    .out (net214)
  );
  and_cell and159 (
    .a (net4),
    .b (net19),
    .out (net215)
  );
  and_cell and160 (
    .a (net214),
    .b (net215),
    .out (net216)
  );
  or_cell or40 (
    .a (net216),
    .b (net217),
    .out (net218)
  );
  and_cell and161 (
    .a (net6),
    .b (net21),
    .out (net219)
  );
  and_cell and162 (
    .a (net4),
    .b (net2),
    .out (net220)
  );
  and_cell and163 (
    .a (net219),
    .b (net220),
    .out (net217)
  );
  and_cell and164 (
    .a (net22),
    .b (net5),
    .out (net221)
  );
  and_cell and165 (
    .a (net20),
    .b (net18),
    .out (net222)
  );
  and_cell and166 (
    .a (net221),
    .b (net222),
    .out (net223)
  );
  and_cell and167 (
    .a (net223),
    .b (net17),
    .out (net224)
  );
  and_cell and168 (
    .a (net22),
    .b (net5),
    .out (net225)
  );
  and_cell and169 (
    .a (net20),
    .b (net3),
    .out (net226)
  );
  and_cell and170 (
    .a (net225),
    .b (net226),
    .out (net227)
  );
  and_cell and171 (
    .a (net227),
    .b (net18),
    .out (net228)
  );
  or_cell or41 (
    .a (net224),
    .b (net228),
    .out (net229)
  );
  and_cell and172 (
    .a (net22),
    .b (net5),
    .out (net230)
  );
  and_cell and173 (
    .a (net20),
    .b (net3),
    .out (net231)
  );
  and_cell and174 (
    .a (net230),
    .b (net231),
    .out (net232)
  );
  and_cell and175 (
    .a (net232),
    .b (net17),
    .out (net233)
  );
  and_cell and176 (
    .a (net22),
    .b (net5),
    .out (net234)
  );
  and_cell and177 (
    .a (net4),
    .b (net19),
    .out (net235)
  );
  and_cell and178 (
    .a (net234),
    .b (net235),
    .out (net236)
  );
  and_cell and179 (
    .a (net236),
    .b (net18),
    .out (net237)
  );
  or_cell or42 (
    .a (net233),
    .b (net237),
    .out (net238)
  );
  and_cell and180 (
    .a (net6),
    .b (net21),
    .out (net239)
  );
  and_cell and181 (
    .a (net20),
    .b (net3),
    .out (net240)
  );
  and_cell and182 (
    .a (net239),
    .b (net240),
    .out (net241)
  );
  and_cell and183 (
    .a (net241),
    .b (net18),
    .out (net242)
  );
  or_cell or43 (
    .a (net238),
    .b (net242),
    .out (net243)
  );
  or_cell or44 (
    .a (net229),
    .b (net243),
    .out (net244)
  );
  or_cell or45 (
    .a (net211),
    .b (net218),
    .out (net245)
  );
  or_cell or46 (
    .a (net245),
    .b (net244),
    .out (net12)
  );
  and_cell and184 (
    .a (net6),
    .b (net21),
    .out (net246)
  );
  and_cell and185 (
    .a (net19),
    .b (net2),
    .out (net247)
  );
  and_cell and186 (
    .a (net246),
    .b (net247),
    .out (net248)
  );
  or_cell or47 (
    .a (net248),
    .b (net249),
    .out (net250)
  );
  and_cell and187 (
    .a (net6),
    .b (net21),
    .out (net251)
  );
  and_cell and188 (
    .a (net2),
    .b (net17),
    .out (net252)
  );
  and_cell and189 (
    .a (net251),
    .b (net252),
    .out (net249)
  );
  and_cell and190 (
    .a (net6),
    .b (net21),
    .out (net253)
  );
  and_cell and191 (
    .a (net4),
    .b (net19),
    .out (net254)
  );
  and_cell and192 (
    .a (net253),
    .b (net254),
    .out (net255)
  );
  or_cell or48 (
    .a (net255),
    .b (net256),
    .out (net257)
  );
  and_cell and193 (
    .a (net6),
    .b (net21),
    .out (net258)
  );
  and_cell and194 (
    .a (net4),
    .b (net1),
    .out (net259)
  );
  and_cell and195 (
    .a (net258),
    .b (net259),
    .out (net256)
  );
  and_cell and196 (
    .a (net22),
    .b (net5),
    .out (net260)
  );
  and_cell and197 (
    .a (net20),
    .b (net19),
    .out (net261)
  );
  and_cell and198 (
    .a (net260),
    .b (net261),
    .out (net262)
  );
  and_cell and199 (
    .a (net262),
    .b (net2),
    .out (net263)
  );
  and_cell and200 (
    .a (net22),
    .b (net5),
    .out (net264)
  );
  and_cell and201 (
    .a (net20),
    .b (net2),
    .out (net265)
  );
  and_cell and202 (
    .a (net264),
    .b (net265),
    .out (net266)
  );
  and_cell and203 (
    .a (net266),
    .b (net17),
    .out (net267)
  );
  or_cell or49 (
    .a (net263),
    .b (net267),
    .out (net268)
  );
  and_cell and204 (
    .a (net22),
    .b (net5),
    .out (net269)
  );
  and_cell and205 (
    .a (net20),
    .b (net3),
    .out (net270)
  );
  and_cell and206 (
    .a (net269),
    .b (net270),
    .out (net271)
  );
  and_cell and207 (
    .a (net271),
    .b (net18),
    .out (net272)
  );
  and_cell and208 (
    .a (net22),
    .b (net5),
    .out (net273)
  );
  and_cell and209 (
    .a (net4),
    .b (net19),
    .out (net274)
  );
  and_cell and210 (
    .a (net273),
    .b (net274),
    .out (net275)
  );
  and_cell and211 (
    .a (net275),
    .b (net18),
    .out (net276)
  );
  or_cell or50 (
    .a (net272),
    .b (net276),
    .out (net277)
  );
  and_cell and212 (
    .a (net6),
    .b (net21),
    .out (net278)
  );
  and_cell and213 (
    .a (net20),
    .b (net3),
    .out (net279)
  );
  and_cell and214 (
    .a (net278),
    .b (net279),
    .out (net280)
  );
  and_cell and215 (
    .a (net280),
    .b (net18),
    .out (net281)
  );
  or_cell or51 (
    .a (net277),
    .b (net281),
    .out (net282)
  );
  or_cell or52 (
    .a (net268),
    .b (net282),
    .out (net283)
  );
  or_cell or53 (
    .a (net250),
    .b (net257),
    .out (net284)
  );
  or_cell or54 (
    .a (net284),
    .b (net283),
    .out (net13)
  );
  and_cell and216 (
    .a (net22),
    .b (net5),
    .out (net14)
  );
endmodule
