magic
tech sky130A
magscale 1 2
timestamp 1682329530
<< viali >>
rect 2421 17221 2455 17255
rect 3249 17221 3283 17255
rect 11805 17221 11839 17255
rect 38853 17221 38887 17255
rect 1593 17153 1627 17187
rect 4629 17153 4663 17187
rect 6745 17153 6779 17187
rect 8033 17153 8067 17187
rect 9965 17153 9999 17187
rect 13185 17153 13219 17187
rect 14473 17153 14507 17187
rect 16865 17153 16899 17187
rect 19625 17153 19659 17187
rect 22845 17153 22879 17187
rect 24777 17153 24811 17187
rect 26065 17153 26099 17187
rect 27997 17153 28031 17187
rect 29929 17153 29963 17187
rect 31217 17153 31251 17187
rect 32321 17153 32355 17187
rect 35081 17153 35115 17187
rect 35725 17153 35759 17187
rect 37657 17153 37691 17187
rect 42809 17153 42843 17187
rect 43453 17153 43487 17187
rect 44097 17153 44131 17187
rect 4905 17085 4939 17119
rect 32597 17085 32631 17119
rect 3433 17017 3467 17051
rect 11989 17017 12023 17051
rect 1777 16949 1811 16983
rect 2513 16949 2547 16983
rect 9781 16949 9815 16983
rect 17049 16949 17083 16983
rect 24593 16949 24627 16983
rect 31033 16949 31067 16983
rect 34897 16949 34931 16983
rect 38945 16949 38979 16983
rect 44373 16745 44407 16779
rect 1869 16609 1903 16643
rect 1685 16541 1719 16575
rect 7021 16541 7055 16575
rect 19993 16541 20027 16575
rect 20913 16541 20947 16575
rect 8125 16473 8159 16507
rect 1777 16065 1811 16099
rect 36001 16065 36035 16099
rect 36093 15997 36127 16031
rect 36185 15997 36219 16031
rect 35633 15861 35667 15895
rect 44373 15861 44407 15895
rect 19533 15657 19567 15691
rect 35725 15657 35759 15691
rect 11529 15589 11563 15623
rect 11989 15521 12023 15555
rect 20085 15521 20119 15555
rect 36277 15521 36311 15555
rect 44005 15521 44039 15555
rect 10149 15453 10183 15487
rect 10405 15453 10439 15487
rect 17601 15453 17635 15487
rect 17785 15453 17819 15487
rect 25237 15453 25271 15487
rect 42809 15453 42843 15487
rect 19901 15385 19935 15419
rect 36093 15385 36127 15419
rect 12633 15317 12667 15351
rect 17969 15317 18003 15351
rect 19993 15317 20027 15351
rect 25053 15317 25087 15351
rect 36185 15317 36219 15351
rect 16313 15113 16347 15147
rect 18521 15113 18555 15147
rect 20361 15113 20395 15147
rect 32321 15113 32355 15147
rect 32689 15113 32723 15147
rect 33977 15113 34011 15147
rect 19226 15045 19260 15079
rect 34866 15045 34900 15079
rect 6745 14977 6779 15011
rect 7389 14977 7423 15011
rect 11897 14977 11931 15011
rect 12164 14977 12198 15011
rect 14933 14977 14967 15011
rect 15200 14977 15234 15011
rect 17141 14977 17175 15011
rect 17397 14977 17431 15011
rect 18981 14977 19015 15011
rect 21005 14977 21039 15011
rect 23029 14977 23063 15011
rect 23285 14977 23319 15011
rect 24869 14977 24903 15011
rect 25136 14977 25170 15011
rect 28805 14977 28839 15011
rect 30757 14977 30791 15011
rect 31401 14977 31435 15011
rect 32781 14977 32815 15011
rect 34161 14977 34195 15011
rect 36645 14977 36679 15011
rect 40049 14977 40083 15011
rect 28549 14909 28583 14943
rect 32873 14909 32907 14943
rect 34621 14909 34655 14943
rect 39865 14909 39899 14943
rect 20821 14841 20855 14875
rect 36001 14841 36035 14875
rect 6561 14773 6595 14807
rect 7205 14773 7239 14807
rect 13277 14773 13311 14807
rect 24409 14773 24443 14807
rect 26249 14773 26283 14807
rect 29929 14773 29963 14807
rect 30573 14773 30607 14807
rect 31217 14773 31251 14807
rect 36461 14773 36495 14807
rect 40233 14773 40267 14807
rect 5641 14569 5675 14603
rect 6469 14569 6503 14603
rect 17509 14569 17543 14603
rect 25053 14569 25087 14603
rect 30113 14569 30147 14603
rect 33609 14569 33643 14603
rect 36737 14569 36771 14603
rect 41429 14569 41463 14603
rect 6653 14501 6687 14535
rect 12909 14501 12943 14535
rect 15301 14501 15335 14535
rect 18153 14501 18187 14535
rect 29193 14501 29227 14535
rect 36277 14501 36311 14535
rect 11529 14433 11563 14467
rect 15945 14433 15979 14467
rect 18797 14433 18831 14467
rect 20085 14433 20119 14467
rect 23765 14433 23799 14467
rect 23857 14433 23891 14467
rect 25605 14433 25639 14467
rect 26709 14433 26743 14467
rect 26801 14433 26835 14467
rect 34069 14433 34103 14467
rect 34161 14433 34195 14467
rect 37381 14433 37415 14467
rect 4721 14365 4755 14399
rect 4905 14365 4939 14399
rect 5641 14365 5675 14399
rect 5825 14365 5859 14399
rect 7113 14365 7147 14399
rect 7369 14365 7403 14399
rect 11069 14365 11103 14399
rect 13369 14365 13403 14399
rect 14289 14365 14323 14399
rect 14473 14365 14507 14399
rect 15669 14365 15703 14399
rect 17693 14365 17727 14399
rect 19809 14365 19843 14399
rect 22109 14365 22143 14399
rect 25421 14365 25455 14399
rect 26617 14365 26651 14399
rect 27813 14365 27847 14399
rect 29745 14365 29779 14399
rect 29929 14365 29963 14399
rect 31033 14365 31067 14399
rect 31289 14365 31323 14399
rect 34897 14365 34931 14399
rect 37105 14365 37139 14399
rect 39497 14365 39531 14399
rect 40049 14365 40083 14399
rect 42809 14365 42843 14399
rect 6285 14297 6319 14331
rect 11774 14297 11808 14331
rect 14381 14297 14415 14331
rect 15761 14297 15795 14331
rect 23673 14297 23707 14331
rect 28058 14297 28092 14331
rect 33977 14297 34011 14331
rect 35164 14297 35198 14331
rect 40294 14297 40328 14331
rect 44005 14297 44039 14331
rect 4813 14229 4847 14263
rect 6495 14229 6529 14263
rect 8493 14229 8527 14263
rect 10885 14229 10919 14263
rect 13461 14229 13495 14263
rect 18521 14229 18555 14263
rect 18613 14229 18647 14263
rect 19441 14229 19475 14263
rect 19901 14229 19935 14263
rect 21925 14229 21959 14263
rect 23305 14229 23339 14263
rect 25513 14229 25547 14263
rect 26249 14229 26283 14263
rect 32413 14229 32447 14263
rect 37197 14229 37231 14263
rect 39313 14229 39347 14263
rect 5273 14025 5307 14059
rect 6009 14025 6043 14059
rect 7941 14025 7975 14059
rect 12265 14025 12299 14059
rect 14933 14025 14967 14059
rect 15393 14025 15427 14059
rect 17877 14025 17911 14059
rect 19901 14025 19935 14059
rect 20729 14025 20763 14059
rect 20821 14025 20855 14059
rect 23397 14025 23431 14059
rect 24225 14025 24259 14059
rect 24317 14025 24351 14059
rect 30205 14025 30239 14059
rect 31309 14025 31343 14059
rect 34437 14025 34471 14059
rect 36277 14025 36311 14059
rect 36369 14025 36403 14059
rect 37473 14025 37507 14059
rect 37841 14025 37875 14059
rect 40141 14025 40175 14059
rect 41337 14025 41371 14059
rect 6828 13957 6862 13991
rect 8401 13957 8435 13991
rect 12081 13957 12115 13991
rect 13820 13957 13854 13991
rect 18766 13957 18800 13991
rect 22262 13957 22296 13991
rect 41705 13957 41739 13991
rect 3065 13889 3099 13923
rect 4997 13889 5031 13923
rect 5733 13889 5767 13923
rect 6561 13889 6595 13923
rect 8585 13889 8619 13923
rect 10977 13889 11011 13923
rect 11161 13889 11195 13923
rect 11713 13889 11747 13923
rect 12909 13889 12943 13923
rect 13553 13889 13587 13923
rect 15577 13889 15611 13923
rect 18061 13889 18095 13923
rect 22017 13889 22051 13923
rect 30021 13889 30055 13923
rect 31493 13889 31527 13923
rect 33057 13889 33091 13923
rect 33313 13889 33347 13923
rect 35449 13889 35483 13923
rect 38761 13889 38795 13923
rect 39017 13889 39051 13923
rect 1777 13821 1811 13855
rect 3341 13821 3375 13855
rect 5273 13821 5307 13855
rect 6009 13821 6043 13855
rect 12725 13821 12759 13855
rect 18521 13821 18555 13855
rect 21005 13821 21039 13855
rect 24501 13821 24535 13855
rect 29837 13821 29871 13855
rect 36461 13821 36495 13855
rect 37933 13821 37967 13855
rect 38117 13821 38151 13855
rect 41797 13821 41831 13855
rect 41889 13821 41923 13855
rect 5089 13753 5123 13787
rect 23857 13753 23891 13787
rect 35265 13753 35299 13787
rect 35909 13753 35943 13787
rect 5825 13685 5859 13719
rect 8769 13685 8803 13719
rect 11069 13685 11103 13719
rect 12081 13685 12115 13719
rect 13093 13685 13127 13719
rect 20361 13685 20395 13719
rect 5365 13481 5399 13515
rect 6009 13481 6043 13515
rect 7021 13481 7055 13515
rect 12541 13481 12575 13515
rect 13645 13481 13679 13515
rect 14657 13481 14691 13515
rect 15301 13481 15335 13515
rect 15485 13481 15519 13515
rect 18889 13481 18923 13515
rect 19441 13481 19475 13515
rect 21649 13481 21683 13515
rect 37749 13481 37783 13515
rect 7205 13413 7239 13447
rect 11253 13413 11287 13447
rect 8033 13345 8067 13379
rect 12633 13345 12667 13379
rect 19993 13345 20027 13379
rect 22201 13345 22235 13379
rect 23949 13345 23983 13379
rect 3433 13277 3467 13311
rect 3985 13277 4019 13311
rect 6653 13277 6687 13311
rect 7757 13277 7791 13311
rect 7849 13277 7883 13311
rect 11253 13277 11287 13311
rect 11437 13277 11471 13311
rect 12081 13277 12115 13311
rect 12817 13277 12851 13311
rect 13553 13277 13587 13311
rect 14289 13277 14323 13311
rect 14473 13277 14507 13311
rect 17509 13277 17543 13311
rect 19901 13277 19935 13311
rect 22109 13277 22143 13311
rect 23673 13277 23707 13311
rect 24777 13277 24811 13311
rect 27905 13277 27939 13311
rect 28181 13277 28215 13311
rect 28825 13277 28859 13311
rect 30757 13277 30791 13311
rect 32781 13277 32815 13311
rect 36369 13277 36403 13311
rect 36625 13277 36659 13311
rect 38393 13277 38427 13311
rect 4230 13209 4264 13243
rect 5825 13209 5859 13243
rect 6025 13209 6059 13243
rect 7021 13209 7055 13243
rect 12541 13209 12575 13243
rect 15117 13209 15151 13243
rect 15317 13209 15351 13243
rect 17776 13209 17810 13243
rect 25044 13209 25078 13243
rect 27721 13209 27755 13243
rect 31024 13209 31058 13243
rect 3249 13141 3283 13175
rect 6193 13141 6227 13175
rect 11897 13141 11931 13175
rect 13001 13141 13035 13175
rect 19809 13141 19843 13175
rect 22017 13141 22051 13175
rect 23305 13141 23339 13175
rect 23765 13141 23799 13175
rect 26157 13141 26191 13175
rect 28089 13141 28123 13175
rect 28641 13141 28675 13175
rect 32137 13141 32171 13175
rect 32597 13141 32631 13175
rect 38209 13141 38243 13175
rect 3525 12937 3559 12971
rect 4537 12937 4571 12971
rect 11069 12937 11103 12971
rect 12541 12937 12575 12971
rect 14381 12937 14415 12971
rect 18889 12937 18923 12971
rect 30205 12937 30239 12971
rect 31493 12937 31527 12971
rect 5641 12869 5675 12903
rect 5857 12869 5891 12903
rect 6929 12869 6963 12903
rect 9505 12869 9539 12903
rect 12173 12869 12207 12903
rect 12265 12869 12299 12903
rect 28273 12869 28307 12903
rect 31309 12869 31343 12903
rect 40417 12869 40451 12903
rect 3341 12801 3375 12835
rect 4353 12801 4387 12835
rect 4537 12801 4571 12835
rect 5181 12801 5215 12835
rect 6561 12801 6595 12835
rect 6745 12801 6779 12835
rect 7389 12801 7423 12835
rect 9413 12801 9447 12835
rect 10977 12801 11011 12835
rect 11161 12801 11195 12835
rect 11897 12801 11931 12835
rect 11990 12801 12024 12835
rect 12362 12801 12396 12835
rect 13001 12801 13035 12835
rect 13257 12801 13291 12835
rect 14841 12801 14875 12835
rect 17509 12801 17543 12835
rect 17776 12801 17810 12835
rect 19349 12801 19383 12835
rect 19605 12801 19639 12835
rect 22753 12801 22787 12835
rect 23213 12801 23247 12835
rect 26617 12801 26651 12835
rect 27169 12801 27203 12835
rect 27997 12801 28031 12835
rect 30389 12801 30423 12835
rect 32505 12801 32539 12835
rect 33333 12801 33367 12835
rect 36093 12801 36127 12835
rect 36185 12801 36219 12835
rect 36829 12801 36863 12835
rect 37657 12801 37691 12835
rect 38393 12801 38427 12835
rect 41061 12801 41095 12835
rect 3157 12733 3191 12767
rect 23489 12733 23523 12767
rect 27261 12733 27295 12767
rect 31585 12733 31619 12767
rect 32321 12733 32355 12767
rect 38669 12733 38703 12767
rect 6009 12665 6043 12699
rect 7481 12665 7515 12699
rect 20729 12665 20763 12699
rect 22569 12665 22603 12699
rect 29745 12665 29779 12699
rect 32689 12665 32723 12699
rect 4997 12597 5031 12631
rect 5825 12597 5859 12631
rect 14933 12597 14967 12631
rect 24961 12597 24995 12631
rect 26433 12597 26467 12631
rect 31033 12597 31067 12631
rect 33149 12597 33183 12631
rect 36645 12597 36679 12631
rect 37473 12597 37507 12631
rect 40877 12597 40911 12631
rect 44373 12597 44407 12631
rect 6929 12393 6963 12427
rect 10609 12393 10643 12427
rect 11713 12393 11747 12427
rect 13277 12393 13311 12427
rect 14289 12393 14323 12427
rect 16681 12393 16715 12427
rect 17877 12393 17911 12427
rect 23305 12393 23339 12427
rect 24593 12393 24627 12427
rect 27905 12393 27939 12427
rect 28641 12393 28675 12427
rect 30297 12393 30331 12427
rect 33425 12393 33459 12427
rect 38945 12393 38979 12427
rect 40049 12393 40083 12427
rect 10149 12325 10183 12359
rect 13185 12325 13219 12359
rect 14841 12325 14875 12359
rect 17049 12325 17083 12359
rect 28825 12325 28859 12359
rect 9873 12257 9907 12291
rect 10793 12257 10827 12291
rect 11897 12257 11931 12291
rect 12265 12257 12299 12291
rect 13369 12257 13403 12291
rect 13737 12257 13771 12291
rect 23857 12257 23891 12291
rect 25329 12257 25363 12291
rect 26157 12257 26191 12291
rect 37197 12257 37231 12291
rect 41521 12257 41555 12291
rect 3433 12189 3467 12223
rect 3985 12189 4019 12223
rect 4169 12189 4203 12223
rect 4813 12189 4847 12223
rect 4997 12189 5031 12223
rect 5089 12189 5123 12223
rect 5549 12189 5583 12223
rect 5816 12189 5850 12223
rect 7665 12189 7699 12223
rect 9781 12189 9815 12223
rect 10885 12189 10919 12223
rect 11989 12189 12023 12223
rect 12817 12189 12851 12223
rect 14414 12189 14448 12223
rect 14933 12189 14967 12223
rect 16865 12189 16899 12223
rect 17141 12189 17175 12223
rect 18061 12189 18095 12223
rect 21005 12189 21039 12223
rect 21465 12189 21499 12223
rect 21741 12189 21775 12223
rect 22385 12189 22419 12223
rect 24777 12189 24811 12223
rect 25237 12189 25271 12223
rect 28365 12189 28399 12223
rect 28549 12189 28583 12223
rect 28641 12189 28675 12223
rect 30481 12189 30515 12223
rect 30757 12189 30791 12223
rect 31217 12189 31251 12223
rect 33609 12189 33643 12223
rect 34345 12189 34379 12223
rect 34897 12189 34931 12223
rect 40233 12189 40267 12223
rect 41245 12189 41279 12223
rect 4629 12121 4663 12155
rect 11161 12121 11195 12155
rect 11253 12121 11287 12155
rect 12357 12121 12391 12155
rect 23673 12121 23707 12155
rect 26433 12121 26467 12155
rect 30665 12121 30699 12155
rect 31493 12121 31527 12155
rect 35173 12121 35207 12155
rect 37473 12121 37507 12155
rect 3249 12053 3283 12087
rect 4077 12053 4111 12087
rect 7757 12053 7791 12087
rect 14473 12053 14507 12087
rect 20821 12053 20855 12087
rect 22201 12053 22235 12087
rect 23765 12053 23799 12087
rect 32965 12053 32999 12087
rect 34161 12053 34195 12087
rect 36645 12053 36679 12087
rect 6009 11849 6043 11883
rect 11161 11849 11195 11883
rect 12725 11849 12759 11883
rect 16865 11849 16899 11883
rect 18061 11849 18095 11883
rect 18705 11849 18739 11883
rect 20729 11849 20763 11883
rect 21097 11849 21131 11883
rect 22017 11849 22051 11883
rect 22477 11849 22511 11883
rect 26433 11849 26467 11883
rect 32689 11849 32723 11883
rect 36553 11849 36587 11883
rect 10793 11781 10827 11815
rect 27813 11781 27847 11815
rect 29193 11781 29227 11815
rect 30941 11781 30975 11815
rect 35725 11781 35759 11815
rect 40960 11781 40994 11815
rect 2145 11713 2179 11747
rect 3801 11713 3835 11747
rect 4057 11713 4091 11747
rect 5733 11713 5767 11747
rect 5825 11713 5859 11747
rect 6929 11713 6963 11747
rect 7021 11713 7055 11747
rect 10609 11713 10643 11747
rect 10885 11713 10919 11747
rect 10977 11713 11011 11747
rect 11989 11713 12023 11747
rect 12173 11713 12207 11747
rect 12357 11713 12391 11747
rect 12541 11713 12575 11747
rect 13553 11713 13587 11747
rect 13645 11713 13679 11747
rect 17233 11713 17267 11747
rect 17325 11713 17359 11747
rect 18245 11713 18279 11747
rect 18889 11713 18923 11747
rect 22385 11713 22419 11747
rect 26617 11713 26651 11747
rect 27445 11713 27479 11747
rect 27629 11713 27663 11747
rect 29009 11713 29043 11747
rect 30021 11713 30055 11747
rect 30665 11713 30699 11747
rect 30849 11713 30883 11747
rect 31033 11713 31067 11747
rect 32321 11713 32355 11747
rect 32505 11713 32539 11747
rect 35633 11713 35667 11747
rect 36277 11713 36311 11747
rect 36369 11713 36403 11747
rect 36645 11713 36679 11747
rect 37473 11713 37507 11747
rect 38393 11713 38427 11747
rect 38660 11713 38694 11747
rect 40693 11713 40727 11747
rect 2789 11645 2823 11679
rect 7113 11645 7147 11679
rect 12265 11645 12299 11679
rect 13737 11645 13771 11679
rect 17509 11645 17543 11679
rect 21189 11645 21223 11679
rect 21373 11645 21407 11679
rect 22661 11645 22695 11679
rect 36461 11645 36495 11679
rect 37565 11645 37599 11679
rect 5181 11577 5215 11611
rect 13185 11577 13219 11611
rect 6561 11509 6595 11543
rect 30113 11509 30147 11543
rect 31217 11509 31251 11543
rect 32505 11509 32539 11543
rect 39773 11509 39807 11543
rect 42073 11509 42107 11543
rect 3433 11305 3467 11339
rect 5365 11305 5399 11339
rect 7297 11305 7331 11339
rect 10793 11305 10827 11339
rect 11989 11305 12023 11339
rect 13461 11305 13495 11339
rect 17693 11305 17727 11339
rect 20085 11305 20119 11339
rect 23213 11305 23247 11339
rect 32689 11305 32723 11339
rect 38853 11305 38887 11339
rect 40417 11305 40451 11339
rect 41429 11305 41463 11339
rect 7757 11237 7791 11271
rect 16865 11237 16899 11271
rect 22477 11237 22511 11271
rect 30297 11237 30331 11271
rect 37749 11237 37783 11271
rect 38301 11237 38335 11271
rect 4629 11169 4663 11203
rect 11253 11169 11287 11203
rect 11437 11169 11471 11203
rect 12633 11169 12667 11203
rect 17325 11169 17359 11203
rect 20729 11169 20763 11203
rect 21005 11169 21039 11203
rect 25145 11169 25179 11203
rect 25421 11169 25455 11203
rect 26893 11169 26927 11203
rect 27353 11169 27387 11203
rect 29101 11169 29135 11203
rect 31217 11169 31251 11203
rect 41889 11169 41923 11203
rect 41981 11169 42015 11203
rect 2053 11101 2087 11135
rect 4353 11101 4387 11135
rect 5181 11101 5215 11135
rect 5917 11101 5951 11135
rect 6184 11101 6218 11135
rect 7941 11101 7975 11135
rect 9965 11101 9999 11135
rect 13461 11101 13495 11135
rect 13645 11101 13679 11135
rect 16497 11101 16531 11135
rect 16681 11101 16715 11135
rect 17509 11101 17543 11135
rect 20269 11101 20303 11135
rect 23397 11101 23431 11135
rect 27537 11101 27571 11135
rect 28641 11101 28675 11135
rect 28825 11101 28859 11135
rect 28943 11101 28977 11135
rect 30481 11101 30515 11135
rect 30941 11101 30975 11135
rect 33333 11101 33367 11135
rect 33977 11101 34011 11135
rect 35081 11101 35115 11135
rect 36001 11101 36035 11135
rect 37197 11101 37231 11135
rect 37565 11101 37599 11135
rect 38209 11101 38243 11135
rect 39037 11101 39071 11135
rect 40233 11101 40267 11135
rect 44373 11101 44407 11135
rect 2320 11033 2354 11067
rect 4445 11033 4479 11067
rect 12357 11033 12391 11067
rect 27721 11033 27755 11067
rect 28733 11033 28767 11067
rect 35817 11033 35851 11067
rect 37381 11033 37415 11067
rect 37473 11033 37507 11067
rect 40049 11033 40083 11067
rect 41797 11033 41831 11067
rect 3985 10965 4019 10999
rect 9781 10965 9815 10999
rect 11161 10965 11195 10999
rect 12449 10965 12483 10999
rect 28457 10965 28491 10999
rect 33149 10965 33183 10999
rect 33793 10965 33827 10999
rect 35265 10965 35299 10999
rect 36185 10965 36219 10999
rect 2697 10761 2731 10795
rect 5733 10761 5767 10795
rect 10425 10761 10459 10795
rect 10793 10761 10827 10795
rect 11805 10761 11839 10795
rect 12173 10761 12207 10795
rect 14289 10761 14323 10795
rect 15393 10761 15427 10795
rect 18613 10761 18647 10795
rect 21097 10761 21131 10795
rect 25605 10761 25639 10795
rect 30941 10761 30975 10795
rect 37565 10761 37599 10795
rect 40065 10761 40099 10795
rect 42073 10761 42107 10795
rect 42625 10761 42659 10795
rect 3586 10693 3620 10727
rect 7849 10693 7883 10727
rect 25513 10693 25547 10727
rect 34713 10693 34747 10727
rect 39865 10693 39899 10727
rect 40960 10693 40994 10727
rect 2881 10625 2915 10659
rect 3341 10625 3375 10659
rect 5365 10625 5399 10659
rect 5549 10625 5583 10659
rect 12265 10625 12299 10659
rect 13001 10625 13035 10659
rect 15577 10625 15611 10659
rect 16037 10625 16071 10659
rect 16865 10625 16899 10659
rect 20269 10625 20303 10659
rect 21189 10625 21223 10659
rect 22560 10625 22594 10659
rect 26341 10625 26375 10659
rect 29653 10625 29687 10659
rect 37473 10625 37507 10659
rect 37657 10625 37691 10659
rect 39405 10625 39439 10659
rect 40693 10625 40727 10659
rect 42809 10625 42843 10659
rect 10885 10557 10919 10591
rect 10977 10557 11011 10591
rect 12449 10557 12483 10591
rect 17141 10557 17175 10591
rect 21373 10557 21407 10591
rect 22293 10557 22327 10591
rect 27169 10557 27203 10591
rect 27445 10557 27479 10591
rect 29193 10557 29227 10591
rect 32505 10557 32539 10591
rect 32781 10557 32815 10591
rect 4721 10489 4755 10523
rect 16037 10489 16071 10523
rect 20085 10489 20119 10523
rect 36001 10489 36035 10523
rect 9137 10421 9171 10455
rect 20729 10421 20763 10455
rect 23673 10421 23707 10455
rect 26341 10421 26375 10455
rect 34253 10421 34287 10455
rect 39221 10421 39255 10455
rect 40049 10421 40083 10455
rect 40233 10421 40267 10455
rect 2881 10217 2915 10251
rect 3985 10217 4019 10251
rect 12127 10217 12161 10251
rect 16497 10217 16531 10251
rect 18705 10217 18739 10251
rect 22845 10217 22879 10251
rect 26157 10217 26191 10251
rect 26801 10217 26835 10251
rect 28273 10217 28307 10251
rect 30573 10217 30607 10251
rect 33609 10217 33643 10251
rect 38301 10217 38335 10251
rect 40049 10217 40083 10251
rect 42809 10217 42843 10251
rect 13093 10149 13127 10183
rect 31125 10149 31159 10183
rect 4629 10081 4663 10115
rect 10333 10081 10367 10115
rect 10701 10081 10735 10115
rect 17785 10081 17819 10115
rect 20545 10081 20579 10115
rect 23397 10081 23431 10115
rect 31769 10081 31803 10115
rect 32505 10081 32539 10115
rect 34897 10081 34931 10115
rect 35173 10081 35207 10115
rect 37197 10081 37231 10115
rect 37565 10081 37599 10115
rect 39129 10081 39163 10115
rect 40969 10081 41003 10115
rect 43085 10081 43119 10115
rect 3065 10013 3099 10047
rect 4353 10013 4387 10047
rect 6561 10013 6595 10047
rect 6828 10013 6862 10047
rect 13001 10013 13035 10047
rect 13185 10013 13219 10047
rect 14289 10013 14323 10047
rect 14381 10013 14415 10047
rect 15117 10013 15151 10047
rect 16681 10013 16715 10047
rect 17509 10013 17543 10047
rect 17601 10013 17635 10047
rect 18337 10013 18371 10047
rect 18521 10013 18555 10047
rect 19717 10013 19751 10047
rect 20913 10013 20947 10047
rect 23213 10013 23247 10047
rect 26341 10013 26375 10047
rect 26985 10013 27019 10047
rect 27721 10013 27755 10047
rect 27813 10013 27847 10047
rect 28457 10013 28491 10047
rect 29929 10013 29963 10047
rect 30481 10013 30515 10047
rect 30665 10013 30699 10047
rect 31309 10013 31343 10047
rect 31401 10013 31435 10047
rect 32413 10013 32447 10047
rect 33609 10013 33643 10047
rect 34345 10013 34379 10047
rect 37381 10013 37415 10047
rect 37657 10013 37691 10047
rect 38117 10013 38151 10047
rect 39313 10013 39347 10047
rect 40233 10013 40267 10047
rect 40417 10013 40451 10047
rect 40509 10013 40543 10047
rect 41225 10013 41259 10047
rect 42809 10013 42843 10047
rect 42901 10013 42935 10047
rect 31493 9945 31527 9979
rect 31611 9945 31645 9979
rect 4445 9877 4479 9911
rect 7941 9877 7975 9911
rect 14933 9877 14967 9911
rect 17141 9877 17175 9911
rect 19809 9877 19843 9911
rect 22339 9877 22373 9911
rect 23305 9877 23339 9911
rect 29745 9877 29779 9911
rect 34161 9877 34195 9911
rect 36645 9877 36679 9911
rect 39497 9877 39531 9911
rect 42349 9877 42383 9911
rect 13461 9673 13495 9707
rect 27169 9673 27203 9707
rect 40417 9673 40451 9707
rect 5733 9605 5767 9639
rect 6806 9605 6840 9639
rect 10793 9605 10827 9639
rect 32873 9605 32907 9639
rect 36001 9605 36035 9639
rect 37565 9605 37599 9639
rect 39405 9605 39439 9639
rect 2780 9537 2814 9571
rect 5641 9537 5675 9571
rect 14105 9537 14139 9571
rect 15189 9537 15223 9571
rect 17132 9537 17166 9571
rect 19533 9537 19567 9571
rect 20177 9537 20211 9571
rect 21097 9537 21131 9571
rect 21189 9537 21223 9571
rect 22201 9537 22235 9571
rect 25237 9537 25271 9571
rect 26433 9537 26467 9571
rect 27353 9537 27387 9571
rect 27997 9537 28031 9571
rect 28457 9537 28491 9571
rect 28641 9537 28675 9571
rect 29552 9537 29586 9571
rect 31125 9537 31159 9571
rect 31309 9537 31343 9571
rect 32597 9537 32631 9571
rect 33241 9537 33275 9571
rect 33425 9537 33459 9571
rect 34713 9537 34747 9571
rect 34897 9537 34931 9571
rect 35725 9537 35759 9571
rect 35817 9537 35851 9571
rect 36461 9537 36495 9571
rect 36737 9537 36771 9571
rect 36829 9537 36863 9571
rect 37473 9537 37507 9571
rect 39589 9537 39623 9571
rect 39681 9537 39715 9571
rect 41613 9537 41647 9571
rect 41705 9537 41739 9571
rect 42625 9537 42659 9571
rect 42809 9537 42843 9571
rect 2513 9469 2547 9503
rect 5825 9469 5859 9503
rect 6561 9469 6595 9503
rect 10885 9469 10919 9503
rect 10977 9469 11011 9503
rect 11713 9469 11747 9503
rect 11989 9469 12023 9503
rect 14933 9469 14967 9503
rect 16865 9469 16899 9503
rect 21373 9469 21407 9503
rect 23857 9469 23891 9503
rect 28825 9469 28859 9503
rect 29285 9469 29319 9503
rect 33333 9469 33367 9503
rect 35357 9469 35391 9503
rect 36553 9469 36587 9503
rect 40141 9469 40175 9503
rect 40509 9469 40543 9503
rect 40626 9469 40660 9503
rect 41889 9469 41923 9503
rect 3893 9401 3927 9435
rect 7941 9401 7975 9435
rect 16313 9401 16347 9435
rect 32413 9401 32447 9435
rect 34805 9401 34839 9435
rect 39405 9401 39439 9435
rect 41245 9401 41279 9435
rect 5273 9333 5307 9367
rect 10425 9333 10459 9367
rect 13921 9333 13955 9367
rect 18245 9333 18279 9367
rect 19349 9333 19383 9367
rect 20177 9333 20211 9367
rect 20729 9333 20763 9367
rect 25053 9333 25087 9367
rect 26525 9333 26559 9367
rect 27813 9333 27847 9367
rect 30665 9333 30699 9367
rect 31125 9333 31159 9367
rect 36921 9333 36955 9367
rect 40785 9333 40819 9367
rect 42717 9333 42751 9367
rect 12173 9129 12207 9163
rect 14289 9129 14323 9163
rect 17601 9129 17635 9163
rect 26341 9129 26375 9163
rect 29193 9129 29227 9163
rect 35173 9129 35207 9163
rect 40049 9129 40083 9163
rect 7573 9061 7607 9095
rect 12633 9061 12667 9095
rect 23305 9061 23339 9095
rect 32045 9061 32079 9095
rect 39221 9061 39255 9095
rect 13093 8993 13127 9027
rect 13277 8993 13311 9027
rect 20821 8993 20855 9027
rect 21097 8993 21131 9027
rect 23029 8993 23063 9027
rect 30757 8993 30791 9027
rect 31585 8993 31619 9027
rect 33885 8993 33919 9027
rect 35357 8993 35391 9027
rect 35449 8993 35483 9027
rect 5273 8925 5307 8959
rect 9965 8925 9999 8959
rect 10425 8925 10459 8959
rect 13001 8925 13035 8959
rect 14473 8925 14507 8959
rect 16221 8925 16255 8959
rect 18245 8925 18279 8959
rect 19717 8925 19751 8959
rect 20361 8925 20395 8959
rect 24593 8925 24627 8959
rect 26985 8925 27019 8959
rect 27261 8925 27295 8959
rect 27813 8925 27847 8959
rect 30573 8925 30607 8959
rect 31677 8925 31711 8959
rect 33977 8925 34011 8959
rect 35817 8925 35851 8959
rect 36277 8925 36311 8959
rect 38761 8925 38795 8959
rect 39497 8925 39531 8959
rect 40049 8925 40083 8959
rect 40233 8925 40267 8959
rect 40693 8925 40727 8959
rect 42533 8925 42567 8959
rect 7849 8857 7883 8891
rect 8125 8857 8159 8891
rect 10701 8857 10735 8891
rect 16466 8857 16500 8891
rect 24869 8857 24903 8891
rect 28080 8857 28114 8891
rect 39221 8857 39255 8891
rect 40938 8857 40972 8891
rect 42800 8857 42834 8891
rect 6561 8789 6595 8823
rect 8033 8789 8067 8823
rect 9781 8789 9815 8823
rect 18061 8789 18095 8823
rect 19533 8789 19567 8823
rect 20177 8789 20211 8823
rect 22569 8789 22603 8823
rect 23489 8789 23523 8823
rect 26801 8789 26835 8823
rect 27169 8789 27203 8823
rect 30205 8789 30239 8823
rect 30665 8789 30699 8823
rect 34345 8789 34379 8823
rect 35541 8789 35575 8823
rect 35725 8789 35759 8823
rect 36461 8789 36495 8823
rect 38577 8789 38611 8823
rect 39405 8789 39439 8823
rect 42073 8789 42107 8823
rect 43913 8789 43947 8823
rect 9781 8585 9815 8619
rect 10333 8585 10367 8619
rect 10977 8585 11011 8619
rect 13461 8585 13495 8619
rect 20637 8585 20671 8619
rect 21097 8585 21131 8619
rect 25421 8585 25455 8619
rect 31309 8585 31343 8619
rect 34989 8585 35023 8619
rect 35633 8585 35667 8619
rect 35817 8585 35851 8619
rect 39405 8585 39439 8619
rect 42901 8585 42935 8619
rect 44189 8585 44223 8619
rect 4252 8517 4286 8551
rect 6828 8517 6862 8551
rect 8646 8517 8680 8551
rect 11989 8517 12023 8551
rect 15577 8517 15611 8551
rect 26433 8517 26467 8551
rect 28089 8517 28123 8551
rect 31125 8517 31159 8551
rect 35541 8517 35575 8551
rect 36277 8517 36311 8551
rect 36493 8517 36527 8551
rect 40509 8517 40543 8551
rect 41797 8517 41831 8551
rect 41981 8517 42015 8551
rect 42993 8517 43027 8551
rect 2145 8449 2179 8483
rect 2412 8449 2446 8483
rect 3985 8449 4019 8483
rect 10517 8449 10551 8483
rect 11161 8449 11195 8483
rect 11713 8449 11747 8483
rect 15485 8449 15519 8483
rect 17233 8449 17267 8483
rect 17500 8449 17534 8483
rect 19809 8449 19843 8483
rect 21005 8449 21039 8483
rect 22468 8449 22502 8483
rect 25421 8449 25455 8483
rect 26157 8449 26191 8483
rect 27261 8449 27295 8483
rect 28641 8449 28675 8483
rect 31033 8449 31067 8483
rect 31401 8449 31435 8483
rect 34621 8449 34655 8483
rect 35449 8449 35483 8483
rect 35817 8449 35851 8483
rect 38577 8449 38611 8483
rect 39681 8449 39715 8483
rect 39773 8449 39807 8483
rect 39865 8449 39899 8483
rect 40049 8449 40083 8483
rect 40969 8449 41003 8483
rect 41613 8449 41647 8483
rect 42809 8449 42843 8483
rect 44373 8449 44407 8483
rect 6561 8381 6595 8415
rect 8401 8381 8435 8415
rect 15669 8381 15703 8415
rect 19901 8381 19935 8415
rect 20085 8381 20119 8415
rect 21189 8381 21223 8415
rect 22201 8381 22235 8415
rect 31217 8381 31251 8415
rect 34529 8381 34563 8415
rect 40877 8381 40911 8415
rect 3525 8313 3559 8347
rect 7941 8313 7975 8347
rect 15117 8313 15151 8347
rect 19441 8313 19475 8347
rect 23581 8313 23615 8347
rect 29929 8313 29963 8347
rect 36645 8313 36679 8347
rect 41153 8313 41187 8347
rect 42625 8313 42659 8347
rect 5365 8245 5399 8279
rect 18613 8245 18647 8279
rect 36461 8245 36495 8279
rect 38669 8245 38703 8279
rect 40601 8245 40635 8279
rect 43177 8245 43211 8279
rect 6561 8041 6595 8075
rect 9781 8041 9815 8075
rect 16221 8041 16255 8075
rect 17785 8041 17819 8075
rect 22569 8041 22603 8075
rect 28641 8041 28675 8075
rect 32321 8041 32355 8075
rect 32505 8041 32539 8075
rect 34253 8041 34287 8075
rect 36553 8041 36587 8075
rect 37013 8041 37047 8075
rect 37381 8041 37415 8075
rect 41889 8041 41923 8075
rect 42349 8041 42383 8075
rect 1593 7973 1627 8007
rect 11897 7973 11931 8007
rect 31677 7973 31711 8007
rect 3157 7905 3191 7939
rect 3341 7905 3375 7939
rect 8309 7905 8343 7939
rect 8401 7905 8435 7939
rect 13093 7905 13127 7939
rect 18337 7905 18371 7939
rect 19901 7905 19935 7939
rect 26249 7905 26283 7939
rect 28089 7905 28123 7939
rect 34345 7905 34379 7939
rect 40509 7905 40543 7939
rect 1777 7837 1811 7871
rect 5273 7837 5307 7871
rect 9689 7837 9723 7871
rect 10517 7837 10551 7871
rect 12817 7837 12851 7871
rect 14841 7837 14875 7871
rect 16865 7837 16899 7871
rect 18153 7837 18187 7871
rect 20157 7837 20191 7871
rect 21925 7837 21959 7871
rect 22753 7837 22787 7871
rect 23489 7837 23523 7871
rect 25789 7837 25823 7871
rect 26617 7837 26651 7871
rect 28641 7837 28675 7871
rect 30297 7837 30331 7871
rect 34069 7837 34103 7871
rect 34161 7837 34195 7871
rect 35173 7837 35207 7871
rect 37013 7837 37047 7871
rect 37105 7837 37139 7871
rect 38025 7837 38059 7871
rect 39129 7837 39163 7871
rect 39221 7837 39255 7871
rect 39313 7837 39347 7871
rect 39497 7837 39531 7871
rect 42533 7837 42567 7871
rect 44373 7837 44407 7871
rect 8217 7769 8251 7803
rect 10762 7769 10796 7803
rect 15108 7769 15142 7803
rect 18245 7769 18279 7803
rect 30564 7769 30598 7803
rect 32137 7769 32171 7803
rect 35440 7769 35474 7803
rect 40776 7769 40810 7803
rect 2697 7701 2731 7735
rect 3065 7701 3099 7735
rect 7849 7701 7883 7735
rect 12449 7701 12483 7735
rect 12909 7701 12943 7735
rect 16681 7701 16715 7735
rect 21281 7701 21315 7735
rect 21741 7701 21775 7735
rect 23305 7701 23339 7735
rect 25605 7701 25639 7735
rect 32347 7701 32381 7735
rect 37841 7701 37875 7735
rect 38853 7701 38887 7735
rect 44189 7701 44223 7735
rect 3893 7497 3927 7531
rect 5273 7497 5307 7531
rect 9137 7497 9171 7531
rect 11713 7497 11747 7531
rect 12449 7497 12483 7531
rect 31033 7497 31067 7531
rect 31401 7497 31435 7531
rect 37565 7497 37599 7531
rect 38409 7497 38443 7531
rect 38577 7497 38611 7531
rect 39221 7497 39255 7531
rect 39589 7497 39623 7531
rect 40693 7497 40727 7531
rect 41429 7497 41463 7531
rect 2605 7429 2639 7463
rect 20168 7429 20202 7463
rect 23388 7429 23422 7463
rect 31585 7429 31619 7463
rect 33425 7429 33459 7463
rect 38209 7429 38243 7463
rect 40325 7429 40359 7463
rect 33655 7395 33689 7429
rect 2145 7361 2179 7395
rect 5181 7361 5215 7395
rect 7297 7361 7331 7395
rect 7757 7361 7791 7395
rect 8013 7361 8047 7395
rect 9873 7361 9907 7395
rect 10977 7361 11011 7395
rect 11897 7361 11931 7395
rect 12357 7361 12391 7395
rect 13277 7361 13311 7395
rect 13533 7361 13567 7395
rect 15485 7361 15519 7395
rect 17233 7361 17267 7395
rect 19901 7361 19935 7395
rect 25973 7361 26007 7395
rect 29193 7361 29227 7395
rect 29653 7361 29687 7395
rect 30297 7361 30331 7395
rect 31217 7361 31251 7395
rect 31677 7361 31711 7395
rect 32597 7361 32631 7395
rect 32689 7361 32723 7395
rect 32781 7361 32815 7395
rect 32965 7361 32999 7395
rect 34529 7361 34563 7395
rect 35173 7361 35207 7395
rect 36001 7361 36035 7395
rect 37473 7361 37507 7395
rect 39865 7361 39899 7395
rect 40969 7361 41003 7395
rect 41613 7361 41647 7395
rect 42625 7361 42659 7395
rect 42809 7361 42843 7395
rect 5457 7293 5491 7327
rect 15577 7293 15611 7327
rect 15669 7293 15703 7327
rect 23121 7293 23155 7327
rect 26249 7293 26283 7327
rect 27169 7293 27203 7327
rect 27445 7293 27479 7327
rect 31309 7293 31343 7327
rect 35449 7293 35483 7327
rect 36277 7293 36311 7327
rect 36369 7293 36403 7327
rect 36486 7293 36520 7327
rect 39405 7293 39439 7327
rect 39497 7293 39531 7327
rect 39773 7293 39807 7327
rect 40509 7293 40543 7327
rect 40601 7293 40635 7327
rect 40877 7293 40911 7327
rect 4813 7225 4847 7259
rect 7113 7225 7147 7259
rect 21281 7225 21315 7259
rect 34989 7225 35023 7259
rect 35357 7225 35391 7259
rect 1961 7157 1995 7191
rect 9873 7157 9907 7191
rect 11069 7157 11103 7191
rect 14657 7157 14691 7191
rect 15117 7157 15151 7191
rect 17325 7157 17359 7191
rect 24501 7157 24535 7191
rect 29745 7157 29779 7191
rect 30389 7157 30423 7191
rect 32321 7157 32355 7191
rect 33609 7157 33643 7191
rect 33793 7157 33827 7191
rect 34345 7157 34379 7191
rect 36645 7157 36679 7191
rect 38393 7157 38427 7191
rect 42625 7157 42659 7191
rect 3433 6953 3467 6987
rect 9400 6953 9434 6987
rect 12357 6953 12391 6987
rect 31585 6953 31619 6987
rect 35725 6953 35759 6987
rect 13001 6885 13035 6919
rect 9137 6817 9171 6851
rect 13461 6817 13495 6851
rect 13645 6817 13679 6851
rect 15301 6817 15335 6851
rect 17693 6817 17727 6851
rect 18613 6817 18647 6851
rect 20545 6817 20579 6851
rect 23765 6817 23799 6851
rect 23857 6817 23891 6851
rect 24685 6817 24719 6851
rect 25145 6817 25179 6851
rect 31861 6817 31895 6851
rect 32229 6817 32263 6851
rect 43453 6817 43487 6851
rect 2053 6749 2087 6783
rect 3985 6749 4019 6783
rect 4252 6749 4286 6783
rect 6561 6749 6595 6783
rect 8309 6749 8343 6783
rect 11897 6749 11931 6783
rect 12541 6749 12575 6783
rect 13369 6749 13403 6783
rect 14473 6749 14507 6783
rect 18521 6749 18555 6783
rect 20177 6749 20211 6783
rect 20361 6749 20395 6783
rect 20456 6749 20490 6783
rect 20729 6749 20763 6783
rect 21373 6749 21407 6783
rect 21466 6749 21500 6783
rect 21649 6749 21683 6783
rect 21838 6749 21872 6783
rect 23673 6749 23707 6783
rect 24777 6749 24811 6783
rect 25973 6749 26007 6783
rect 26801 6749 26835 6783
rect 27261 6749 27295 6783
rect 29745 6749 29779 6783
rect 31769 6749 31803 6783
rect 32137 6749 32171 6783
rect 32689 6749 32723 6783
rect 33977 6749 34011 6783
rect 34161 6749 34195 6783
rect 35357 6749 35391 6783
rect 35725 6749 35759 6783
rect 36553 6749 36587 6783
rect 36737 6749 36771 6783
rect 36921 6749 36955 6783
rect 37381 6749 37415 6783
rect 39497 6749 39531 6783
rect 40233 6749 40267 6783
rect 40509 6749 40543 6783
rect 40693 6749 40727 6783
rect 41337 6749 41371 6783
rect 43361 6749 43395 6783
rect 2320 6681 2354 6715
rect 15568 6681 15602 6715
rect 17509 6681 17543 6715
rect 21741 6681 21775 6715
rect 28457 6681 28491 6715
rect 30012 6681 30046 6715
rect 36369 6681 36403 6715
rect 41582 6681 41616 6715
rect 5365 6613 5399 6647
rect 6377 6613 6411 6647
rect 8493 6613 8527 6647
rect 10885 6613 10919 6647
rect 11713 6613 11747 6647
rect 14289 6613 14323 6647
rect 16681 6613 16715 6647
rect 17141 6613 17175 6647
rect 17601 6613 17635 6647
rect 18889 6613 18923 6647
rect 20913 6613 20947 6647
rect 22017 6613 22051 6647
rect 23305 6613 23339 6647
rect 25789 6613 25823 6647
rect 26617 6613 26651 6647
rect 31125 6613 31159 6647
rect 32045 6613 32079 6647
rect 32781 6613 32815 6647
rect 34345 6613 34379 6647
rect 35909 6613 35943 6647
rect 36645 6613 36679 6647
rect 37473 6613 37507 6647
rect 39313 6613 39347 6647
rect 40049 6613 40083 6647
rect 42717 6613 42751 6647
rect 43729 6613 43763 6647
rect 3433 6409 3467 6443
rect 5365 6409 5399 6443
rect 10333 6409 10367 6443
rect 10793 6409 10827 6443
rect 15577 6409 15611 6443
rect 17969 6409 18003 6443
rect 23213 6409 23247 6443
rect 27261 6409 27295 6443
rect 30481 6409 30515 6443
rect 31125 6409 31159 6443
rect 4252 6341 4286 6375
rect 9873 6341 9907 6375
rect 13001 6341 13035 6375
rect 14749 6341 14783 6375
rect 23765 6341 23799 6375
rect 23981 6341 24015 6375
rect 33333 6341 33367 6375
rect 34253 6341 34287 6375
rect 40877 6341 40911 6375
rect 41337 6341 41371 6375
rect 2053 6273 2087 6307
rect 2320 6273 2354 6307
rect 6009 6273 6043 6307
rect 8493 6273 8527 6307
rect 9137 6273 9171 6307
rect 10977 6273 11011 6307
rect 15761 6273 15795 6307
rect 17966 6273 18000 6307
rect 19165 6273 19199 6307
rect 19257 6273 19291 6307
rect 19349 6273 19383 6307
rect 19533 6273 19567 6307
rect 19993 6273 20027 6307
rect 20453 6273 20487 6307
rect 23121 6273 23155 6307
rect 27169 6273 27203 6307
rect 27353 6273 27387 6307
rect 28641 6273 28675 6307
rect 29285 6273 29319 6307
rect 29745 6273 29779 6307
rect 30665 6273 30699 6307
rect 31309 6273 31343 6307
rect 33241 6273 33275 6307
rect 33885 6273 33919 6307
rect 33977 6273 34011 6307
rect 34161 6273 34195 6307
rect 34345 6273 34379 6307
rect 35449 6273 35483 6307
rect 35633 6273 35667 6307
rect 35725 6273 35759 6307
rect 36645 6273 36679 6307
rect 37473 6273 37507 6307
rect 37657 6273 37691 6307
rect 38485 6273 38519 6307
rect 38669 6273 38703 6307
rect 39037 6273 39071 6307
rect 40601 6273 40635 6307
rect 41521 6273 41555 6307
rect 41613 6273 41647 6307
rect 42809 6273 42843 6307
rect 3985 6205 4019 6239
rect 8953 6205 8987 6239
rect 18429 6205 18463 6239
rect 20177 6205 20211 6239
rect 20821 6205 20855 6239
rect 24593 6205 24627 6239
rect 24869 6205 24903 6239
rect 30021 6205 30055 6239
rect 35265 6205 35299 6239
rect 36461 6205 36495 6239
rect 36553 6205 36587 6239
rect 38761 6205 38795 6239
rect 38853 6205 38887 6239
rect 40693 6205 40727 6239
rect 40877 6205 40911 6239
rect 41409 6205 41443 6239
rect 5825 6137 5859 6171
rect 10241 6137 10275 6171
rect 17785 6137 17819 6171
rect 20085 6137 20119 6171
rect 35541 6137 35575 6171
rect 8309 6069 8343 6103
rect 9321 6069 9355 6103
rect 18337 6069 18371 6103
rect 18889 6069 18923 6103
rect 23949 6069 23983 6103
rect 24133 6069 24167 6103
rect 26341 6069 26375 6103
rect 28457 6069 28491 6103
rect 29101 6069 29135 6103
rect 29837 6069 29871 6103
rect 29929 6069 29963 6103
rect 33885 6069 33919 6103
rect 36277 6069 36311 6103
rect 37473 6069 37507 6103
rect 39221 6069 39255 6103
rect 42625 6069 42659 6103
rect 1777 5865 1811 5899
rect 5365 5865 5399 5899
rect 11713 5865 11747 5899
rect 15669 5865 15703 5899
rect 17785 5865 17819 5899
rect 18337 5865 18371 5899
rect 19993 5865 20027 5899
rect 20913 5865 20947 5899
rect 23029 5865 23063 5899
rect 23857 5865 23891 5899
rect 24593 5865 24627 5899
rect 26065 5865 26099 5899
rect 27629 5865 27663 5899
rect 28641 5865 28675 5899
rect 34161 5865 34195 5899
rect 34345 5865 34379 5899
rect 36277 5865 36311 5899
rect 36921 5865 36955 5899
rect 18797 5797 18831 5831
rect 24041 5797 24075 5831
rect 8585 5729 8619 5763
rect 13737 5729 13771 5763
rect 30297 5729 30331 5763
rect 32965 5729 32999 5763
rect 34897 5729 34931 5763
rect 40785 5729 40819 5763
rect 2973 5661 3007 5695
rect 3985 5661 4019 5695
rect 5825 5661 5859 5695
rect 6009 5661 6043 5695
rect 7573 5661 7607 5695
rect 8217 5661 8251 5695
rect 8401 5661 8435 5695
rect 10425 5661 10459 5695
rect 12633 5661 12667 5695
rect 13461 5661 13495 5695
rect 13553 5661 13587 5695
rect 14289 5661 14323 5695
rect 16313 5661 16347 5695
rect 17693 5661 17727 5695
rect 18521 5661 18555 5695
rect 18613 5661 18647 5695
rect 18889 5661 18923 5695
rect 19441 5661 19475 5695
rect 19717 5661 19751 5695
rect 19809 5661 19843 5695
rect 20545 5661 20579 5695
rect 20637 5661 20671 5695
rect 20729 5661 20763 5695
rect 21373 5661 21407 5695
rect 22385 5661 22419 5695
rect 23213 5661 23247 5695
rect 24777 5661 24811 5695
rect 25053 5661 25087 5695
rect 25881 5661 25915 5695
rect 27537 5661 27571 5695
rect 28641 5661 28675 5695
rect 28917 5661 28951 5695
rect 30389 5661 30423 5695
rect 31217 5661 31251 5695
rect 34069 5661 34103 5695
rect 34253 5661 34287 5695
rect 35153 5661 35187 5695
rect 38025 5661 38059 5695
rect 38118 5661 38152 5695
rect 38393 5661 38427 5695
rect 38531 5661 38565 5695
rect 41052 5661 41086 5695
rect 4230 5593 4264 5627
rect 7941 5593 7975 5627
rect 14556 5593 14590 5627
rect 19625 5593 19659 5627
rect 21465 5593 21499 5627
rect 23673 5593 23707 5627
rect 23889 5593 23923 5627
rect 33885 5593 33919 5627
rect 36737 5593 36771 5627
rect 36937 5593 36971 5627
rect 38301 5593 38335 5627
rect 2789 5525 2823 5559
rect 6193 5525 6227 5559
rect 7389 5525 7423 5559
rect 12725 5525 12759 5559
rect 13737 5525 13771 5559
rect 16129 5525 16163 5559
rect 22477 5525 22511 5559
rect 24961 5525 24995 5559
rect 28825 5525 28859 5559
rect 30757 5525 30791 5559
rect 37105 5525 37139 5559
rect 38669 5525 38703 5559
rect 42165 5525 42199 5559
rect 4353 5321 4387 5355
rect 4445 5321 4479 5355
rect 10885 5321 10919 5355
rect 13001 5321 13035 5355
rect 16037 5321 16071 5355
rect 17167 5321 17201 5355
rect 17785 5321 17819 5355
rect 22753 5321 22787 5355
rect 41705 5321 41739 5355
rect 7205 5253 7239 5287
rect 12817 5253 12851 5287
rect 16957 5253 16991 5287
rect 18797 5253 18831 5287
rect 19013 5253 19047 5287
rect 19809 5253 19843 5287
rect 26525 5253 26559 5287
rect 37565 5253 37599 5287
rect 38786 5253 38820 5287
rect 5181 5185 5215 5219
rect 5365 5185 5399 5219
rect 6929 5185 6963 5219
rect 9137 5185 9171 5219
rect 12357 5185 12391 5219
rect 13093 5185 13127 5219
rect 13553 5185 13587 5219
rect 15761 5185 15795 5219
rect 18061 5185 18095 5219
rect 18153 5185 18187 5219
rect 18245 5185 18279 5219
rect 19993 5185 20027 5219
rect 20637 5185 20671 5219
rect 20821 5185 20855 5219
rect 21281 5185 21315 5219
rect 21465 5185 21499 5219
rect 22661 5185 22695 5219
rect 23305 5185 23339 5219
rect 23489 5185 23523 5219
rect 23949 5185 23983 5219
rect 24041 5185 24075 5219
rect 24225 5185 24259 5219
rect 24317 5185 24351 5219
rect 24409 5185 24443 5219
rect 24961 5185 24995 5219
rect 25237 5185 25271 5219
rect 25329 5185 25363 5219
rect 25973 5185 26007 5219
rect 26433 5185 26467 5219
rect 33149 5185 33183 5219
rect 33609 5185 33643 5219
rect 33865 5185 33899 5219
rect 35449 5185 35483 5219
rect 35705 5185 35739 5219
rect 37473 5185 37507 5219
rect 38301 5185 38335 5219
rect 41705 5185 41739 5219
rect 42809 5185 42843 5219
rect 1593 5117 1627 5151
rect 1869 5117 1903 5151
rect 4629 5117 4663 5151
rect 8677 5117 8711 5151
rect 9413 5117 9447 5151
rect 13829 5117 13863 5151
rect 15301 5117 15335 5151
rect 15853 5117 15887 5151
rect 16037 5109 16071 5143
rect 17969 5117 18003 5151
rect 24501 5117 24535 5151
rect 28089 5117 28123 5151
rect 28365 5117 28399 5151
rect 29837 5117 29871 5151
rect 38577 5117 38611 5151
rect 38669 5117 38703 5151
rect 44005 5117 44039 5151
rect 3985 5049 4019 5083
rect 20637 5049 20671 5083
rect 32965 5049 32999 5083
rect 38945 5049 38979 5083
rect 5549 4981 5583 5015
rect 12173 4981 12207 5015
rect 12817 4981 12851 5015
rect 17141 4981 17175 5015
rect 17325 4981 17359 5015
rect 18981 4981 19015 5015
rect 19165 4981 19199 5015
rect 20177 4981 20211 5015
rect 21373 4981 21407 5015
rect 23305 4981 23339 5015
rect 25789 4981 25823 5015
rect 34989 4981 35023 5015
rect 36829 4981 36863 5015
rect 10425 4777 10459 4811
rect 14473 4777 14507 4811
rect 18889 4777 18923 4811
rect 21189 4777 21223 4811
rect 27353 4777 27387 4811
rect 34897 4777 34931 4811
rect 37105 4777 37139 4811
rect 38301 4777 38335 4811
rect 13553 4709 13587 4743
rect 21649 4709 21683 4743
rect 23949 4709 23983 4743
rect 11805 4641 11839 4675
rect 12081 4641 12115 4675
rect 17141 4641 17175 4675
rect 19441 4641 19475 4675
rect 19717 4641 19751 4675
rect 25605 4641 25639 4675
rect 36829 4641 36863 4675
rect 38117 4641 38151 4675
rect 4721 4573 4755 4607
rect 4813 4573 4847 4607
rect 9873 4573 9907 4607
rect 9965 4573 9999 4607
rect 10609 4573 10643 4607
rect 14473 4573 14507 4607
rect 15025 4573 15059 4607
rect 15209 4573 15243 4607
rect 21833 4573 21867 4607
rect 23765 4573 23799 4607
rect 24041 4573 24075 4607
rect 24593 4573 24627 4607
rect 24777 4573 24811 4607
rect 25053 4573 25087 4607
rect 29929 4573 29963 4607
rect 30573 4573 30607 4607
rect 35081 4573 35115 4607
rect 36737 4573 36771 4607
rect 38025 4573 38059 4607
rect 17417 4505 17451 4539
rect 25881 4505 25915 4539
rect 4997 4437 5031 4471
rect 15117 4437 15151 4471
rect 23581 4437 23615 4471
rect 24961 4437 24995 4471
rect 29745 4437 29779 4471
rect 30389 4437 30423 4471
rect 12725 4233 12759 4267
rect 14105 4233 14139 4267
rect 17693 4233 17727 4267
rect 18613 4233 18647 4267
rect 20198 4233 20232 4267
rect 25421 4233 25455 4267
rect 25881 4233 25915 4267
rect 19993 4165 20027 4199
rect 9413 4097 9447 4131
rect 12909 4097 12943 4131
rect 14289 4097 14323 4131
rect 16313 4097 16347 4131
rect 16957 4097 16991 4131
rect 17877 4097 17911 4131
rect 18613 4097 18647 4131
rect 19165 4097 19199 4131
rect 21005 4097 21039 4131
rect 23673 4097 23707 4131
rect 26065 4097 26099 4131
rect 27169 4097 27203 4131
rect 28365 4097 28399 4131
rect 28457 4097 28491 4131
rect 29377 4097 29411 4131
rect 31401 4097 31435 4131
rect 23949 4029 23983 4063
rect 29653 4029 29687 4063
rect 9229 3961 9263 3995
rect 16957 3961 16991 3995
rect 20361 3961 20395 3995
rect 16129 3893 16163 3927
rect 19257 3893 19291 3927
rect 20177 3893 20211 3927
rect 20821 3893 20855 3927
rect 27169 3893 27203 3927
rect 19441 3689 19475 3723
rect 20453 3689 20487 3723
rect 23857 3689 23891 3723
rect 24869 3689 24903 3723
rect 26801 3689 26835 3723
rect 30297 3621 30331 3655
rect 6285 3553 6319 3587
rect 30021 3553 30055 3587
rect 1777 3485 1811 3519
rect 5641 3485 5675 3519
rect 13553 3485 13587 3519
rect 14749 3485 14783 3519
rect 15393 3485 15427 3519
rect 15853 3485 15887 3519
rect 16221 3485 16255 3519
rect 18153 3485 18187 3519
rect 19625 3485 19659 3519
rect 20637 3485 20671 3519
rect 24041 3485 24075 3519
rect 24777 3485 24811 3519
rect 26985 3485 27019 3519
rect 29929 3485 29963 3519
rect 44373 3485 44407 3519
rect 17647 3417 17681 3451
rect 13645 3349 13679 3383
rect 15209 3349 15243 3383
rect 18245 3349 18279 3383
rect 17049 3145 17083 3179
rect 44189 3145 44223 3179
rect 19809 3077 19843 3111
rect 7205 3009 7239 3043
rect 13645 3009 13679 3043
rect 14841 3009 14875 3043
rect 16267 3009 16301 3043
rect 16865 3009 16899 3043
rect 18061 3009 18095 3043
rect 20453 3009 20487 3043
rect 22937 3009 22971 3043
rect 34253 3009 34287 3043
rect 44373 3009 44407 3043
rect 8401 2941 8435 2975
rect 14473 2941 14507 2975
rect 17693 2941 17727 2975
rect 23397 2941 23431 2975
rect 35449 2941 35483 2975
rect 13829 2873 13863 2907
rect 20269 2873 20303 2907
rect 1777 2805 1811 2839
rect 12909 2601 12943 2635
rect 14841 2601 14875 2635
rect 16221 2601 16255 2635
rect 27537 2601 27571 2635
rect 32505 2601 32539 2635
rect 37473 2601 37507 2635
rect 43913 2601 43947 2635
rect 13737 2533 13771 2567
rect 16957 2533 16991 2567
rect 2421 2465 2455 2499
rect 42901 2465 42935 2499
rect 1777 2397 1811 2431
rect 4169 2397 4203 2431
rect 4813 2397 4847 2431
rect 8033 2397 8067 2431
rect 11897 2397 11931 2431
rect 13093 2397 13127 2431
rect 14749 2397 14783 2431
rect 15393 2397 15427 2431
rect 15485 2397 15519 2431
rect 16037 2397 16071 2431
rect 16865 2397 16899 2431
rect 17509 2397 17543 2431
rect 17785 2397 17819 2431
rect 19625 2397 19659 2431
rect 20913 2397 20947 2431
rect 24777 2397 24811 2431
rect 26065 2397 26099 2431
rect 29929 2397 29963 2431
rect 30573 2397 30607 2431
rect 37657 2397 37691 2431
rect 38945 2397 38979 2431
rect 40233 2397 40267 2431
rect 44097 2397 44131 2431
rect 27261 2329 27295 2363
rect 32413 2329 32447 2363
rect 42717 2329 42751 2363
rect 25881 2261 25915 2295
<< metal1 >>
rect 16114 19048 16120 19100
rect 16172 19088 16178 19100
rect 16850 19088 16856 19100
rect 16172 19060 16856 19088
rect 16172 19048 16178 19060
rect 16850 19048 16856 19060
rect 16908 19048 16914 19100
rect 34146 19048 34152 19100
rect 34204 19088 34210 19100
rect 35066 19088 35072 19100
rect 34204 19060 35072 19088
rect 34204 19048 34210 19060
rect 35066 19048 35072 19060
rect 35124 19048 35130 19100
rect 41874 19048 41880 19100
rect 41932 19088 41938 19100
rect 42794 19088 42800 19100
rect 41932 19060 42800 19088
rect 41932 19048 41938 19060
rect 42794 19048 42800 19060
rect 42852 19048 42858 19100
rect 43438 18028 43444 18080
rect 43496 18068 43502 18080
rect 45002 18068 45008 18080
rect 43496 18040 45008 18068
rect 43496 18028 43502 18040
rect 45002 18028 45008 18040
rect 45060 18028 45066 18080
rect 43990 17484 43996 17536
rect 44048 17524 44054 17536
rect 45002 17524 45008 17536
rect 44048 17496 45008 17524
rect 44048 17484 44054 17496
rect 45002 17484 45008 17496
rect 45060 17484 45066 17536
rect 1104 17434 45051 17456
rect 1104 17382 11896 17434
rect 11948 17382 11960 17434
rect 12012 17382 12024 17434
rect 12076 17382 12088 17434
rect 12140 17382 12152 17434
rect 12204 17382 22843 17434
rect 22895 17382 22907 17434
rect 22959 17382 22971 17434
rect 23023 17382 23035 17434
rect 23087 17382 23099 17434
rect 23151 17382 33790 17434
rect 33842 17382 33854 17434
rect 33906 17382 33918 17434
rect 33970 17382 33982 17434
rect 34034 17382 34046 17434
rect 34098 17382 44737 17434
rect 44789 17382 44801 17434
rect 44853 17382 44865 17434
rect 44917 17382 44929 17434
rect 44981 17382 44993 17434
rect 45045 17382 45051 17434
rect 1104 17360 45051 17382
rect 934 17212 940 17264
rect 992 17252 998 17264
rect 2409 17255 2467 17261
rect 2409 17252 2421 17255
rect 992 17224 2421 17252
rect 992 17212 998 17224
rect 2409 17221 2421 17224
rect 2455 17221 2467 17255
rect 2409 17215 2467 17221
rect 3234 17212 3240 17264
rect 3292 17212 3298 17264
rect 11054 17212 11060 17264
rect 11112 17252 11118 17264
rect 11793 17255 11851 17261
rect 11793 17252 11805 17255
rect 11112 17224 11805 17252
rect 11112 17212 11118 17224
rect 11793 17221 11805 17224
rect 11839 17221 11851 17255
rect 11793 17215 11851 17221
rect 38654 17212 38660 17264
rect 38712 17252 38718 17264
rect 38841 17255 38899 17261
rect 38841 17252 38853 17255
rect 38712 17224 38853 17252
rect 38712 17212 38718 17224
rect 38841 17221 38853 17224
rect 38887 17221 38899 17255
rect 38841 17215 38899 17221
rect 1302 17144 1308 17196
rect 1360 17184 1366 17196
rect 1581 17187 1639 17193
rect 1581 17184 1593 17187
rect 1360 17156 1593 17184
rect 1360 17144 1366 17156
rect 1581 17153 1593 17156
rect 1627 17153 1639 17187
rect 1581 17147 1639 17153
rect 4522 17144 4528 17196
rect 4580 17184 4586 17196
rect 4617 17187 4675 17193
rect 4617 17184 4629 17187
rect 4580 17156 4629 17184
rect 4580 17144 4586 17156
rect 4617 17153 4629 17156
rect 4663 17153 4675 17187
rect 4617 17147 4675 17153
rect 6454 17144 6460 17196
rect 6512 17184 6518 17196
rect 6733 17187 6791 17193
rect 6733 17184 6745 17187
rect 6512 17156 6745 17184
rect 6512 17144 6518 17156
rect 6733 17153 6745 17156
rect 6779 17153 6791 17187
rect 6733 17147 6791 17153
rect 7742 17144 7748 17196
rect 7800 17184 7806 17196
rect 8021 17187 8079 17193
rect 8021 17184 8033 17187
rect 7800 17156 8033 17184
rect 7800 17144 7806 17156
rect 8021 17153 8033 17156
rect 8067 17153 8079 17187
rect 8021 17147 8079 17153
rect 9674 17144 9680 17196
rect 9732 17184 9738 17196
rect 9953 17187 10011 17193
rect 9953 17184 9965 17187
rect 9732 17156 9965 17184
rect 9732 17144 9738 17156
rect 9953 17153 9965 17156
rect 9999 17153 10011 17187
rect 9953 17147 10011 17153
rect 12894 17144 12900 17196
rect 12952 17184 12958 17196
rect 13173 17187 13231 17193
rect 13173 17184 13185 17187
rect 12952 17156 13185 17184
rect 12952 17144 12958 17156
rect 13173 17153 13185 17156
rect 13219 17153 13231 17187
rect 13173 17147 13231 17153
rect 14182 17144 14188 17196
rect 14240 17184 14246 17196
rect 14461 17187 14519 17193
rect 14461 17184 14473 17187
rect 14240 17156 14473 17184
rect 14240 17144 14246 17156
rect 14461 17153 14473 17156
rect 14507 17153 14519 17187
rect 14461 17147 14519 17153
rect 16850 17144 16856 17196
rect 16908 17144 16914 17196
rect 19334 17144 19340 17196
rect 19392 17184 19398 17196
rect 19613 17187 19671 17193
rect 19613 17184 19625 17187
rect 19392 17156 19625 17184
rect 19392 17144 19398 17156
rect 19613 17153 19625 17156
rect 19659 17153 19671 17187
rect 19613 17147 19671 17153
rect 22554 17144 22560 17196
rect 22612 17184 22618 17196
rect 22833 17187 22891 17193
rect 22833 17184 22845 17187
rect 22612 17156 22845 17184
rect 22612 17144 22618 17156
rect 22833 17153 22845 17156
rect 22879 17153 22891 17187
rect 22833 17147 22891 17153
rect 23842 17144 23848 17196
rect 23900 17184 23906 17196
rect 24765 17187 24823 17193
rect 24765 17184 24777 17187
rect 23900 17156 24777 17184
rect 23900 17144 23906 17156
rect 24765 17153 24777 17156
rect 24811 17153 24823 17187
rect 24765 17147 24823 17153
rect 25774 17144 25780 17196
rect 25832 17184 25838 17196
rect 26053 17187 26111 17193
rect 26053 17184 26065 17187
rect 25832 17156 26065 17184
rect 25832 17144 25838 17156
rect 26053 17153 26065 17156
rect 26099 17153 26111 17187
rect 26053 17147 26111 17153
rect 27706 17144 27712 17196
rect 27764 17184 27770 17196
rect 27985 17187 28043 17193
rect 27985 17184 27997 17187
rect 27764 17156 27997 17184
rect 27764 17144 27770 17156
rect 27985 17153 27997 17156
rect 28031 17153 28043 17187
rect 27985 17147 28043 17153
rect 28994 17144 29000 17196
rect 29052 17184 29058 17196
rect 29917 17187 29975 17193
rect 29917 17184 29929 17187
rect 29052 17156 29929 17184
rect 29052 17144 29058 17156
rect 29917 17153 29929 17156
rect 29963 17153 29975 17187
rect 29917 17147 29975 17153
rect 30926 17144 30932 17196
rect 30984 17184 30990 17196
rect 31205 17187 31263 17193
rect 31205 17184 31217 17187
rect 30984 17156 31217 17184
rect 30984 17144 30990 17156
rect 31205 17153 31217 17156
rect 31251 17153 31263 17187
rect 31205 17147 31263 17153
rect 32214 17144 32220 17196
rect 32272 17184 32278 17196
rect 32309 17187 32367 17193
rect 32309 17184 32321 17187
rect 32272 17156 32321 17184
rect 32272 17144 32278 17156
rect 32309 17153 32321 17156
rect 32355 17153 32367 17187
rect 32309 17147 32367 17153
rect 35066 17144 35072 17196
rect 35124 17144 35130 17196
rect 35434 17144 35440 17196
rect 35492 17184 35498 17196
rect 35713 17187 35771 17193
rect 35713 17184 35725 17187
rect 35492 17156 35725 17184
rect 35492 17144 35498 17156
rect 35713 17153 35725 17156
rect 35759 17153 35771 17187
rect 35713 17147 35771 17153
rect 37366 17144 37372 17196
rect 37424 17184 37430 17196
rect 37645 17187 37703 17193
rect 37645 17184 37657 17187
rect 37424 17156 37657 17184
rect 37424 17144 37430 17156
rect 37645 17153 37657 17156
rect 37691 17153 37703 17187
rect 37645 17147 37703 17153
rect 42794 17144 42800 17196
rect 42852 17144 42858 17196
rect 43438 17144 43444 17196
rect 43496 17144 43502 17196
rect 43806 17144 43812 17196
rect 43864 17184 43870 17196
rect 44085 17187 44143 17193
rect 44085 17184 44097 17187
rect 43864 17156 44097 17184
rect 43864 17144 43870 17156
rect 44085 17153 44097 17156
rect 44131 17153 44143 17187
rect 44085 17147 44143 17153
rect 4893 17119 4951 17125
rect 4893 17085 4905 17119
rect 4939 17116 4951 17119
rect 10870 17116 10876 17128
rect 4939 17088 10876 17116
rect 4939 17085 4951 17088
rect 4893 17079 4951 17085
rect 10870 17076 10876 17088
rect 10928 17076 10934 17128
rect 32582 17076 32588 17128
rect 32640 17076 32646 17128
rect 3421 17051 3479 17057
rect 3421 17017 3433 17051
rect 3467 17048 3479 17051
rect 3602 17048 3608 17060
rect 3467 17020 3608 17048
rect 3467 17017 3479 17020
rect 3421 17011 3479 17017
rect 3602 17008 3608 17020
rect 3660 17008 3666 17060
rect 11977 17051 12035 17057
rect 11977 17017 11989 17051
rect 12023 17048 12035 17051
rect 15654 17048 15660 17060
rect 12023 17020 15660 17048
rect 12023 17017 12035 17020
rect 11977 17011 12035 17017
rect 15654 17008 15660 17020
rect 15712 17008 15718 17060
rect 1762 16940 1768 16992
rect 1820 16940 1826 16992
rect 2498 16940 2504 16992
rect 2556 16940 2562 16992
rect 9769 16983 9827 16989
rect 9769 16949 9781 16983
rect 9815 16980 9827 16983
rect 10226 16980 10232 16992
rect 9815 16952 10232 16980
rect 9815 16949 9827 16952
rect 9769 16943 9827 16949
rect 10226 16940 10232 16952
rect 10284 16940 10290 16992
rect 16574 16940 16580 16992
rect 16632 16980 16638 16992
rect 17037 16983 17095 16989
rect 17037 16980 17049 16983
rect 16632 16952 17049 16980
rect 16632 16940 16638 16952
rect 17037 16949 17049 16952
rect 17083 16949 17095 16983
rect 17037 16943 17095 16949
rect 23750 16940 23756 16992
rect 23808 16980 23814 16992
rect 24581 16983 24639 16989
rect 24581 16980 24593 16983
rect 23808 16952 24593 16980
rect 23808 16940 23814 16952
rect 24581 16949 24593 16952
rect 24627 16949 24639 16983
rect 24581 16943 24639 16949
rect 31021 16983 31079 16989
rect 31021 16949 31033 16983
rect 31067 16980 31079 16983
rect 31294 16980 31300 16992
rect 31067 16952 31300 16980
rect 31067 16949 31079 16952
rect 31021 16943 31079 16949
rect 31294 16940 31300 16952
rect 31352 16940 31358 16992
rect 34514 16940 34520 16992
rect 34572 16980 34578 16992
rect 34885 16983 34943 16989
rect 34885 16980 34897 16983
rect 34572 16952 34897 16980
rect 34572 16940 34578 16952
rect 34885 16949 34897 16952
rect 34931 16949 34943 16983
rect 34885 16943 34943 16949
rect 38838 16940 38844 16992
rect 38896 16980 38902 16992
rect 38933 16983 38991 16989
rect 38933 16980 38945 16983
rect 38896 16952 38945 16980
rect 38896 16940 38902 16952
rect 38933 16949 38945 16952
rect 38979 16949 38991 16983
rect 38933 16943 38991 16949
rect 1104 16890 44896 16912
rect 1104 16838 6423 16890
rect 6475 16838 6487 16890
rect 6539 16838 6551 16890
rect 6603 16838 6615 16890
rect 6667 16838 6679 16890
rect 6731 16838 17370 16890
rect 17422 16838 17434 16890
rect 17486 16838 17498 16890
rect 17550 16838 17562 16890
rect 17614 16838 17626 16890
rect 17678 16838 28317 16890
rect 28369 16838 28381 16890
rect 28433 16838 28445 16890
rect 28497 16838 28509 16890
rect 28561 16838 28573 16890
rect 28625 16838 39264 16890
rect 39316 16838 39328 16890
rect 39380 16838 39392 16890
rect 39444 16838 39456 16890
rect 39508 16838 39520 16890
rect 39572 16838 44896 16890
rect 1104 16816 44896 16838
rect 44361 16779 44419 16785
rect 44361 16745 44373 16779
rect 44407 16776 44419 16779
rect 45094 16776 45100 16788
rect 44407 16748 45100 16776
rect 44407 16745 44419 16748
rect 44361 16739 44419 16745
rect 45094 16736 45100 16748
rect 45152 16736 45158 16788
rect 1857 16643 1915 16649
rect 1857 16609 1869 16643
rect 1903 16640 1915 16643
rect 5166 16640 5172 16652
rect 1903 16612 5172 16640
rect 1903 16609 1915 16612
rect 1857 16603 1915 16609
rect 5166 16600 5172 16612
rect 5224 16600 5230 16652
rect 14 16532 20 16584
rect 72 16572 78 16584
rect 1673 16575 1731 16581
rect 1673 16572 1685 16575
rect 72 16544 1685 16572
rect 72 16532 78 16544
rect 1673 16541 1685 16544
rect 1719 16541 1731 16575
rect 1673 16535 1731 16541
rect 7006 16532 7012 16584
rect 7064 16532 7070 16584
rect 19518 16532 19524 16584
rect 19576 16572 19582 16584
rect 19981 16575 20039 16581
rect 19981 16572 19993 16575
rect 19576 16544 19993 16572
rect 19576 16532 19582 16544
rect 19981 16541 19993 16544
rect 20027 16541 20039 16575
rect 19981 16535 20039 16541
rect 20622 16532 20628 16584
rect 20680 16572 20686 16584
rect 20901 16575 20959 16581
rect 20901 16572 20913 16575
rect 20680 16544 20913 16572
rect 20680 16532 20686 16544
rect 20901 16541 20913 16544
rect 20947 16541 20959 16575
rect 20901 16535 20959 16541
rect 8113 16507 8171 16513
rect 8113 16473 8125 16507
rect 8159 16504 8171 16507
rect 17218 16504 17224 16516
rect 8159 16476 17224 16504
rect 8159 16473 8171 16476
rect 8113 16467 8171 16473
rect 17218 16464 17224 16476
rect 17276 16464 17282 16516
rect 1104 16346 45051 16368
rect 1104 16294 11896 16346
rect 11948 16294 11960 16346
rect 12012 16294 12024 16346
rect 12076 16294 12088 16346
rect 12140 16294 12152 16346
rect 12204 16294 22843 16346
rect 22895 16294 22907 16346
rect 22959 16294 22971 16346
rect 23023 16294 23035 16346
rect 23087 16294 23099 16346
rect 23151 16294 33790 16346
rect 33842 16294 33854 16346
rect 33906 16294 33918 16346
rect 33970 16294 33982 16346
rect 34034 16294 34046 16346
rect 34098 16294 44737 16346
rect 44789 16294 44801 16346
rect 44853 16294 44865 16346
rect 44917 16294 44929 16346
rect 44981 16294 44993 16346
rect 45045 16294 45051 16346
rect 1104 16272 45051 16294
rect 1026 16056 1032 16108
rect 1084 16096 1090 16108
rect 1765 16099 1823 16105
rect 1765 16096 1777 16099
rect 1084 16068 1777 16096
rect 1084 16056 1090 16068
rect 1765 16065 1777 16068
rect 1811 16065 1823 16099
rect 1765 16059 1823 16065
rect 35989 16099 36047 16105
rect 35989 16065 36001 16099
rect 36035 16096 36047 16099
rect 41598 16096 41604 16108
rect 36035 16068 41604 16096
rect 36035 16065 36047 16068
rect 35989 16059 36047 16065
rect 41598 16056 41604 16068
rect 41656 16056 41662 16108
rect 35710 15988 35716 16040
rect 35768 16028 35774 16040
rect 36081 16031 36139 16037
rect 36081 16028 36093 16031
rect 35768 16000 36093 16028
rect 35768 15988 35774 16000
rect 36081 15997 36093 16000
rect 36127 15997 36139 16031
rect 36081 15991 36139 15997
rect 36170 15988 36176 16040
rect 36228 15988 36234 16040
rect 40586 15988 40592 16040
rect 40644 16028 40650 16040
rect 41506 16028 41512 16040
rect 40644 16000 41512 16028
rect 40644 15988 40650 16000
rect 41506 15988 41512 16000
rect 41564 15988 41570 16040
rect 35621 15895 35679 15901
rect 35621 15861 35633 15895
rect 35667 15892 35679 15895
rect 36630 15892 36636 15904
rect 35667 15864 36636 15892
rect 35667 15861 35679 15864
rect 35621 15855 35679 15861
rect 36630 15852 36636 15864
rect 36688 15852 36694 15904
rect 44358 15852 44364 15904
rect 44416 15852 44422 15904
rect 1104 15802 44896 15824
rect 1104 15750 6423 15802
rect 6475 15750 6487 15802
rect 6539 15750 6551 15802
rect 6603 15750 6615 15802
rect 6667 15750 6679 15802
rect 6731 15750 17370 15802
rect 17422 15750 17434 15802
rect 17486 15750 17498 15802
rect 17550 15750 17562 15802
rect 17614 15750 17626 15802
rect 17678 15750 28317 15802
rect 28369 15750 28381 15802
rect 28433 15750 28445 15802
rect 28497 15750 28509 15802
rect 28561 15750 28573 15802
rect 28625 15750 39264 15802
rect 39316 15750 39328 15802
rect 39380 15750 39392 15802
rect 39444 15750 39456 15802
rect 39508 15750 39520 15802
rect 39572 15750 44896 15802
rect 1104 15728 44896 15750
rect 19518 15648 19524 15700
rect 19576 15648 19582 15700
rect 35710 15648 35716 15700
rect 35768 15648 35774 15700
rect 11517 15623 11575 15629
rect 11517 15589 11529 15623
rect 11563 15620 11575 15623
rect 11563 15592 12020 15620
rect 11563 15589 11575 15592
rect 11517 15583 11575 15589
rect 11992 15561 12020 15592
rect 11977 15555 12035 15561
rect 11977 15521 11989 15555
rect 12023 15521 12035 15555
rect 20073 15555 20131 15561
rect 20073 15552 20085 15555
rect 11977 15515 12035 15521
rect 17604 15524 20085 15552
rect 10134 15444 10140 15496
rect 10192 15444 10198 15496
rect 10226 15444 10232 15496
rect 10284 15484 10290 15496
rect 10393 15487 10451 15493
rect 10393 15484 10405 15487
rect 10284 15456 10405 15484
rect 10284 15444 10290 15456
rect 10393 15453 10405 15456
rect 10439 15453 10451 15487
rect 10393 15447 10451 15453
rect 17126 15444 17132 15496
rect 17184 15484 17190 15496
rect 17604 15493 17632 15524
rect 20073 15521 20085 15524
rect 20119 15521 20131 15555
rect 20073 15515 20131 15521
rect 35894 15512 35900 15564
rect 35952 15552 35958 15564
rect 36265 15555 36323 15561
rect 36265 15552 36277 15555
rect 35952 15524 36277 15552
rect 35952 15512 35958 15524
rect 36265 15521 36277 15524
rect 36311 15521 36323 15555
rect 36265 15515 36323 15521
rect 43990 15512 43996 15564
rect 44048 15512 44054 15564
rect 17589 15487 17647 15493
rect 17589 15484 17601 15487
rect 17184 15456 17601 15484
rect 17184 15444 17190 15456
rect 17589 15453 17601 15456
rect 17635 15453 17647 15487
rect 17589 15447 17647 15453
rect 17770 15444 17776 15496
rect 17828 15444 17834 15496
rect 25222 15444 25228 15496
rect 25280 15444 25286 15496
rect 41414 15444 41420 15496
rect 41472 15484 41478 15496
rect 42797 15487 42855 15493
rect 42797 15484 42809 15487
rect 41472 15456 42809 15484
rect 41472 15444 41478 15456
rect 42797 15453 42809 15456
rect 42843 15453 42855 15487
rect 42797 15447 42855 15453
rect 19886 15376 19892 15428
rect 19944 15376 19950 15428
rect 36081 15419 36139 15425
rect 36081 15385 36093 15419
rect 36127 15416 36139 15419
rect 36262 15416 36268 15428
rect 36127 15388 36268 15416
rect 36127 15385 36139 15388
rect 36081 15379 36139 15385
rect 36262 15376 36268 15388
rect 36320 15376 36326 15428
rect 12618 15308 12624 15360
rect 12676 15308 12682 15360
rect 17957 15351 18015 15357
rect 17957 15317 17969 15351
rect 18003 15348 18015 15351
rect 19794 15348 19800 15360
rect 18003 15320 19800 15348
rect 18003 15317 18015 15320
rect 17957 15311 18015 15317
rect 19794 15308 19800 15320
rect 19852 15308 19858 15360
rect 19978 15308 19984 15360
rect 20036 15308 20042 15360
rect 25041 15351 25099 15357
rect 25041 15317 25053 15351
rect 25087 15348 25099 15351
rect 25130 15348 25136 15360
rect 25087 15320 25136 15348
rect 25087 15317 25099 15320
rect 25041 15311 25099 15317
rect 25130 15308 25136 15320
rect 25188 15308 25194 15360
rect 36170 15308 36176 15360
rect 36228 15308 36234 15360
rect 1104 15258 45051 15280
rect 1104 15206 11896 15258
rect 11948 15206 11960 15258
rect 12012 15206 12024 15258
rect 12076 15206 12088 15258
rect 12140 15206 12152 15258
rect 12204 15206 22843 15258
rect 22895 15206 22907 15258
rect 22959 15206 22971 15258
rect 23023 15206 23035 15258
rect 23087 15206 23099 15258
rect 23151 15206 33790 15258
rect 33842 15206 33854 15258
rect 33906 15206 33918 15258
rect 33970 15206 33982 15258
rect 34034 15206 34046 15258
rect 34098 15206 44737 15258
rect 44789 15206 44801 15258
rect 44853 15206 44865 15258
rect 44917 15206 44929 15258
rect 44981 15206 44993 15258
rect 45045 15206 45051 15258
rect 1104 15184 45051 15206
rect 16301 15147 16359 15153
rect 16301 15113 16313 15147
rect 16347 15144 16359 15147
rect 17770 15144 17776 15156
rect 16347 15116 17776 15144
rect 16347 15113 16359 15116
rect 16301 15107 16359 15113
rect 17770 15104 17776 15116
rect 17828 15104 17834 15156
rect 18509 15147 18567 15153
rect 18509 15113 18521 15147
rect 18555 15113 18567 15147
rect 18509 15107 18567 15113
rect 18524 15076 18552 15107
rect 19978 15104 19984 15156
rect 20036 15144 20042 15156
rect 20349 15147 20407 15153
rect 20349 15144 20361 15147
rect 20036 15116 20361 15144
rect 20036 15104 20042 15116
rect 20349 15113 20361 15116
rect 20395 15113 20407 15147
rect 20349 15107 20407 15113
rect 32309 15147 32367 15153
rect 32309 15113 32321 15147
rect 32355 15113 32367 15147
rect 32309 15107 32367 15113
rect 19214 15079 19272 15085
rect 19214 15076 19226 15079
rect 11900 15048 13860 15076
rect 5626 14968 5632 15020
rect 5684 15008 5690 15020
rect 6733 15011 6791 15017
rect 6733 15008 6745 15011
rect 5684 14980 6745 15008
rect 5684 14968 5690 14980
rect 6733 14977 6745 14980
rect 6779 14977 6791 15011
rect 6733 14971 6791 14977
rect 7374 14968 7380 15020
rect 7432 14968 7438 15020
rect 11900 15017 11928 15048
rect 13832 15020 13860 15048
rect 14936 15048 17908 15076
rect 18524 15048 19226 15076
rect 11885 15011 11943 15017
rect 11885 14977 11897 15011
rect 11931 14977 11943 15011
rect 11885 14971 11943 14977
rect 12152 15011 12210 15017
rect 12152 14977 12164 15011
rect 12198 15008 12210 15011
rect 12618 15008 12624 15020
rect 12198 14980 12624 15008
rect 12198 14977 12210 14980
rect 12152 14971 12210 14977
rect 12618 14968 12624 14980
rect 12676 14968 12682 15020
rect 13814 14968 13820 15020
rect 13872 15008 13878 15020
rect 14936 15017 14964 15048
rect 15194 15017 15200 15020
rect 14921 15011 14979 15017
rect 14921 15008 14933 15011
rect 13872 14980 14933 15008
rect 13872 14968 13878 14980
rect 14921 14977 14933 14980
rect 14967 14977 14979 15011
rect 14921 14971 14979 14977
rect 15188 14971 15200 15017
rect 15194 14968 15200 14971
rect 15252 14968 15258 15020
rect 17144 15017 17172 15048
rect 17880 15020 17908 15048
rect 19214 15045 19226 15048
rect 19260 15076 19272 15079
rect 19702 15076 19708 15088
rect 19260 15048 19708 15076
rect 19260 15045 19272 15048
rect 19214 15039 19272 15045
rect 19702 15036 19708 15048
rect 19760 15036 19766 15088
rect 23032 15048 24900 15076
rect 17129 15011 17187 15017
rect 17129 14977 17141 15011
rect 17175 14977 17187 15011
rect 17129 14971 17187 14977
rect 17218 14968 17224 15020
rect 17276 15008 17282 15020
rect 17385 15011 17443 15017
rect 17385 15008 17397 15011
rect 17276 14980 17397 15008
rect 17276 14968 17282 14980
rect 17385 14977 17397 14980
rect 17431 14977 17443 15011
rect 17385 14971 17443 14977
rect 17862 14968 17868 15020
rect 17920 15008 17926 15020
rect 18969 15011 19027 15017
rect 18969 15008 18981 15011
rect 17920 14980 18981 15008
rect 17920 14968 17926 14980
rect 18969 14977 18981 14980
rect 19015 14977 19027 15011
rect 18969 14971 19027 14977
rect 19794 14968 19800 15020
rect 19852 15008 19858 15020
rect 20993 15011 21051 15017
rect 20993 15008 21005 15011
rect 19852 14980 21005 15008
rect 19852 14968 19858 14980
rect 20993 14977 21005 14980
rect 21039 14977 21051 15011
rect 20993 14971 21051 14977
rect 22094 14968 22100 15020
rect 22152 15008 22158 15020
rect 23032 15017 23060 15048
rect 24872 15020 24900 15048
rect 30116 15048 31754 15076
rect 23017 15011 23075 15017
rect 23017 15008 23029 15011
rect 22152 14980 23029 15008
rect 22152 14968 22158 14980
rect 23017 14977 23029 14980
rect 23063 14977 23075 15011
rect 23273 15011 23331 15017
rect 23273 15008 23285 15011
rect 23017 14971 23075 14977
rect 23124 14980 23285 15008
rect 23124 14940 23152 14980
rect 23273 14977 23285 14980
rect 23319 14977 23331 15011
rect 23273 14971 23331 14977
rect 24854 14968 24860 15020
rect 24912 14968 24918 15020
rect 25130 15017 25136 15020
rect 25124 15008 25136 15017
rect 25091 14980 25136 15008
rect 25124 14971 25136 14980
rect 25130 14968 25136 14971
rect 25188 14968 25194 15020
rect 27706 14968 27712 15020
rect 27764 15008 27770 15020
rect 28793 15011 28851 15017
rect 28793 15008 28805 15011
rect 27764 14980 28805 15008
rect 27764 14968 27770 14980
rect 28793 14977 28805 14980
rect 28839 15008 28851 15011
rect 30116 15008 30144 15048
rect 28839 14980 30144 15008
rect 28839 14977 28851 14980
rect 28793 14971 28851 14977
rect 30190 14968 30196 15020
rect 30248 15008 30254 15020
rect 30745 15011 30803 15017
rect 30745 15008 30757 15011
rect 30248 14980 30757 15008
rect 30248 14968 30254 14980
rect 30745 14977 30757 14980
rect 30791 14977 30803 15011
rect 30745 14971 30803 14977
rect 31386 14968 31392 15020
rect 31444 14968 31450 15020
rect 31726 15008 31754 15048
rect 32030 15036 32036 15088
rect 32088 15076 32094 15088
rect 32324 15076 32352 15107
rect 32582 15104 32588 15156
rect 32640 15144 32646 15156
rect 32677 15147 32735 15153
rect 32677 15144 32689 15147
rect 32640 15116 32689 15144
rect 32640 15104 32646 15116
rect 32677 15113 32689 15116
rect 32723 15113 32735 15147
rect 32677 15107 32735 15113
rect 33965 15147 34023 15153
rect 33965 15113 33977 15147
rect 34011 15113 34023 15147
rect 33965 15107 34023 15113
rect 32088 15048 32352 15076
rect 32088 15036 32094 15048
rect 32600 15008 32628 15104
rect 33980 15076 34008 15107
rect 34854 15079 34912 15085
rect 34854 15076 34866 15079
rect 33980 15048 34866 15076
rect 34854 15045 34866 15048
rect 34900 15045 34912 15079
rect 34854 15039 34912 15045
rect 31726 14980 32628 15008
rect 32769 15011 32827 15017
rect 32769 14977 32781 15011
rect 32815 15008 32827 15011
rect 32815 14980 33548 15008
rect 32815 14977 32827 14980
rect 32769 14971 32827 14977
rect 22066 14912 23152 14940
rect 28537 14943 28595 14949
rect 20809 14875 20867 14881
rect 18340 14844 18644 14872
rect 6549 14807 6607 14813
rect 6549 14773 6561 14807
rect 6595 14804 6607 14807
rect 6822 14804 6828 14816
rect 6595 14776 6828 14804
rect 6595 14773 6607 14776
rect 6549 14767 6607 14773
rect 6822 14764 6828 14776
rect 6880 14764 6886 14816
rect 7190 14764 7196 14816
rect 7248 14764 7254 14816
rect 13265 14807 13323 14813
rect 13265 14773 13277 14807
rect 13311 14804 13323 14807
rect 18340 14804 18368 14844
rect 13311 14776 18368 14804
rect 18616 14804 18644 14844
rect 20809 14841 20821 14875
rect 20855 14872 20867 14875
rect 22066 14872 22094 14912
rect 28537 14909 28549 14943
rect 28583 14909 28595 14943
rect 28537 14903 28595 14909
rect 20855 14844 22094 14872
rect 20855 14841 20867 14844
rect 20809 14835 20867 14841
rect 22370 14804 22376 14816
rect 18616 14776 22376 14804
rect 13311 14773 13323 14776
rect 13265 14767 13323 14773
rect 22370 14764 22376 14776
rect 22428 14764 22434 14816
rect 24394 14764 24400 14816
rect 24452 14764 24458 14816
rect 26237 14807 26295 14813
rect 26237 14773 26249 14807
rect 26283 14804 26295 14807
rect 26602 14804 26608 14816
rect 26283 14776 26608 14804
rect 26283 14773 26295 14776
rect 26237 14767 26295 14773
rect 26602 14764 26608 14776
rect 26660 14764 26666 14816
rect 28552 14804 28580 14903
rect 29546 14900 29552 14952
rect 29604 14940 29610 14952
rect 32861 14943 32919 14949
rect 29604 14912 32352 14940
rect 29604 14900 29610 14912
rect 29638 14832 29644 14884
rect 29696 14872 29702 14884
rect 32324 14872 32352 14912
rect 32861 14909 32873 14943
rect 32907 14909 32919 14943
rect 33520 14940 33548 14980
rect 33594 14968 33600 15020
rect 33652 15008 33658 15020
rect 34149 15011 34207 15017
rect 34149 15008 34161 15011
rect 33652 14980 34161 15008
rect 33652 14968 33658 14980
rect 34149 14977 34161 14980
rect 34195 14977 34207 15011
rect 34149 14971 34207 14977
rect 36630 14968 36636 15020
rect 36688 14968 36694 15020
rect 40037 15011 40095 15017
rect 40037 14977 40049 15011
rect 40083 15008 40095 15011
rect 40126 15008 40132 15020
rect 40083 14980 40132 15008
rect 40083 14977 40095 14980
rect 40037 14971 40095 14977
rect 40126 14968 40132 14980
rect 40184 14968 40190 15020
rect 34514 14940 34520 14952
rect 33520 14912 34520 14940
rect 32861 14903 32919 14909
rect 32876 14872 32904 14903
rect 34514 14900 34520 14912
rect 34572 14900 34578 14952
rect 34606 14900 34612 14952
rect 34664 14900 34670 14952
rect 38930 14900 38936 14952
rect 38988 14940 38994 14952
rect 39853 14943 39911 14949
rect 39853 14940 39865 14943
rect 38988 14912 39865 14940
rect 38988 14900 38994 14912
rect 39853 14909 39865 14912
rect 39899 14909 39911 14943
rect 39853 14903 39911 14909
rect 29696 14844 32260 14872
rect 32324 14844 32904 14872
rect 35989 14875 36047 14881
rect 29696 14832 29702 14844
rect 28902 14804 28908 14816
rect 28552 14776 28908 14804
rect 28902 14764 28908 14776
rect 28960 14764 28966 14816
rect 29917 14807 29975 14813
rect 29917 14773 29929 14807
rect 29963 14804 29975 14807
rect 30006 14804 30012 14816
rect 29963 14776 30012 14804
rect 29963 14773 29975 14776
rect 29917 14767 29975 14773
rect 30006 14764 30012 14776
rect 30064 14764 30070 14816
rect 30561 14807 30619 14813
rect 30561 14773 30573 14807
rect 30607 14804 30619 14807
rect 31110 14804 31116 14816
rect 30607 14776 31116 14804
rect 30607 14773 30619 14776
rect 30561 14767 30619 14773
rect 31110 14764 31116 14776
rect 31168 14764 31174 14816
rect 31202 14764 31208 14816
rect 31260 14764 31266 14816
rect 32232 14804 32260 14844
rect 35989 14841 36001 14875
rect 36035 14872 36047 14875
rect 36170 14872 36176 14884
rect 36035 14844 36176 14872
rect 36035 14841 36047 14844
rect 35989 14835 36047 14841
rect 36170 14832 36176 14844
rect 36228 14872 36234 14884
rect 37090 14872 37096 14884
rect 36228 14844 37096 14872
rect 36228 14832 36234 14844
rect 37090 14832 37096 14844
rect 37148 14832 37154 14884
rect 36262 14804 36268 14816
rect 32232 14776 36268 14804
rect 36262 14764 36268 14776
rect 36320 14764 36326 14816
rect 36446 14764 36452 14816
rect 36504 14764 36510 14816
rect 39666 14764 39672 14816
rect 39724 14804 39730 14816
rect 40221 14807 40279 14813
rect 40221 14804 40233 14807
rect 39724 14776 40233 14804
rect 39724 14764 39730 14776
rect 40221 14773 40233 14776
rect 40267 14773 40279 14807
rect 40221 14767 40279 14773
rect 1104 14714 44896 14736
rect 1104 14662 6423 14714
rect 6475 14662 6487 14714
rect 6539 14662 6551 14714
rect 6603 14662 6615 14714
rect 6667 14662 6679 14714
rect 6731 14662 17370 14714
rect 17422 14662 17434 14714
rect 17486 14662 17498 14714
rect 17550 14662 17562 14714
rect 17614 14662 17626 14714
rect 17678 14662 28317 14714
rect 28369 14662 28381 14714
rect 28433 14662 28445 14714
rect 28497 14662 28509 14714
rect 28561 14662 28573 14714
rect 28625 14662 39264 14714
rect 39316 14662 39328 14714
rect 39380 14662 39392 14714
rect 39444 14662 39456 14714
rect 39508 14662 39520 14714
rect 39572 14662 44896 14714
rect 1104 14640 44896 14662
rect 5626 14560 5632 14612
rect 5684 14560 5690 14612
rect 5810 14560 5816 14612
rect 5868 14600 5874 14612
rect 6457 14603 6515 14609
rect 6457 14600 6469 14603
rect 5868 14572 6469 14600
rect 5868 14560 5874 14572
rect 6457 14569 6469 14572
rect 6503 14600 6515 14603
rect 7834 14600 7840 14612
rect 6503 14572 7840 14600
rect 6503 14569 6515 14572
rect 6457 14563 6515 14569
rect 7834 14560 7840 14572
rect 7892 14560 7898 14612
rect 17218 14560 17224 14612
rect 17276 14600 17282 14612
rect 17497 14603 17555 14609
rect 17497 14600 17509 14603
rect 17276 14572 17509 14600
rect 17276 14560 17282 14572
rect 17497 14569 17509 14572
rect 17543 14569 17555 14603
rect 25041 14603 25099 14609
rect 17497 14563 17555 14569
rect 18064 14572 22094 14600
rect 6641 14535 6699 14541
rect 6641 14501 6653 14535
rect 6687 14501 6699 14535
rect 6641 14495 6699 14501
rect 12897 14535 12955 14541
rect 12897 14501 12909 14535
rect 12943 14501 12955 14535
rect 12897 14495 12955 14501
rect 15289 14535 15347 14541
rect 15289 14501 15301 14535
rect 15335 14532 15347 14535
rect 15335 14504 15884 14532
rect 15335 14501 15347 14504
rect 15289 14495 15347 14501
rect 6656 14464 6684 14495
rect 5828 14436 6684 14464
rect 4706 14356 4712 14408
rect 4764 14356 4770 14408
rect 4893 14399 4951 14405
rect 4893 14365 4905 14399
rect 4939 14365 4951 14399
rect 4893 14359 4951 14365
rect 4338 14288 4344 14340
rect 4396 14328 4402 14340
rect 4908 14328 4936 14359
rect 5626 14356 5632 14408
rect 5684 14356 5690 14408
rect 5718 14356 5724 14408
rect 5776 14396 5782 14408
rect 5828 14405 5856 14436
rect 10134 14424 10140 14476
rect 10192 14464 10198 14476
rect 11517 14467 11575 14473
rect 11517 14464 11529 14467
rect 10192 14436 11529 14464
rect 10192 14424 10198 14436
rect 11517 14433 11529 14436
rect 11563 14433 11575 14467
rect 11517 14427 11575 14433
rect 5813 14399 5871 14405
rect 5813 14396 5825 14399
rect 5776 14368 5825 14396
rect 5776 14356 5782 14368
rect 5813 14365 5825 14368
rect 5859 14365 5871 14399
rect 5813 14359 5871 14365
rect 6546 14356 6552 14408
rect 6604 14396 6610 14408
rect 7101 14399 7159 14405
rect 7101 14396 7113 14399
rect 6604 14368 7113 14396
rect 6604 14356 6610 14368
rect 7101 14365 7113 14368
rect 7147 14365 7159 14399
rect 7101 14359 7159 14365
rect 7190 14356 7196 14408
rect 7248 14396 7254 14408
rect 7357 14399 7415 14405
rect 7357 14396 7369 14399
rect 7248 14368 7369 14396
rect 7248 14356 7254 14368
rect 7357 14365 7369 14368
rect 7403 14365 7415 14399
rect 7357 14359 7415 14365
rect 11057 14399 11115 14405
rect 11057 14365 11069 14399
rect 11103 14396 11115 14399
rect 12250 14396 12256 14408
rect 11103 14368 12256 14396
rect 11103 14365 11115 14368
rect 11057 14359 11115 14365
rect 12250 14356 12256 14368
rect 12308 14356 12314 14408
rect 12912 14396 12940 14495
rect 13357 14399 13415 14405
rect 13357 14396 13369 14399
rect 12912 14368 13369 14396
rect 13357 14365 13369 14368
rect 13403 14365 13415 14399
rect 13357 14359 13415 14365
rect 14274 14356 14280 14408
rect 14332 14356 14338 14408
rect 14458 14356 14464 14408
rect 14516 14356 14522 14408
rect 15654 14356 15660 14408
rect 15712 14356 15718 14408
rect 15856 14396 15884 14504
rect 15933 14467 15991 14473
rect 15933 14433 15945 14467
rect 15979 14464 15991 14467
rect 18064 14464 18092 14572
rect 18141 14535 18199 14541
rect 18141 14501 18153 14535
rect 18187 14501 18199 14535
rect 19886 14532 19892 14544
rect 18141 14495 18199 14501
rect 18248 14504 19892 14532
rect 15979 14436 18092 14464
rect 15979 14433 15991 14436
rect 15933 14427 15991 14433
rect 17681 14399 17739 14405
rect 15856 14368 17632 14396
rect 4396 14300 4936 14328
rect 6273 14331 6331 14337
rect 4396 14288 4402 14300
rect 6273 14297 6285 14331
rect 6319 14328 6331 14331
rect 11762 14331 11820 14337
rect 11762 14328 11774 14331
rect 6319 14300 8524 14328
rect 6319 14297 6331 14300
rect 6273 14291 6331 14297
rect 8496 14272 8524 14300
rect 10888 14300 11774 14328
rect 4154 14220 4160 14272
rect 4212 14260 4218 14272
rect 4801 14263 4859 14269
rect 4801 14260 4813 14263
rect 4212 14232 4813 14260
rect 4212 14220 4218 14232
rect 4801 14229 4813 14232
rect 4847 14229 4859 14263
rect 4801 14223 4859 14229
rect 6483 14263 6541 14269
rect 6483 14229 6495 14263
rect 6529 14260 6541 14263
rect 8202 14260 8208 14272
rect 6529 14232 8208 14260
rect 6529 14229 6541 14232
rect 6483 14223 6541 14229
rect 8202 14220 8208 14232
rect 8260 14220 8266 14272
rect 8478 14220 8484 14272
rect 8536 14220 8542 14272
rect 10888 14269 10916 14300
rect 11762 14297 11774 14300
rect 11808 14297 11820 14331
rect 14369 14331 14427 14337
rect 14369 14328 14381 14331
rect 11762 14291 11820 14297
rect 11900 14300 14381 14328
rect 10873 14263 10931 14269
rect 10873 14229 10885 14263
rect 10919 14229 10931 14263
rect 10873 14223 10931 14229
rect 11330 14220 11336 14272
rect 11388 14260 11394 14272
rect 11900 14260 11928 14300
rect 14369 14297 14381 14300
rect 14415 14328 14427 14331
rect 15286 14328 15292 14340
rect 14415 14300 15292 14328
rect 14415 14297 14427 14300
rect 14369 14291 14427 14297
rect 15286 14288 15292 14300
rect 15344 14288 15350 14340
rect 15470 14288 15476 14340
rect 15528 14328 15534 14340
rect 15749 14331 15807 14337
rect 15749 14328 15761 14331
rect 15528 14300 15761 14328
rect 15528 14288 15534 14300
rect 15749 14297 15761 14300
rect 15795 14297 15807 14331
rect 17604 14328 17632 14368
rect 17681 14365 17693 14399
rect 17727 14396 17739 14399
rect 18156 14396 18184 14495
rect 17727 14368 18184 14396
rect 17727 14365 17739 14368
rect 17681 14359 17739 14365
rect 18248 14328 18276 14504
rect 19886 14492 19892 14504
rect 19944 14492 19950 14544
rect 22066 14532 22094 14572
rect 25041 14569 25053 14603
rect 25087 14600 25099 14603
rect 25222 14600 25228 14612
rect 25087 14572 25228 14600
rect 25087 14569 25099 14572
rect 25041 14563 25099 14569
rect 25222 14560 25228 14572
rect 25280 14560 25286 14612
rect 29638 14600 29644 14612
rect 26712 14572 29644 14600
rect 22066 14504 23888 14532
rect 23860 14476 23888 14504
rect 18785 14467 18843 14473
rect 18785 14433 18797 14467
rect 18831 14464 18843 14467
rect 19978 14464 19984 14476
rect 18831 14436 19984 14464
rect 18831 14433 18843 14436
rect 18785 14427 18843 14433
rect 19978 14424 19984 14436
rect 20036 14424 20042 14476
rect 20073 14467 20131 14473
rect 20073 14433 20085 14467
rect 20119 14464 20131 14467
rect 20990 14464 20996 14476
rect 20119 14436 20996 14464
rect 20119 14433 20131 14436
rect 20073 14427 20131 14433
rect 20990 14424 20996 14436
rect 21048 14424 21054 14476
rect 23750 14424 23756 14476
rect 23808 14424 23814 14476
rect 23842 14424 23848 14476
rect 23900 14424 23906 14476
rect 25498 14424 25504 14476
rect 25556 14464 25562 14476
rect 26712 14473 26740 14572
rect 29638 14560 29644 14572
rect 29696 14560 29702 14612
rect 30101 14603 30159 14609
rect 30101 14569 30113 14603
rect 30147 14600 30159 14603
rect 31386 14600 31392 14612
rect 30147 14572 31392 14600
rect 30147 14569 30159 14572
rect 30101 14563 30159 14569
rect 31386 14560 31392 14572
rect 31444 14560 31450 14612
rect 33594 14560 33600 14612
rect 33652 14560 33658 14612
rect 36725 14603 36783 14609
rect 36725 14600 36737 14603
rect 34072 14572 36737 14600
rect 29181 14535 29239 14541
rect 29181 14501 29193 14535
rect 29227 14501 29239 14535
rect 29181 14495 29239 14501
rect 25593 14467 25651 14473
rect 25593 14464 25605 14467
rect 25556 14436 25605 14464
rect 25556 14424 25562 14436
rect 25593 14433 25605 14436
rect 25639 14433 25651 14467
rect 25593 14427 25651 14433
rect 26697 14467 26755 14473
rect 26697 14433 26709 14467
rect 26743 14433 26755 14467
rect 26697 14427 26755 14433
rect 26786 14424 26792 14476
rect 26844 14424 26850 14476
rect 29196 14464 29224 14495
rect 34072 14473 34100 14572
rect 36725 14569 36737 14572
rect 36771 14569 36783 14603
rect 36725 14563 36783 14569
rect 41417 14603 41475 14609
rect 41417 14569 41429 14603
rect 41463 14600 41475 14603
rect 41598 14600 41604 14612
rect 41463 14572 41604 14600
rect 41463 14569 41475 14572
rect 41417 14563 41475 14569
rect 41598 14560 41604 14572
rect 41656 14560 41662 14612
rect 36262 14492 36268 14544
rect 36320 14492 36326 14544
rect 34057 14467 34115 14473
rect 29196 14436 29960 14464
rect 17604 14300 18276 14328
rect 18432 14368 19472 14396
rect 15749 14291 15807 14297
rect 11388 14232 11928 14260
rect 11388 14220 11394 14232
rect 12342 14220 12348 14272
rect 12400 14260 12406 14272
rect 13449 14263 13507 14269
rect 13449 14260 13461 14263
rect 12400 14232 13461 14260
rect 12400 14220 12406 14232
rect 13449 14229 13461 14232
rect 13495 14260 13507 14263
rect 13538 14260 13544 14272
rect 13495 14232 13544 14260
rect 13495 14229 13507 14232
rect 13449 14223 13507 14229
rect 13538 14220 13544 14232
rect 13596 14220 13602 14272
rect 15654 14220 15660 14272
rect 15712 14260 15718 14272
rect 18432 14260 18460 14368
rect 19444 14328 19472 14368
rect 19702 14356 19708 14408
rect 19760 14396 19766 14408
rect 19797 14399 19855 14405
rect 19797 14396 19809 14399
rect 19760 14368 19809 14396
rect 19760 14356 19766 14368
rect 19797 14365 19809 14368
rect 19843 14365 19855 14399
rect 19797 14359 19855 14365
rect 22097 14399 22155 14405
rect 22097 14365 22109 14399
rect 22143 14396 22155 14399
rect 22186 14396 22192 14408
rect 22143 14368 22192 14396
rect 22143 14365 22155 14368
rect 22097 14359 22155 14365
rect 22186 14356 22192 14368
rect 22244 14356 22250 14408
rect 23584 14368 23796 14396
rect 20622 14328 20628 14340
rect 19444 14300 20628 14328
rect 20622 14288 20628 14300
rect 20680 14328 20686 14340
rect 23584 14328 23612 14368
rect 20680 14300 23612 14328
rect 20680 14288 20686 14300
rect 23658 14288 23664 14340
rect 23716 14288 23722 14340
rect 23768 14328 23796 14368
rect 24394 14356 24400 14408
rect 24452 14396 24458 14408
rect 25409 14399 25467 14405
rect 25409 14396 25421 14399
rect 24452 14368 25421 14396
rect 24452 14356 24458 14368
rect 25409 14365 25421 14368
rect 25455 14365 25467 14399
rect 25409 14359 25467 14365
rect 26602 14356 26608 14408
rect 26660 14356 26666 14408
rect 27798 14356 27804 14408
rect 27856 14396 27862 14408
rect 28902 14396 28908 14408
rect 27856 14368 28908 14396
rect 27856 14356 27862 14368
rect 28902 14356 28908 14368
rect 28960 14356 28966 14408
rect 29730 14356 29736 14408
rect 29788 14356 29794 14408
rect 29932 14405 29960 14436
rect 34057 14433 34069 14467
rect 34103 14433 34115 14467
rect 34057 14427 34115 14433
rect 34149 14467 34207 14473
rect 34149 14433 34161 14467
rect 34195 14433 34207 14467
rect 34149 14427 34207 14433
rect 29917 14399 29975 14405
rect 29917 14365 29929 14399
rect 29963 14365 29975 14399
rect 29917 14359 29975 14365
rect 30926 14356 30932 14408
rect 30984 14396 30990 14408
rect 31021 14399 31079 14405
rect 31021 14396 31033 14399
rect 30984 14368 31033 14396
rect 30984 14356 30990 14368
rect 31021 14365 31033 14368
rect 31067 14365 31079 14399
rect 31021 14359 31079 14365
rect 31110 14356 31116 14408
rect 31168 14396 31174 14408
rect 31277 14399 31335 14405
rect 31277 14396 31289 14399
rect 31168 14368 31289 14396
rect 31168 14356 31174 14368
rect 31277 14365 31289 14368
rect 31323 14365 31335 14399
rect 31277 14359 31335 14365
rect 32398 14356 32404 14408
rect 32456 14396 32462 14408
rect 34164 14396 34192 14427
rect 35894 14424 35900 14476
rect 35952 14464 35958 14476
rect 37369 14467 37427 14473
rect 37369 14464 37381 14467
rect 35952 14436 37381 14464
rect 35952 14424 35958 14436
rect 37369 14433 37381 14436
rect 37415 14464 37427 14467
rect 38194 14464 38200 14476
rect 37415 14436 38200 14464
rect 37415 14433 37427 14436
rect 37369 14427 37427 14433
rect 38194 14424 38200 14436
rect 38252 14424 38258 14476
rect 32456 14368 34192 14396
rect 32456 14356 32462 14368
rect 28046 14331 28104 14337
rect 28046 14328 28058 14331
rect 23768 14300 28058 14328
rect 28046 14297 28058 14300
rect 28092 14297 28104 14331
rect 33965 14331 34023 14337
rect 33965 14328 33977 14331
rect 28046 14291 28104 14297
rect 32416 14300 33977 14328
rect 15712 14232 18460 14260
rect 15712 14220 15718 14232
rect 18506 14220 18512 14272
rect 18564 14220 18570 14272
rect 18601 14263 18659 14269
rect 18601 14229 18613 14263
rect 18647 14260 18659 14263
rect 19429 14263 19487 14269
rect 19429 14260 19441 14263
rect 18647 14232 19441 14260
rect 18647 14229 18659 14232
rect 18601 14223 18659 14229
rect 19429 14229 19441 14232
rect 19475 14229 19487 14263
rect 19429 14223 19487 14229
rect 19886 14220 19892 14272
rect 19944 14220 19950 14272
rect 21910 14220 21916 14272
rect 21968 14220 21974 14272
rect 23293 14263 23351 14269
rect 23293 14229 23305 14263
rect 23339 14260 23351 14263
rect 23566 14260 23572 14272
rect 23339 14232 23572 14260
rect 23339 14229 23351 14232
rect 23293 14223 23351 14229
rect 23566 14220 23572 14232
rect 23624 14220 23630 14272
rect 25501 14263 25559 14269
rect 25501 14229 25513 14263
rect 25547 14260 25559 14263
rect 26237 14263 26295 14269
rect 26237 14260 26249 14263
rect 25547 14232 26249 14260
rect 25547 14229 25559 14232
rect 25501 14223 25559 14229
rect 26237 14229 26249 14232
rect 26283 14229 26295 14263
rect 26237 14223 26295 14229
rect 26786 14220 26792 14272
rect 26844 14260 26850 14272
rect 31110 14260 31116 14272
rect 26844 14232 31116 14260
rect 26844 14220 26850 14232
rect 31110 14220 31116 14232
rect 31168 14220 31174 14272
rect 32416 14269 32444 14300
rect 33965 14297 33977 14300
rect 34011 14297 34023 14331
rect 33965 14291 34023 14297
rect 32401 14263 32459 14269
rect 32401 14229 32413 14263
rect 32447 14229 32459 14263
rect 34164 14260 34192 14368
rect 34606 14356 34612 14408
rect 34664 14396 34670 14408
rect 34885 14399 34943 14405
rect 34885 14396 34897 14399
rect 34664 14368 34897 14396
rect 34664 14356 34670 14368
rect 34885 14365 34897 14368
rect 34931 14396 34943 14399
rect 36354 14396 36360 14408
rect 34931 14368 36360 14396
rect 34931 14365 34943 14368
rect 34885 14359 34943 14365
rect 36354 14356 36360 14368
rect 36412 14356 36418 14408
rect 37090 14356 37096 14408
rect 37148 14356 37154 14408
rect 39485 14399 39543 14405
rect 39485 14365 39497 14399
rect 39531 14396 39543 14399
rect 39666 14396 39672 14408
rect 39531 14368 39672 14396
rect 39531 14365 39543 14368
rect 39485 14359 39543 14365
rect 39666 14356 39672 14368
rect 39724 14356 39730 14408
rect 40034 14356 40040 14408
rect 40092 14356 40098 14408
rect 41690 14356 41696 14408
rect 41748 14396 41754 14408
rect 42797 14399 42855 14405
rect 42797 14396 42809 14399
rect 41748 14368 42809 14396
rect 41748 14356 41754 14368
rect 42797 14365 42809 14368
rect 42843 14365 42855 14399
rect 42797 14359 42855 14365
rect 35152 14331 35210 14337
rect 35152 14297 35164 14331
rect 35198 14328 35210 14331
rect 36446 14328 36452 14340
rect 35198 14300 36452 14328
rect 35198 14297 35210 14300
rect 35152 14291 35210 14297
rect 36446 14288 36452 14300
rect 36504 14288 36510 14340
rect 40282 14331 40340 14337
rect 40282 14328 40294 14331
rect 39316 14300 40294 14328
rect 36078 14260 36084 14272
rect 34164 14232 36084 14260
rect 32401 14223 32459 14229
rect 36078 14220 36084 14232
rect 36136 14260 36142 14272
rect 36262 14260 36268 14272
rect 36136 14232 36268 14260
rect 36136 14220 36142 14232
rect 36262 14220 36268 14232
rect 36320 14220 36326 14272
rect 37185 14263 37243 14269
rect 37185 14229 37197 14263
rect 37231 14260 37243 14263
rect 37826 14260 37832 14272
rect 37231 14232 37832 14260
rect 37231 14229 37243 14232
rect 37185 14223 37243 14229
rect 37826 14220 37832 14232
rect 37884 14220 37890 14272
rect 39316 14269 39344 14300
rect 40282 14297 40294 14300
rect 40328 14297 40340 14331
rect 40282 14291 40340 14297
rect 43993 14331 44051 14337
rect 43993 14297 44005 14331
rect 44039 14328 44051 14331
rect 45002 14328 45008 14340
rect 44039 14300 45008 14328
rect 44039 14297 44051 14300
rect 43993 14291 44051 14297
rect 45002 14288 45008 14300
rect 45060 14288 45066 14340
rect 39301 14263 39359 14269
rect 39301 14229 39313 14263
rect 39347 14229 39359 14263
rect 39301 14223 39359 14229
rect 1104 14170 45051 14192
rect 1104 14118 11896 14170
rect 11948 14118 11960 14170
rect 12012 14118 12024 14170
rect 12076 14118 12088 14170
rect 12140 14118 12152 14170
rect 12204 14118 22843 14170
rect 22895 14118 22907 14170
rect 22959 14118 22971 14170
rect 23023 14118 23035 14170
rect 23087 14118 23099 14170
rect 23151 14118 33790 14170
rect 33842 14118 33854 14170
rect 33906 14118 33918 14170
rect 33970 14118 33982 14170
rect 34034 14118 34046 14170
rect 34098 14118 44737 14170
rect 44789 14118 44801 14170
rect 44853 14118 44865 14170
rect 44917 14118 44929 14170
rect 44981 14118 44993 14170
rect 45045 14118 45051 14170
rect 1104 14096 45051 14118
rect 4706 14016 4712 14068
rect 4764 14056 4770 14068
rect 5261 14059 5319 14065
rect 5261 14056 5273 14059
rect 4764 14028 5273 14056
rect 4764 14016 4770 14028
rect 5261 14025 5273 14028
rect 5307 14025 5319 14059
rect 5261 14019 5319 14025
rect 5626 14016 5632 14068
rect 5684 14056 5690 14068
rect 5997 14059 6055 14065
rect 5997 14056 6009 14059
rect 5684 14028 6009 14056
rect 5684 14016 5690 14028
rect 5997 14025 6009 14028
rect 6043 14025 6055 14059
rect 5997 14019 6055 14025
rect 7834 14016 7840 14068
rect 7892 14056 7898 14068
rect 7929 14059 7987 14065
rect 7929 14056 7941 14059
rect 7892 14028 7941 14056
rect 7892 14016 7898 14028
rect 7929 14025 7941 14028
rect 7975 14056 7987 14059
rect 9766 14056 9772 14068
rect 7975 14028 9772 14056
rect 7975 14025 7987 14028
rect 7929 14019 7987 14025
rect 9766 14016 9772 14028
rect 9824 14016 9830 14068
rect 12250 14016 12256 14068
rect 12308 14016 12314 14068
rect 14274 14016 14280 14068
rect 14332 14056 14338 14068
rect 14921 14059 14979 14065
rect 14921 14056 14933 14059
rect 14332 14028 14933 14056
rect 14332 14016 14338 14028
rect 14921 14025 14933 14028
rect 14967 14025 14979 14059
rect 14921 14019 14979 14025
rect 15381 14059 15439 14065
rect 15381 14025 15393 14059
rect 15427 14025 15439 14059
rect 15381 14019 15439 14025
rect 17865 14059 17923 14065
rect 17865 14025 17877 14059
rect 17911 14025 17923 14059
rect 17865 14019 17923 14025
rect 5534 13948 5540 14000
rect 5592 13988 5598 14000
rect 6822 13997 6828 14000
rect 6816 13988 6828 13997
rect 5592 13960 6592 13988
rect 6783 13960 6828 13988
rect 5592 13948 5598 13960
rect 6564 13932 6592 13960
rect 6816 13951 6828 13960
rect 6822 13948 6828 13951
rect 6880 13948 6886 14000
rect 8202 13948 8208 14000
rect 8260 13988 8266 14000
rect 8389 13991 8447 13997
rect 8389 13988 8401 13991
rect 8260 13960 8401 13988
rect 8260 13948 8266 13960
rect 8389 13957 8401 13960
rect 8435 13988 8447 13991
rect 11238 13988 11244 14000
rect 8435 13960 11244 13988
rect 8435 13957 8447 13960
rect 8389 13951 8447 13957
rect 11238 13948 11244 13960
rect 11296 13948 11302 14000
rect 12069 13991 12127 13997
rect 12069 13957 12081 13991
rect 12115 13988 12127 13991
rect 13808 13991 13866 13997
rect 12115 13960 13768 13988
rect 12115 13957 12127 13960
rect 12069 13951 12127 13957
rect 1026 13880 1032 13932
rect 1084 13920 1090 13932
rect 1084 13892 1900 13920
rect 1084 13880 1090 13892
rect 934 13812 940 13864
rect 992 13852 998 13864
rect 1765 13855 1823 13861
rect 1765 13852 1777 13855
rect 992 13824 1777 13852
rect 992 13812 998 13824
rect 1765 13821 1777 13824
rect 1811 13821 1823 13855
rect 1872 13852 1900 13892
rect 3050 13880 3056 13932
rect 3108 13880 3114 13932
rect 4982 13880 4988 13932
rect 5040 13880 5046 13932
rect 5721 13923 5779 13929
rect 5721 13889 5733 13923
rect 5767 13920 5779 13923
rect 5810 13920 5816 13932
rect 5767 13892 5816 13920
rect 5767 13889 5779 13892
rect 5721 13883 5779 13889
rect 5810 13880 5816 13892
rect 5868 13880 5874 13932
rect 6546 13880 6552 13932
rect 6604 13880 6610 13932
rect 7098 13920 7104 13932
rect 6656 13892 7104 13920
rect 3329 13855 3387 13861
rect 3329 13852 3341 13855
rect 1872 13824 3341 13852
rect 1765 13815 1823 13821
rect 3329 13821 3341 13824
rect 3375 13821 3387 13855
rect 3329 13815 3387 13821
rect 5258 13812 5264 13864
rect 5316 13852 5322 13864
rect 5997 13855 6055 13861
rect 5997 13852 6009 13855
rect 5316 13824 6009 13852
rect 5316 13812 5322 13824
rect 5997 13821 6009 13824
rect 6043 13852 6055 13855
rect 6656 13852 6684 13892
rect 7098 13880 7104 13892
rect 7156 13920 7162 13932
rect 7156 13892 7696 13920
rect 7156 13880 7162 13892
rect 6043 13824 6684 13852
rect 7668 13852 7696 13892
rect 8478 13880 8484 13932
rect 8536 13920 8542 13932
rect 8573 13923 8631 13929
rect 8573 13920 8585 13923
rect 8536 13892 8585 13920
rect 8536 13880 8542 13892
rect 8573 13889 8585 13892
rect 8619 13920 8631 13923
rect 9398 13920 9404 13932
rect 8619 13892 9404 13920
rect 8619 13889 8631 13892
rect 8573 13883 8631 13889
rect 9398 13880 9404 13892
rect 9456 13880 9462 13932
rect 10965 13923 11023 13929
rect 10965 13889 10977 13923
rect 11011 13889 11023 13923
rect 10965 13883 11023 13889
rect 10980 13852 11008 13883
rect 11146 13880 11152 13932
rect 11204 13880 11210 13932
rect 11256 13920 11284 13948
rect 11701 13923 11759 13929
rect 11701 13920 11713 13923
rect 11256 13892 11713 13920
rect 11701 13889 11713 13892
rect 11747 13889 11759 13923
rect 11701 13883 11759 13889
rect 11330 13852 11336 13864
rect 7668 13824 10916 13852
rect 10980 13824 11336 13852
rect 6043 13821 6055 13824
rect 5997 13815 6055 13821
rect 5077 13787 5135 13793
rect 5077 13753 5089 13787
rect 5123 13784 5135 13787
rect 5718 13784 5724 13796
rect 5123 13756 5724 13784
rect 5123 13753 5135 13756
rect 5077 13747 5135 13753
rect 5718 13744 5724 13756
rect 5776 13744 5782 13796
rect 10888 13784 10916 13824
rect 11330 13812 11336 13824
rect 11388 13812 11394 13864
rect 12084 13852 12112 13951
rect 12912 13929 12940 13960
rect 12897 13923 12955 13929
rect 12897 13889 12909 13923
rect 12943 13889 12955 13923
rect 12897 13883 12955 13889
rect 13541 13923 13599 13929
rect 13541 13889 13553 13923
rect 13587 13920 13599 13923
rect 13630 13920 13636 13932
rect 13587 13892 13636 13920
rect 13587 13889 13599 13892
rect 13541 13883 13599 13889
rect 13630 13880 13636 13892
rect 13688 13880 13694 13932
rect 13740 13920 13768 13960
rect 13808 13957 13820 13991
rect 13854 13988 13866 13991
rect 15396 13988 15424 14019
rect 13854 13960 15424 13988
rect 17880 13988 17908 14019
rect 19886 14016 19892 14068
rect 19944 14056 19950 14068
rect 20717 14059 20775 14065
rect 20717 14056 20729 14059
rect 19944 14028 20729 14056
rect 19944 14016 19950 14028
rect 20717 14025 20729 14028
rect 20763 14025 20775 14059
rect 20717 14019 20775 14025
rect 20809 14059 20867 14065
rect 20809 14025 20821 14059
rect 20855 14056 20867 14059
rect 23385 14059 23443 14065
rect 23385 14056 23397 14059
rect 20855 14028 23397 14056
rect 20855 14025 20867 14028
rect 20809 14019 20867 14025
rect 23385 14025 23397 14028
rect 23431 14056 23443 14059
rect 24213 14059 24271 14065
rect 24213 14056 24225 14059
rect 23431 14028 24225 14056
rect 23431 14025 23443 14028
rect 23385 14019 23443 14025
rect 24213 14025 24225 14028
rect 24259 14025 24271 14059
rect 24213 14019 24271 14025
rect 24305 14059 24363 14065
rect 24305 14025 24317 14059
rect 24351 14056 24363 14059
rect 26602 14056 26608 14068
rect 24351 14028 26608 14056
rect 24351 14025 24363 14028
rect 24305 14019 24363 14025
rect 26602 14016 26608 14028
rect 26660 14016 26666 14068
rect 30190 14016 30196 14068
rect 30248 14016 30254 14068
rect 31297 14059 31355 14065
rect 31297 14025 31309 14059
rect 31343 14056 31355 14059
rect 31386 14056 31392 14068
rect 31343 14028 31392 14056
rect 31343 14025 31355 14028
rect 31297 14019 31355 14025
rect 31386 14016 31392 14028
rect 31444 14016 31450 14068
rect 34425 14059 34483 14065
rect 34425 14025 34437 14059
rect 34471 14056 34483 14059
rect 36265 14059 36323 14065
rect 36265 14056 36277 14059
rect 34471 14028 36277 14056
rect 34471 14025 34483 14028
rect 34425 14019 34483 14025
rect 36265 14025 36277 14028
rect 36311 14025 36323 14059
rect 36265 14019 36323 14025
rect 36357 14059 36415 14065
rect 36357 14025 36369 14059
rect 36403 14056 36415 14059
rect 37461 14059 37519 14065
rect 37461 14056 37473 14059
rect 36403 14028 37473 14056
rect 36403 14025 36415 14028
rect 36357 14019 36415 14025
rect 37461 14025 37473 14028
rect 37507 14025 37519 14059
rect 37461 14019 37519 14025
rect 37826 14016 37832 14068
rect 37884 14016 37890 14068
rect 40126 14016 40132 14068
rect 40184 14016 40190 14068
rect 41325 14059 41383 14065
rect 41325 14025 41337 14059
rect 41371 14056 41383 14059
rect 41414 14056 41420 14068
rect 41371 14028 41420 14056
rect 41371 14025 41383 14028
rect 41325 14019 41383 14025
rect 41414 14016 41420 14028
rect 41472 14016 41478 14068
rect 18754 13991 18812 13997
rect 18754 13988 18766 13991
rect 17880 13960 18766 13988
rect 13854 13957 13866 13960
rect 13808 13951 13866 13957
rect 18754 13957 18766 13960
rect 18800 13957 18812 13991
rect 18754 13951 18812 13957
rect 21910 13948 21916 14000
rect 21968 13988 21974 14000
rect 22250 13991 22308 13997
rect 22250 13988 22262 13991
rect 21968 13960 22262 13988
rect 21968 13948 21974 13960
rect 22250 13957 22262 13960
rect 22296 13957 22308 13991
rect 22250 13951 22308 13957
rect 25498 13948 25504 14000
rect 25556 13988 25562 14000
rect 25556 13960 30236 13988
rect 25556 13948 25562 13960
rect 15102 13920 15108 13932
rect 13740 13892 15108 13920
rect 15102 13880 15108 13892
rect 15160 13880 15166 13932
rect 15562 13880 15568 13932
rect 15620 13880 15626 13932
rect 18049 13923 18107 13929
rect 18049 13889 18061 13923
rect 18095 13920 18107 13923
rect 19334 13920 19340 13932
rect 18095 13892 19340 13920
rect 18095 13889 18107 13892
rect 18049 13883 18107 13889
rect 19334 13880 19340 13892
rect 19392 13880 19398 13932
rect 22005 13923 22063 13929
rect 22005 13889 22017 13923
rect 22051 13920 22063 13923
rect 22094 13920 22100 13932
rect 22051 13892 22100 13920
rect 22051 13889 22063 13892
rect 22005 13883 22063 13889
rect 22094 13880 22100 13892
rect 22152 13880 22158 13932
rect 23842 13880 23848 13932
rect 23900 13920 23906 13932
rect 29546 13920 29552 13932
rect 23900 13892 29552 13920
rect 23900 13880 23906 13892
rect 29546 13880 29552 13892
rect 29604 13880 29610 13932
rect 30006 13880 30012 13932
rect 30064 13880 30070 13932
rect 11440 13824 12112 13852
rect 11440 13784 11468 13824
rect 12618 13812 12624 13864
rect 12676 13852 12682 13864
rect 12713 13855 12771 13861
rect 12713 13852 12725 13855
rect 12676 13824 12725 13852
rect 12676 13812 12682 13824
rect 12713 13821 12725 13824
rect 12759 13821 12771 13855
rect 12713 13815 12771 13821
rect 17862 13812 17868 13864
rect 17920 13852 17926 13864
rect 18509 13855 18567 13861
rect 18509 13852 18521 13855
rect 17920 13824 18521 13852
rect 17920 13812 17926 13824
rect 18509 13821 18521 13824
rect 18555 13821 18567 13855
rect 18509 13815 18567 13821
rect 20990 13812 20996 13864
rect 21048 13852 21054 13864
rect 21048 13824 21128 13852
rect 21048 13812 21054 13824
rect 10888 13756 11468 13784
rect 5813 13719 5871 13725
rect 5813 13685 5825 13719
rect 5859 13716 5871 13719
rect 5994 13716 6000 13728
rect 5859 13688 6000 13716
rect 5859 13685 5871 13688
rect 5813 13679 5871 13685
rect 5994 13676 6000 13688
rect 6052 13676 6058 13728
rect 8754 13676 8760 13728
rect 8812 13676 8818 13728
rect 11057 13719 11115 13725
rect 11057 13685 11069 13719
rect 11103 13716 11115 13719
rect 12069 13719 12127 13725
rect 12069 13716 12081 13719
rect 11103 13688 12081 13716
rect 11103 13685 11115 13688
rect 11057 13679 11115 13685
rect 12069 13685 12081 13688
rect 12115 13685 12127 13719
rect 12069 13679 12127 13685
rect 12710 13676 12716 13728
rect 12768 13716 12774 13728
rect 13081 13719 13139 13725
rect 13081 13716 13093 13719
rect 12768 13688 13093 13716
rect 12768 13676 12774 13688
rect 13081 13685 13093 13688
rect 13127 13685 13139 13719
rect 13081 13679 13139 13685
rect 20346 13676 20352 13728
rect 20404 13676 20410 13728
rect 21100 13716 21128 13824
rect 23014 13812 23020 13864
rect 23072 13852 23078 13864
rect 24489 13855 24547 13861
rect 23072 13824 23888 13852
rect 23072 13812 23078 13824
rect 23860 13793 23888 13824
rect 24489 13821 24501 13855
rect 24535 13821 24547 13855
rect 24489 13815 24547 13821
rect 23845 13787 23903 13793
rect 23845 13753 23857 13787
rect 23891 13753 23903 13787
rect 23845 13747 23903 13753
rect 24504 13784 24532 13815
rect 24854 13812 24860 13864
rect 24912 13852 24918 13864
rect 26142 13852 26148 13864
rect 24912 13824 26148 13852
rect 24912 13812 24918 13824
rect 26142 13812 26148 13824
rect 26200 13852 26206 13864
rect 27798 13852 27804 13864
rect 26200 13824 27804 13852
rect 26200 13812 26206 13824
rect 27798 13812 27804 13824
rect 27856 13812 27862 13864
rect 28994 13812 29000 13864
rect 29052 13852 29058 13864
rect 29730 13852 29736 13864
rect 29052 13824 29736 13852
rect 29052 13812 29058 13824
rect 29730 13812 29736 13824
rect 29788 13852 29794 13864
rect 29825 13855 29883 13861
rect 29825 13852 29837 13855
rect 29788 13824 29837 13852
rect 29788 13812 29794 13824
rect 29825 13821 29837 13824
rect 29871 13821 29883 13855
rect 30208 13852 30236 13960
rect 31202 13948 31208 14000
rect 31260 13988 31266 14000
rect 34606 13988 34612 14000
rect 31260 13960 32536 13988
rect 31260 13948 31266 13960
rect 30282 13880 30288 13932
rect 30340 13920 30346 13932
rect 31481 13923 31539 13929
rect 31481 13920 31493 13923
rect 30340 13892 31493 13920
rect 30340 13880 30346 13892
rect 31481 13889 31493 13892
rect 31527 13889 31539 13923
rect 31481 13883 31539 13889
rect 32398 13852 32404 13864
rect 30208 13824 32404 13852
rect 29825 13815 29883 13821
rect 32398 13812 32404 13824
rect 32456 13812 32462 13864
rect 32508 13852 32536 13960
rect 33060 13960 34612 13988
rect 33060 13929 33088 13960
rect 34606 13948 34612 13960
rect 34664 13948 34670 14000
rect 40034 13988 40040 14000
rect 38764 13960 40040 13988
rect 33045 13923 33103 13929
rect 33045 13889 33057 13923
rect 33091 13889 33103 13923
rect 33301 13923 33359 13929
rect 33301 13920 33313 13923
rect 33045 13883 33103 13889
rect 33152 13892 33313 13920
rect 33152 13852 33180 13892
rect 33301 13889 33313 13892
rect 33347 13889 33359 13923
rect 33301 13883 33359 13889
rect 35437 13923 35495 13929
rect 35437 13889 35449 13923
rect 35483 13920 35495 13923
rect 35483 13892 35940 13920
rect 35483 13889 35495 13892
rect 35437 13883 35495 13889
rect 32508 13824 33180 13852
rect 35268 13824 35848 13852
rect 26786 13784 26792 13796
rect 24504 13756 26792 13784
rect 24504 13716 24532 13756
rect 26786 13744 26792 13756
rect 26844 13744 26850 13796
rect 35268 13793 35296 13824
rect 35253 13787 35311 13793
rect 35253 13753 35265 13787
rect 35299 13753 35311 13787
rect 35253 13747 35311 13753
rect 21100 13688 24532 13716
rect 35820 13716 35848 13824
rect 35912 13793 35940 13892
rect 38378 13880 38384 13932
rect 38436 13920 38442 13932
rect 38764 13929 38792 13960
rect 40034 13948 40040 13960
rect 40092 13948 40098 14000
rect 41690 13948 41696 14000
rect 41748 13948 41754 14000
rect 38749 13923 38807 13929
rect 38749 13920 38761 13923
rect 38436 13892 38761 13920
rect 38436 13880 38442 13892
rect 38749 13889 38761 13892
rect 38795 13889 38807 13923
rect 38749 13883 38807 13889
rect 38838 13880 38844 13932
rect 38896 13920 38902 13932
rect 39005 13923 39063 13929
rect 39005 13920 39017 13923
rect 38896 13892 39017 13920
rect 38896 13880 38902 13892
rect 39005 13889 39017 13892
rect 39051 13889 39063 13923
rect 39005 13883 39063 13889
rect 36262 13812 36268 13864
rect 36320 13852 36326 13864
rect 36446 13852 36452 13864
rect 36320 13824 36452 13852
rect 36320 13812 36326 13824
rect 36446 13812 36452 13824
rect 36504 13812 36510 13864
rect 37918 13812 37924 13864
rect 37976 13812 37982 13864
rect 38105 13855 38163 13861
rect 38105 13821 38117 13855
rect 38151 13852 38163 13855
rect 38194 13852 38200 13864
rect 38151 13824 38200 13852
rect 38151 13821 38163 13824
rect 38105 13815 38163 13821
rect 38194 13812 38200 13824
rect 38252 13812 38258 13864
rect 41782 13812 41788 13864
rect 41840 13812 41846 13864
rect 41877 13855 41935 13861
rect 41877 13821 41889 13855
rect 41923 13821 41935 13855
rect 41877 13815 41935 13821
rect 35897 13787 35955 13793
rect 35897 13753 35909 13787
rect 35943 13753 35955 13787
rect 41892 13784 41920 13815
rect 41966 13784 41972 13796
rect 35897 13747 35955 13753
rect 41386 13756 41972 13784
rect 36630 13716 36636 13728
rect 35820 13688 36636 13716
rect 36630 13676 36636 13688
rect 36688 13676 36694 13728
rect 38930 13676 38936 13728
rect 38988 13716 38994 13728
rect 41386 13716 41414 13756
rect 41966 13744 41972 13756
rect 42024 13744 42030 13796
rect 38988 13688 41414 13716
rect 38988 13676 38994 13688
rect 1104 13626 44896 13648
rect 1104 13574 6423 13626
rect 6475 13574 6487 13626
rect 6539 13574 6551 13626
rect 6603 13574 6615 13626
rect 6667 13574 6679 13626
rect 6731 13574 17370 13626
rect 17422 13574 17434 13626
rect 17486 13574 17498 13626
rect 17550 13574 17562 13626
rect 17614 13574 17626 13626
rect 17678 13574 28317 13626
rect 28369 13574 28381 13626
rect 28433 13574 28445 13626
rect 28497 13574 28509 13626
rect 28561 13574 28573 13626
rect 28625 13574 39264 13626
rect 39316 13574 39328 13626
rect 39380 13574 39392 13626
rect 39444 13574 39456 13626
rect 39508 13574 39520 13626
rect 39572 13574 44896 13626
rect 1104 13552 44896 13574
rect 4154 13512 4160 13524
rect 3436 13484 4160 13512
rect 3436 13317 3464 13484
rect 4154 13472 4160 13484
rect 4212 13472 4218 13524
rect 4982 13472 4988 13524
rect 5040 13512 5046 13524
rect 5353 13515 5411 13521
rect 5353 13512 5365 13515
rect 5040 13484 5365 13512
rect 5040 13472 5046 13484
rect 5353 13481 5365 13484
rect 5399 13512 5411 13515
rect 5997 13515 6055 13521
rect 5997 13512 6009 13515
rect 5399 13484 6009 13512
rect 5399 13481 5411 13484
rect 5353 13475 5411 13481
rect 5997 13481 6009 13484
rect 6043 13512 6055 13515
rect 6822 13512 6828 13524
rect 6043 13484 6828 13512
rect 6043 13481 6055 13484
rect 5997 13475 6055 13481
rect 6822 13472 6828 13484
rect 6880 13472 6886 13524
rect 7009 13515 7067 13521
rect 7009 13481 7021 13515
rect 7055 13512 7067 13515
rect 8754 13512 8760 13524
rect 7055 13484 8760 13512
rect 7055 13481 7067 13484
rect 7009 13475 7067 13481
rect 8754 13472 8760 13484
rect 8812 13472 8818 13524
rect 11054 13472 11060 13524
rect 11112 13512 11118 13524
rect 12529 13515 12587 13521
rect 12529 13512 12541 13515
rect 11112 13484 12541 13512
rect 11112 13472 11118 13484
rect 12529 13481 12541 13484
rect 12575 13481 12587 13515
rect 12529 13475 12587 13481
rect 12618 13472 12624 13524
rect 12676 13512 12682 13524
rect 13633 13515 13691 13521
rect 13633 13512 13645 13515
rect 12676 13484 13645 13512
rect 12676 13472 12682 13484
rect 13633 13481 13645 13484
rect 13679 13481 13691 13515
rect 13633 13475 13691 13481
rect 14645 13515 14703 13521
rect 14645 13481 14657 13515
rect 14691 13512 14703 13515
rect 15289 13515 15347 13521
rect 15289 13512 15301 13515
rect 14691 13484 15301 13512
rect 14691 13481 14703 13484
rect 14645 13475 14703 13481
rect 15289 13481 15301 13484
rect 15335 13481 15347 13515
rect 15289 13475 15347 13481
rect 15473 13515 15531 13521
rect 15473 13481 15485 13515
rect 15519 13512 15531 13515
rect 15562 13512 15568 13524
rect 15519 13484 15568 13512
rect 15519 13481 15531 13484
rect 15473 13475 15531 13481
rect 15562 13472 15568 13484
rect 15620 13472 15626 13524
rect 18506 13472 18512 13524
rect 18564 13512 18570 13524
rect 18877 13515 18935 13521
rect 18877 13512 18889 13515
rect 18564 13484 18889 13512
rect 18564 13472 18570 13484
rect 18877 13481 18889 13484
rect 18923 13481 18935 13515
rect 18877 13475 18935 13481
rect 19334 13472 19340 13524
rect 19392 13512 19398 13524
rect 19429 13515 19487 13521
rect 19429 13512 19441 13515
rect 19392 13484 19441 13512
rect 19392 13472 19398 13484
rect 19429 13481 19441 13484
rect 19475 13481 19487 13515
rect 19429 13475 19487 13481
rect 21637 13515 21695 13521
rect 21637 13481 21649 13515
rect 21683 13512 21695 13515
rect 22186 13512 22192 13524
rect 21683 13484 22192 13512
rect 21683 13481 21695 13484
rect 21637 13475 21695 13481
rect 22186 13472 22192 13484
rect 22244 13472 22250 13524
rect 25498 13512 25504 13524
rect 24780 13484 25504 13512
rect 7193 13447 7251 13453
rect 7193 13413 7205 13447
rect 7239 13444 7251 13447
rect 7374 13444 7380 13456
rect 7239 13416 7380 13444
rect 7239 13413 7251 13416
rect 7193 13407 7251 13413
rect 7374 13404 7380 13416
rect 7432 13404 7438 13456
rect 11238 13404 11244 13456
rect 11296 13404 11302 13456
rect 12342 13444 12348 13456
rect 11440 13416 12348 13444
rect 8021 13379 8079 13385
rect 8021 13376 8033 13379
rect 6886 13348 8033 13376
rect 3421 13311 3479 13317
rect 3421 13277 3433 13311
rect 3467 13277 3479 13311
rect 3421 13271 3479 13277
rect 3973 13311 4031 13317
rect 3973 13277 3985 13311
rect 4019 13308 4031 13311
rect 4062 13308 4068 13320
rect 4019 13280 4068 13308
rect 4019 13277 4031 13280
rect 3973 13271 4031 13277
rect 4062 13268 4068 13280
rect 4120 13268 4126 13320
rect 6641 13311 6699 13317
rect 6641 13277 6653 13311
rect 6687 13308 6699 13311
rect 6886 13308 6914 13348
rect 8021 13345 8033 13348
rect 8067 13345 8079 13379
rect 8021 13339 8079 13345
rect 11146 13336 11152 13388
rect 11204 13376 11210 13388
rect 11440 13376 11468 13416
rect 12342 13404 12348 13416
rect 12400 13404 12406 13456
rect 24780 13444 24808 13484
rect 25498 13472 25504 13484
rect 25556 13472 25562 13524
rect 36354 13472 36360 13524
rect 36412 13512 36418 13524
rect 37737 13515 37795 13521
rect 36412 13484 37320 13512
rect 36412 13472 36418 13484
rect 22204 13416 24808 13444
rect 11204 13348 11468 13376
rect 11204 13336 11210 13348
rect 6687 13280 6914 13308
rect 7745 13311 7803 13317
rect 6687 13277 6699 13280
rect 6641 13271 6699 13277
rect 7745 13277 7757 13311
rect 7791 13277 7803 13311
rect 7745 13271 7803 13277
rect 7837 13311 7895 13317
rect 7837 13277 7849 13311
rect 7883 13308 7895 13311
rect 8202 13308 8208 13320
rect 7883 13280 8208 13308
rect 7883 13277 7895 13280
rect 7837 13271 7895 13277
rect 4218 13243 4276 13249
rect 4218 13240 4230 13243
rect 3252 13212 4230 13240
rect 3252 13181 3280 13212
rect 4218 13209 4230 13212
rect 4264 13209 4276 13243
rect 4218 13203 4276 13209
rect 5810 13200 5816 13252
rect 5868 13200 5874 13252
rect 5994 13200 6000 13252
rect 6052 13249 6058 13252
rect 6052 13243 6071 13249
rect 6059 13240 6071 13243
rect 6656 13240 6684 13271
rect 6059 13212 6684 13240
rect 7009 13243 7067 13249
rect 6059 13209 6071 13212
rect 6052 13203 6071 13209
rect 7009 13209 7021 13243
rect 7055 13240 7067 13243
rect 7098 13240 7104 13252
rect 7055 13212 7104 13240
rect 7055 13209 7067 13212
rect 7009 13203 7067 13209
rect 6052 13200 6058 13203
rect 7098 13200 7104 13212
rect 7156 13200 7162 13252
rect 7760 13240 7788 13271
rect 8202 13268 8208 13280
rect 8260 13268 8266 13320
rect 11241 13311 11299 13317
rect 11241 13277 11253 13311
rect 11287 13308 11299 13311
rect 11330 13308 11336 13320
rect 11287 13280 11336 13308
rect 11287 13277 11299 13280
rect 11241 13271 11299 13277
rect 11330 13268 11336 13280
rect 11388 13268 11394 13320
rect 11440 13317 11468 13348
rect 11514 13336 11520 13388
rect 11572 13376 11578 13388
rect 12621 13379 12679 13385
rect 12621 13376 12633 13379
rect 11572 13348 12633 13376
rect 11572 13336 11578 13348
rect 12621 13345 12633 13348
rect 12667 13345 12679 13379
rect 12621 13339 12679 13345
rect 19978 13336 19984 13388
rect 20036 13376 20042 13388
rect 22204 13385 22232 13416
rect 22189 13379 22247 13385
rect 22189 13376 22201 13379
rect 20036 13348 22201 13376
rect 20036 13336 20042 13348
rect 22189 13345 22201 13348
rect 22235 13345 22247 13379
rect 22189 13339 22247 13345
rect 23937 13379 23995 13385
rect 23937 13345 23949 13379
rect 23983 13376 23995 13379
rect 24670 13376 24676 13388
rect 23983 13348 24676 13376
rect 23983 13345 23995 13348
rect 23937 13339 23995 13345
rect 24670 13336 24676 13348
rect 24728 13336 24734 13388
rect 11425 13311 11483 13317
rect 11425 13277 11437 13311
rect 11471 13277 11483 13311
rect 11425 13271 11483 13277
rect 12069 13311 12127 13317
rect 12069 13277 12081 13311
rect 12115 13308 12127 13311
rect 12710 13308 12716 13320
rect 12115 13280 12716 13308
rect 12115 13277 12127 13280
rect 12069 13271 12127 13277
rect 12710 13268 12716 13280
rect 12768 13268 12774 13320
rect 12802 13268 12808 13320
rect 12860 13268 12866 13320
rect 13541 13311 13599 13317
rect 13541 13277 13553 13311
rect 13587 13277 13599 13311
rect 13541 13271 13599 13277
rect 8478 13240 8484 13252
rect 7760 13212 8484 13240
rect 8478 13200 8484 13212
rect 8536 13200 8542 13252
rect 12526 13200 12532 13252
rect 12584 13200 12590 13252
rect 13078 13240 13084 13252
rect 12820 13212 13084 13240
rect 3237 13175 3295 13181
rect 3237 13141 3249 13175
rect 3283 13141 3295 13175
rect 3237 13135 3295 13141
rect 4338 13132 4344 13184
rect 4396 13172 4402 13184
rect 6181 13175 6239 13181
rect 6181 13172 6193 13175
rect 4396 13144 6193 13172
rect 4396 13132 4402 13144
rect 6181 13141 6193 13144
rect 6227 13172 6239 13175
rect 6546 13172 6552 13184
rect 6227 13144 6552 13172
rect 6227 13141 6239 13144
rect 6181 13135 6239 13141
rect 6546 13132 6552 13144
rect 6604 13132 6610 13184
rect 11885 13175 11943 13181
rect 11885 13141 11897 13175
rect 11931 13172 11943 13175
rect 12820 13172 12848 13212
rect 13078 13200 13084 13212
rect 13136 13200 13142 13252
rect 13556 13240 13584 13271
rect 14274 13268 14280 13320
rect 14332 13268 14338 13320
rect 14458 13268 14464 13320
rect 14516 13268 14522 13320
rect 17497 13311 17555 13317
rect 17497 13277 17509 13311
rect 17543 13308 17555 13311
rect 19889 13311 19947 13317
rect 17543 13280 17908 13308
rect 17543 13277 17555 13280
rect 17497 13271 17555 13277
rect 14476 13240 14504 13268
rect 17880 13252 17908 13280
rect 19889 13277 19901 13311
rect 19935 13308 19947 13311
rect 20346 13308 20352 13320
rect 19935 13280 20352 13308
rect 19935 13277 19947 13280
rect 19889 13271 19947 13277
rect 20346 13268 20352 13280
rect 20404 13268 20410 13320
rect 22097 13311 22155 13317
rect 22097 13277 22109 13311
rect 22143 13308 22155 13311
rect 23014 13308 23020 13320
rect 22143 13280 23020 13308
rect 22143 13277 22155 13280
rect 22097 13271 22155 13277
rect 23014 13268 23020 13280
rect 23072 13268 23078 13320
rect 23566 13268 23572 13320
rect 23624 13308 23630 13320
rect 23661 13311 23719 13317
rect 23661 13308 23673 13311
rect 23624 13280 23673 13308
rect 23624 13268 23630 13280
rect 23661 13277 23673 13280
rect 23707 13277 23719 13311
rect 23661 13271 23719 13277
rect 24765 13311 24823 13317
rect 24765 13277 24777 13311
rect 24811 13308 24823 13311
rect 24854 13308 24860 13320
rect 24811 13280 24860 13308
rect 24811 13277 24823 13280
rect 24765 13271 24823 13277
rect 24854 13268 24860 13280
rect 24912 13268 24918 13320
rect 27890 13308 27896 13320
rect 26206 13280 27896 13308
rect 13556 13212 14504 13240
rect 15102 13200 15108 13252
rect 15160 13200 15166 13252
rect 15286 13200 15292 13252
rect 15344 13249 15350 13252
rect 17770 13249 17776 13252
rect 15344 13243 15363 13249
rect 15351 13209 15363 13243
rect 15344 13203 15363 13209
rect 17764 13203 17776 13249
rect 15344 13200 15350 13203
rect 17770 13200 17776 13203
rect 17828 13200 17834 13252
rect 17862 13200 17868 13252
rect 17920 13200 17926 13252
rect 25032 13243 25090 13249
rect 25032 13209 25044 13243
rect 25078 13240 25090 13243
rect 26206 13240 26234 13280
rect 27890 13268 27896 13280
rect 27948 13268 27954 13320
rect 28166 13268 28172 13320
rect 28224 13268 28230 13320
rect 28813 13311 28871 13317
rect 28813 13277 28825 13311
rect 28859 13277 28871 13311
rect 28813 13271 28871 13277
rect 25078 13212 26234 13240
rect 27709 13243 27767 13249
rect 25078 13209 25090 13212
rect 25032 13203 25090 13209
rect 27709 13209 27721 13243
rect 27755 13240 27767 13243
rect 28828 13240 28856 13271
rect 28902 13268 28908 13320
rect 28960 13308 28966 13320
rect 30745 13311 30803 13317
rect 30745 13308 30757 13311
rect 28960 13280 30757 13308
rect 28960 13268 28966 13280
rect 30745 13277 30757 13280
rect 30791 13308 30803 13311
rect 30834 13308 30840 13320
rect 30791 13280 30840 13308
rect 30791 13277 30803 13280
rect 30745 13271 30803 13277
rect 30834 13268 30840 13280
rect 30892 13268 30898 13320
rect 32766 13268 32772 13320
rect 32824 13268 32830 13320
rect 36372 13317 36400 13472
rect 37292 13444 37320 13484
rect 37737 13481 37749 13515
rect 37783 13512 37795 13515
rect 37826 13512 37832 13524
rect 37783 13484 37832 13512
rect 37783 13481 37795 13484
rect 37737 13475 37795 13481
rect 37826 13472 37832 13484
rect 37884 13472 37890 13524
rect 38378 13444 38384 13456
rect 37292 13416 38384 13444
rect 38378 13404 38384 13416
rect 38436 13404 38442 13456
rect 36630 13317 36636 13320
rect 36357 13311 36415 13317
rect 36357 13277 36369 13311
rect 36403 13277 36415 13311
rect 36357 13271 36415 13277
rect 36613 13311 36636 13317
rect 36613 13277 36625 13311
rect 36613 13271 36636 13277
rect 36630 13268 36636 13271
rect 36688 13268 36694 13320
rect 38381 13311 38439 13317
rect 38381 13277 38393 13311
rect 38427 13277 38439 13311
rect 38381 13271 38439 13277
rect 27755 13212 28856 13240
rect 31012 13243 31070 13249
rect 27755 13209 27767 13212
rect 27709 13203 27767 13209
rect 31012 13209 31024 13243
rect 31058 13240 31070 13243
rect 31058 13212 32628 13240
rect 31058 13209 31070 13212
rect 31012 13203 31070 13209
rect 11931 13144 12848 13172
rect 11931 13141 11943 13144
rect 11885 13135 11943 13141
rect 12986 13132 12992 13184
rect 13044 13132 13050 13184
rect 18874 13132 18880 13184
rect 18932 13172 18938 13184
rect 19797 13175 19855 13181
rect 19797 13172 19809 13175
rect 18932 13144 19809 13172
rect 18932 13132 18938 13144
rect 19797 13141 19809 13144
rect 19843 13141 19855 13175
rect 19797 13135 19855 13141
rect 22002 13132 22008 13184
rect 22060 13132 22066 13184
rect 22646 13132 22652 13184
rect 22704 13172 22710 13184
rect 23293 13175 23351 13181
rect 23293 13172 23305 13175
rect 22704 13144 23305 13172
rect 22704 13132 22710 13144
rect 23293 13141 23305 13144
rect 23339 13141 23351 13175
rect 23293 13135 23351 13141
rect 23753 13175 23811 13181
rect 23753 13141 23765 13175
rect 23799 13172 23811 13175
rect 26145 13175 26203 13181
rect 26145 13172 26157 13175
rect 23799 13144 26157 13172
rect 23799 13141 23811 13144
rect 23753 13135 23811 13141
rect 26145 13141 26157 13144
rect 26191 13141 26203 13175
rect 26145 13135 26203 13141
rect 28074 13132 28080 13184
rect 28132 13132 28138 13184
rect 28258 13132 28264 13184
rect 28316 13172 28322 13184
rect 28629 13175 28687 13181
rect 28629 13172 28641 13175
rect 28316 13144 28641 13172
rect 28316 13132 28322 13144
rect 28629 13141 28641 13144
rect 28675 13141 28687 13175
rect 28629 13135 28687 13141
rect 31478 13132 31484 13184
rect 31536 13172 31542 13184
rect 32600 13181 32628 13212
rect 37090 13200 37096 13252
rect 37148 13240 37154 13252
rect 38396 13240 38424 13271
rect 37148 13212 38424 13240
rect 37148 13200 37154 13212
rect 32125 13175 32183 13181
rect 32125 13172 32137 13175
rect 31536 13144 32137 13172
rect 31536 13132 31542 13144
rect 32125 13141 32137 13144
rect 32171 13141 32183 13175
rect 32125 13135 32183 13141
rect 32585 13175 32643 13181
rect 32585 13141 32597 13175
rect 32631 13141 32643 13175
rect 32585 13135 32643 13141
rect 38102 13132 38108 13184
rect 38160 13172 38166 13184
rect 38197 13175 38255 13181
rect 38197 13172 38209 13175
rect 38160 13144 38209 13172
rect 38160 13132 38166 13144
rect 38197 13141 38209 13144
rect 38243 13141 38255 13175
rect 38197 13135 38255 13141
rect 1104 13082 45051 13104
rect 1104 13030 11896 13082
rect 11948 13030 11960 13082
rect 12012 13030 12024 13082
rect 12076 13030 12088 13082
rect 12140 13030 12152 13082
rect 12204 13030 22843 13082
rect 22895 13030 22907 13082
rect 22959 13030 22971 13082
rect 23023 13030 23035 13082
rect 23087 13030 23099 13082
rect 23151 13030 33790 13082
rect 33842 13030 33854 13082
rect 33906 13030 33918 13082
rect 33970 13030 33982 13082
rect 34034 13030 34046 13082
rect 34098 13030 44737 13082
rect 44789 13030 44801 13082
rect 44853 13030 44865 13082
rect 44917 13030 44929 13082
rect 44981 13030 44993 13082
rect 45045 13030 45051 13082
rect 1104 13008 45051 13030
rect 3050 12928 3056 12980
rect 3108 12968 3114 12980
rect 3513 12971 3571 12977
rect 3513 12968 3525 12971
rect 3108 12940 3525 12968
rect 3108 12928 3114 12940
rect 3513 12937 3525 12940
rect 3559 12937 3571 12971
rect 3513 12931 3571 12937
rect 4522 12928 4528 12980
rect 4580 12968 4586 12980
rect 5718 12968 5724 12980
rect 4580 12940 5724 12968
rect 4580 12928 4586 12940
rect 5718 12928 5724 12940
rect 5776 12928 5782 12980
rect 11054 12928 11060 12980
rect 11112 12928 11118 12980
rect 12529 12971 12587 12977
rect 11256 12940 12296 12968
rect 4890 12860 4896 12912
rect 4948 12900 4954 12912
rect 5258 12900 5264 12912
rect 4948 12872 5264 12900
rect 4948 12860 4954 12872
rect 5258 12860 5264 12872
rect 5316 12900 5322 12912
rect 5629 12903 5687 12909
rect 5629 12900 5641 12903
rect 5316 12872 5641 12900
rect 5316 12860 5322 12872
rect 5629 12869 5641 12872
rect 5675 12869 5687 12903
rect 5629 12863 5687 12869
rect 5845 12903 5903 12909
rect 5845 12869 5857 12903
rect 5891 12900 5903 12903
rect 6917 12903 6975 12909
rect 6917 12900 6929 12903
rect 5891 12872 6929 12900
rect 5891 12869 5903 12872
rect 5845 12863 5903 12869
rect 6917 12869 6929 12872
rect 6963 12869 6975 12903
rect 6917 12863 6975 12869
rect 9493 12903 9551 12909
rect 9493 12869 9505 12903
rect 9539 12900 9551 12903
rect 11256 12900 11284 12940
rect 9539 12872 11284 12900
rect 9539 12869 9551 12872
rect 9493 12863 9551 12869
rect 11330 12860 11336 12912
rect 11388 12900 11394 12912
rect 12268 12909 12296 12940
rect 12529 12937 12541 12971
rect 12575 12968 12587 12971
rect 12802 12968 12808 12980
rect 12575 12940 12808 12968
rect 12575 12937 12587 12940
rect 12529 12931 12587 12937
rect 12802 12928 12808 12940
rect 12860 12928 12866 12980
rect 14369 12971 14427 12977
rect 14369 12937 14381 12971
rect 14415 12968 14427 12971
rect 14458 12968 14464 12980
rect 14415 12940 14464 12968
rect 14415 12937 14427 12940
rect 14369 12931 14427 12937
rect 14458 12928 14464 12940
rect 14516 12928 14522 12980
rect 18874 12928 18880 12980
rect 18932 12928 18938 12980
rect 24854 12968 24860 12980
rect 23216 12940 24860 12968
rect 12161 12903 12219 12909
rect 12161 12900 12173 12903
rect 11388 12872 12173 12900
rect 11388 12860 11394 12872
rect 12161 12869 12173 12872
rect 12207 12869 12219 12903
rect 12161 12863 12219 12869
rect 12253 12903 12311 12909
rect 12253 12869 12265 12903
rect 12299 12900 12311 12903
rect 12434 12900 12440 12912
rect 12299 12872 12440 12900
rect 12299 12869 12311 12872
rect 12253 12863 12311 12869
rect 12434 12860 12440 12872
rect 12492 12860 12498 12912
rect 13722 12900 13728 12912
rect 13004 12872 13728 12900
rect 3329 12835 3387 12841
rect 3329 12801 3341 12835
rect 3375 12832 3387 12835
rect 3418 12832 3424 12844
rect 3375 12804 3424 12832
rect 3375 12801 3387 12804
rect 3329 12795 3387 12801
rect 3418 12792 3424 12804
rect 3476 12792 3482 12844
rect 4338 12792 4344 12844
rect 4396 12792 4402 12844
rect 4525 12835 4583 12841
rect 4525 12801 4537 12835
rect 4571 12801 4583 12835
rect 4525 12795 4583 12801
rect 5169 12835 5227 12841
rect 5169 12801 5181 12835
rect 5215 12832 5227 12835
rect 5215 12804 6040 12832
rect 5215 12801 5227 12804
rect 5169 12795 5227 12801
rect 3145 12767 3203 12773
rect 3145 12733 3157 12767
rect 3191 12764 3203 12767
rect 4430 12764 4436 12776
rect 3191 12736 4436 12764
rect 3191 12733 3203 12736
rect 3145 12727 3203 12733
rect 4430 12724 4436 12736
rect 4488 12724 4494 12776
rect 4540 12696 4568 12795
rect 6012 12705 6040 12804
rect 6546 12792 6552 12844
rect 6604 12792 6610 12844
rect 6733 12835 6791 12841
rect 6733 12801 6745 12835
rect 6779 12801 6791 12835
rect 6733 12795 6791 12801
rect 5997 12699 6055 12705
rect 4540 12668 5948 12696
rect 4985 12631 5043 12637
rect 4985 12597 4997 12631
rect 5031 12628 5043 12631
rect 5718 12628 5724 12640
rect 5031 12600 5724 12628
rect 5031 12597 5043 12600
rect 4985 12591 5043 12597
rect 5718 12588 5724 12600
rect 5776 12588 5782 12640
rect 5810 12588 5816 12640
rect 5868 12588 5874 12640
rect 5920 12628 5948 12668
rect 5997 12665 6009 12699
rect 6043 12665 6055 12699
rect 5997 12659 6055 12665
rect 6748 12628 6776 12795
rect 6822 12792 6828 12844
rect 6880 12832 6886 12844
rect 7377 12835 7435 12841
rect 7377 12832 7389 12835
rect 6880 12804 7389 12832
rect 6880 12792 6886 12804
rect 7377 12801 7389 12804
rect 7423 12801 7435 12835
rect 7377 12795 7435 12801
rect 9398 12792 9404 12844
rect 9456 12792 9462 12844
rect 10965 12835 11023 12841
rect 10965 12801 10977 12835
rect 11011 12832 11023 12835
rect 11054 12832 11060 12844
rect 11011 12804 11060 12832
rect 11011 12801 11023 12804
rect 10965 12795 11023 12801
rect 11054 12792 11060 12804
rect 11112 12792 11118 12844
rect 11146 12792 11152 12844
rect 11204 12792 11210 12844
rect 11238 12792 11244 12844
rect 11296 12832 11302 12844
rect 11885 12835 11943 12841
rect 11885 12832 11897 12835
rect 11296 12804 11897 12832
rect 11296 12792 11302 12804
rect 11885 12801 11897 12804
rect 11931 12801 11943 12835
rect 11885 12795 11943 12801
rect 11978 12835 12036 12841
rect 11978 12801 11990 12835
rect 12024 12801 12036 12835
rect 11978 12795 12036 12801
rect 11992 12764 12020 12795
rect 12342 12792 12348 12844
rect 12400 12841 12406 12844
rect 13004 12841 13032 12872
rect 13722 12860 13728 12872
rect 13780 12860 13786 12912
rect 17862 12900 17868 12912
rect 17512 12872 17868 12900
rect 12400 12795 12408 12841
rect 12989 12835 13047 12841
rect 12989 12801 13001 12835
rect 13035 12801 13047 12835
rect 12989 12795 13047 12801
rect 12400 12792 12406 12795
rect 13078 12792 13084 12844
rect 13136 12832 13142 12844
rect 13245 12835 13303 12841
rect 13245 12832 13257 12835
rect 13136 12804 13257 12832
rect 13136 12792 13142 12804
rect 13245 12801 13257 12804
rect 13291 12801 13303 12835
rect 13245 12795 13303 12801
rect 14274 12792 14280 12844
rect 14332 12832 14338 12844
rect 17512 12841 17540 12872
rect 17862 12860 17868 12872
rect 17920 12900 17926 12912
rect 20714 12900 20720 12912
rect 17920 12872 20720 12900
rect 17920 12860 17926 12872
rect 14829 12835 14887 12841
rect 14829 12832 14841 12835
rect 14332 12804 14841 12832
rect 14332 12792 14338 12804
rect 14829 12801 14841 12804
rect 14875 12801 14887 12835
rect 14829 12795 14887 12801
rect 17497 12835 17555 12841
rect 17497 12801 17509 12835
rect 17543 12801 17555 12835
rect 17497 12795 17555 12801
rect 17764 12835 17822 12841
rect 17764 12801 17776 12835
rect 17810 12832 17822 12835
rect 18046 12832 18052 12844
rect 17810 12804 18052 12832
rect 17810 12801 17822 12804
rect 17764 12795 17822 12801
rect 18046 12792 18052 12804
rect 18104 12792 18110 12844
rect 19352 12841 19380 12872
rect 20714 12860 20720 12872
rect 20772 12860 20778 12912
rect 19337 12835 19395 12841
rect 19337 12801 19349 12835
rect 19383 12801 19395 12835
rect 19337 12795 19395 12801
rect 19426 12792 19432 12844
rect 19484 12832 19490 12844
rect 19593 12835 19651 12841
rect 19593 12832 19605 12835
rect 19484 12804 19605 12832
rect 19484 12792 19490 12804
rect 19593 12801 19605 12804
rect 19639 12801 19651 12835
rect 19593 12795 19651 12801
rect 22738 12792 22744 12844
rect 22796 12792 22802 12844
rect 23216 12841 23244 12940
rect 24854 12928 24860 12940
rect 24912 12928 24918 12980
rect 28902 12968 28908 12980
rect 28000 12940 28908 12968
rect 23201 12835 23259 12841
rect 23201 12801 23213 12835
rect 23247 12801 23259 12835
rect 23201 12795 23259 12801
rect 24578 12792 24584 12844
rect 24636 12792 24642 12844
rect 26605 12835 26663 12841
rect 26605 12801 26617 12835
rect 26651 12801 26663 12835
rect 26605 12795 26663 12801
rect 23477 12767 23535 12773
rect 23477 12764 23489 12767
rect 10796 12736 12020 12764
rect 22572 12736 23489 12764
rect 10796 12708 10824 12736
rect 7469 12699 7527 12705
rect 7469 12665 7481 12699
rect 7515 12696 7527 12699
rect 10778 12696 10784 12708
rect 7515 12668 10784 12696
rect 7515 12665 7527 12668
rect 7469 12659 7527 12665
rect 10778 12656 10784 12668
rect 10836 12656 10842 12708
rect 20717 12699 20775 12705
rect 20717 12665 20729 12699
rect 20763 12696 20775 12699
rect 22002 12696 22008 12708
rect 20763 12668 22008 12696
rect 20763 12665 20775 12668
rect 20717 12659 20775 12665
rect 22002 12656 22008 12668
rect 22060 12656 22066 12708
rect 22572 12705 22600 12736
rect 23477 12733 23489 12736
rect 23523 12733 23535 12767
rect 26620 12764 26648 12795
rect 27154 12792 27160 12844
rect 27212 12792 27218 12844
rect 28000 12841 28028 12940
rect 28902 12928 28908 12940
rect 28960 12928 28966 12980
rect 30193 12971 30251 12977
rect 30193 12937 30205 12971
rect 30239 12937 30251 12971
rect 30193 12931 30251 12937
rect 28258 12860 28264 12912
rect 28316 12860 28322 12912
rect 30208 12900 30236 12931
rect 31478 12928 31484 12980
rect 31536 12928 31542 12980
rect 38194 12928 38200 12980
rect 38252 12968 38258 12980
rect 38252 12940 40448 12968
rect 38252 12928 38258 12940
rect 29486 12872 30236 12900
rect 31297 12903 31355 12909
rect 31297 12869 31309 12903
rect 31343 12900 31355 12903
rect 32030 12900 32036 12912
rect 31343 12872 32036 12900
rect 31343 12869 31355 12872
rect 31297 12863 31355 12869
rect 32030 12860 32036 12872
rect 32088 12860 32094 12912
rect 38930 12900 38936 12912
rect 32600 12872 38936 12900
rect 27985 12835 28043 12841
rect 27985 12801 27997 12835
rect 28031 12801 28043 12835
rect 27985 12795 28043 12801
rect 30374 12792 30380 12844
rect 30432 12792 30438 12844
rect 31202 12792 31208 12844
rect 31260 12832 31266 12844
rect 32493 12835 32551 12841
rect 32493 12832 32505 12835
rect 31260 12804 32505 12832
rect 31260 12792 31266 12804
rect 32493 12801 32505 12804
rect 32539 12801 32551 12835
rect 32493 12795 32551 12801
rect 27249 12767 27307 12773
rect 27249 12764 27261 12767
rect 26620 12736 27261 12764
rect 23477 12727 23535 12733
rect 27249 12733 27261 12736
rect 27295 12733 27307 12767
rect 27249 12727 27307 12733
rect 31478 12724 31484 12776
rect 31536 12764 31542 12776
rect 31573 12767 31631 12773
rect 31573 12764 31585 12767
rect 31536 12736 31585 12764
rect 31536 12724 31542 12736
rect 31573 12733 31585 12736
rect 31619 12733 31631 12767
rect 32306 12764 32312 12776
rect 31573 12727 31631 12733
rect 31726 12736 32312 12764
rect 22557 12699 22615 12705
rect 22557 12665 22569 12699
rect 22603 12665 22615 12699
rect 22557 12659 22615 12665
rect 29733 12699 29791 12705
rect 29733 12665 29745 12699
rect 29779 12696 29791 12699
rect 31726 12696 31754 12736
rect 32306 12724 32312 12736
rect 32364 12724 32370 12776
rect 29779 12668 31754 12696
rect 29779 12665 29791 12668
rect 29733 12659 29791 12665
rect 6914 12628 6920 12640
rect 5920 12600 6920 12628
rect 6914 12588 6920 12600
rect 6972 12588 6978 12640
rect 14826 12588 14832 12640
rect 14884 12628 14890 12640
rect 14921 12631 14979 12637
rect 14921 12628 14933 12631
rect 14884 12600 14933 12628
rect 14884 12588 14890 12600
rect 14921 12597 14933 12600
rect 14967 12597 14979 12631
rect 14921 12591 14979 12597
rect 24946 12588 24952 12640
rect 25004 12588 25010 12640
rect 26421 12631 26479 12637
rect 26421 12597 26433 12631
rect 26467 12628 26479 12631
rect 26878 12628 26884 12640
rect 26467 12600 26884 12628
rect 26467 12597 26479 12600
rect 26421 12591 26479 12597
rect 26878 12588 26884 12600
rect 26936 12588 26942 12640
rect 28074 12588 28080 12640
rect 28132 12628 28138 12640
rect 29748 12628 29776 12659
rect 28132 12600 29776 12628
rect 28132 12588 28138 12600
rect 31018 12588 31024 12640
rect 31076 12588 31082 12640
rect 31478 12588 31484 12640
rect 31536 12628 31542 12640
rect 32600 12628 32628 12872
rect 38930 12860 38936 12872
rect 38988 12860 38994 12912
rect 40034 12900 40040 12912
rect 39882 12872 40040 12900
rect 40034 12860 40040 12872
rect 40092 12860 40098 12912
rect 40420 12909 40448 12940
rect 40405 12903 40463 12909
rect 40405 12869 40417 12903
rect 40451 12869 40463 12903
rect 40405 12863 40463 12869
rect 33318 12792 33324 12844
rect 33376 12792 33382 12844
rect 36078 12792 36084 12844
rect 36136 12792 36142 12844
rect 36173 12835 36231 12841
rect 36173 12801 36185 12835
rect 36219 12832 36231 12835
rect 36817 12835 36875 12841
rect 36817 12832 36829 12835
rect 36219 12804 36829 12832
rect 36219 12801 36231 12804
rect 36173 12795 36231 12801
rect 36817 12801 36829 12804
rect 36863 12801 36875 12835
rect 36817 12795 36875 12801
rect 37642 12792 37648 12844
rect 37700 12792 37706 12844
rect 38378 12792 38384 12844
rect 38436 12792 38442 12844
rect 41046 12792 41052 12844
rect 41104 12792 41110 12844
rect 38654 12724 38660 12776
rect 38712 12724 38718 12776
rect 32677 12699 32735 12705
rect 32677 12665 32689 12699
rect 32723 12696 32735 12699
rect 34330 12696 34336 12708
rect 32723 12668 34336 12696
rect 32723 12665 32735 12668
rect 32677 12659 32735 12665
rect 34330 12656 34336 12668
rect 34388 12656 34394 12708
rect 31536 12600 32628 12628
rect 31536 12588 31542 12600
rect 33134 12588 33140 12640
rect 33192 12588 33198 12640
rect 36538 12588 36544 12640
rect 36596 12628 36602 12640
rect 36633 12631 36691 12637
rect 36633 12628 36645 12631
rect 36596 12600 36645 12628
rect 36596 12588 36602 12600
rect 36633 12597 36645 12600
rect 36679 12597 36691 12631
rect 36633 12591 36691 12597
rect 37458 12588 37464 12640
rect 37516 12588 37522 12640
rect 40865 12631 40923 12637
rect 40865 12597 40877 12631
rect 40911 12628 40923 12631
rect 40954 12628 40960 12640
rect 40911 12600 40960 12628
rect 40911 12597 40923 12600
rect 40865 12591 40923 12597
rect 40954 12588 40960 12600
rect 41012 12588 41018 12640
rect 44361 12631 44419 12637
rect 44361 12597 44373 12631
rect 44407 12628 44419 12631
rect 45002 12628 45008 12640
rect 44407 12600 45008 12628
rect 44407 12597 44419 12600
rect 44361 12591 44419 12597
rect 45002 12588 45008 12600
rect 45060 12588 45066 12640
rect 1104 12538 44896 12560
rect 1104 12486 6423 12538
rect 6475 12486 6487 12538
rect 6539 12486 6551 12538
rect 6603 12486 6615 12538
rect 6667 12486 6679 12538
rect 6731 12486 17370 12538
rect 17422 12486 17434 12538
rect 17486 12486 17498 12538
rect 17550 12486 17562 12538
rect 17614 12486 17626 12538
rect 17678 12486 28317 12538
rect 28369 12486 28381 12538
rect 28433 12486 28445 12538
rect 28497 12486 28509 12538
rect 28561 12486 28573 12538
rect 28625 12486 39264 12538
rect 39316 12486 39328 12538
rect 39380 12486 39392 12538
rect 39444 12486 39456 12538
rect 39508 12486 39520 12538
rect 39572 12486 44896 12538
rect 1104 12464 44896 12486
rect 6914 12384 6920 12436
rect 6972 12384 6978 12436
rect 10597 12427 10655 12433
rect 10597 12393 10609 12427
rect 10643 12424 10655 12427
rect 11514 12424 11520 12436
rect 10643 12396 11520 12424
rect 10643 12393 10655 12396
rect 10597 12387 10655 12393
rect 11514 12384 11520 12396
rect 11572 12384 11578 12436
rect 11701 12427 11759 12433
rect 11701 12393 11713 12427
rect 11747 12424 11759 12427
rect 12526 12424 12532 12436
rect 11747 12396 12532 12424
rect 11747 12393 11759 12396
rect 11701 12387 11759 12393
rect 12526 12384 12532 12396
rect 12584 12384 12590 12436
rect 12986 12384 12992 12436
rect 13044 12424 13050 12436
rect 13265 12427 13323 12433
rect 13265 12424 13277 12427
rect 13044 12396 13277 12424
rect 13044 12384 13050 12396
rect 13265 12393 13277 12396
rect 13311 12393 13323 12427
rect 13265 12387 13323 12393
rect 13354 12384 13360 12436
rect 13412 12424 13418 12436
rect 14277 12427 14335 12433
rect 14277 12424 14289 12427
rect 13412 12396 14289 12424
rect 13412 12384 13418 12396
rect 14277 12393 14289 12396
rect 14323 12393 14335 12427
rect 14277 12387 14335 12393
rect 15102 12384 15108 12436
rect 15160 12424 15166 12436
rect 16669 12427 16727 12433
rect 16669 12424 16681 12427
rect 15160 12396 16681 12424
rect 15160 12384 15166 12396
rect 16669 12393 16681 12396
rect 16715 12393 16727 12427
rect 16669 12387 16727 12393
rect 17770 12384 17776 12436
rect 17828 12424 17834 12436
rect 17865 12427 17923 12433
rect 17865 12424 17877 12427
rect 17828 12396 17877 12424
rect 17828 12384 17834 12396
rect 17865 12393 17877 12396
rect 17911 12393 17923 12427
rect 17865 12387 17923 12393
rect 20622 12384 20628 12436
rect 20680 12424 20686 12436
rect 22462 12424 22468 12436
rect 20680 12396 22468 12424
rect 20680 12384 20686 12396
rect 22462 12384 22468 12396
rect 22520 12384 22526 12436
rect 22738 12384 22744 12436
rect 22796 12424 22802 12436
rect 23293 12427 23351 12433
rect 23293 12424 23305 12427
rect 22796 12396 23305 12424
rect 22796 12384 22802 12396
rect 23293 12393 23305 12396
rect 23339 12393 23351 12427
rect 23293 12387 23351 12393
rect 24578 12384 24584 12436
rect 24636 12384 24642 12436
rect 24688 12396 27476 12424
rect 4522 12356 4528 12368
rect 3988 12328 4528 12356
rect 3988 12229 4016 12328
rect 4522 12316 4528 12328
rect 4580 12316 4586 12368
rect 10137 12359 10195 12365
rect 10137 12325 10149 12359
rect 10183 12356 10195 12359
rect 13173 12359 13231 12365
rect 13173 12356 13185 12359
rect 10183 12328 13185 12356
rect 10183 12325 10195 12328
rect 10137 12319 10195 12325
rect 13173 12325 13185 12328
rect 13219 12325 13231 12359
rect 14826 12356 14832 12368
rect 13173 12319 13231 12325
rect 13280 12328 14832 12356
rect 4062 12248 4068 12300
rect 4120 12288 4126 12300
rect 4120 12260 5580 12288
rect 4120 12248 4126 12260
rect 5552 12232 5580 12260
rect 9858 12248 9864 12300
rect 9916 12248 9922 12300
rect 10778 12248 10784 12300
rect 10836 12248 10842 12300
rect 10962 12248 10968 12300
rect 11020 12288 11026 12300
rect 11885 12291 11943 12297
rect 11885 12288 11897 12291
rect 11020 12260 11897 12288
rect 11020 12248 11026 12260
rect 11885 12257 11897 12260
rect 11931 12288 11943 12291
rect 12253 12291 12311 12297
rect 11931 12260 12204 12288
rect 11931 12257 11943 12260
rect 11885 12251 11943 12257
rect 3421 12223 3479 12229
rect 3421 12189 3433 12223
rect 3467 12189 3479 12223
rect 3421 12183 3479 12189
rect 3973 12223 4031 12229
rect 3973 12189 3985 12223
rect 4019 12189 4031 12223
rect 3973 12183 4031 12189
rect 4157 12223 4215 12229
rect 4157 12189 4169 12223
rect 4203 12220 4215 12223
rect 4338 12220 4344 12232
rect 4203 12192 4344 12220
rect 4203 12189 4215 12192
rect 4157 12183 4215 12189
rect 3436 12152 3464 12183
rect 4338 12180 4344 12192
rect 4396 12180 4402 12232
rect 4801 12223 4859 12229
rect 4801 12189 4813 12223
rect 4847 12220 4859 12223
rect 4890 12220 4896 12232
rect 4847 12192 4896 12220
rect 4847 12189 4859 12192
rect 4801 12183 4859 12189
rect 4890 12180 4896 12192
rect 4948 12180 4954 12232
rect 4982 12180 4988 12232
rect 5040 12180 5046 12232
rect 5077 12223 5135 12229
rect 5077 12189 5089 12223
rect 5123 12220 5135 12223
rect 5123 12192 5212 12220
rect 5123 12189 5135 12192
rect 5077 12183 5135 12189
rect 4617 12155 4675 12161
rect 4617 12152 4629 12155
rect 3436 12124 4629 12152
rect 4617 12121 4629 12124
rect 4663 12121 4675 12155
rect 4617 12115 4675 12121
rect 3237 12087 3295 12093
rect 3237 12053 3249 12087
rect 3283 12084 3295 12087
rect 3878 12084 3884 12096
rect 3283 12056 3884 12084
rect 3283 12053 3295 12056
rect 3237 12047 3295 12053
rect 3878 12044 3884 12056
rect 3936 12044 3942 12096
rect 4065 12087 4123 12093
rect 4065 12053 4077 12087
rect 4111 12084 4123 12087
rect 5184 12084 5212 12192
rect 5534 12180 5540 12232
rect 5592 12180 5598 12232
rect 5804 12223 5862 12229
rect 5804 12189 5816 12223
rect 5850 12189 5862 12223
rect 5804 12183 5862 12189
rect 5718 12112 5724 12164
rect 5776 12152 5782 12164
rect 5828 12152 5856 12183
rect 6914 12180 6920 12232
rect 6972 12220 6978 12232
rect 7653 12223 7711 12229
rect 7653 12220 7665 12223
rect 6972 12192 7665 12220
rect 6972 12180 6978 12192
rect 7653 12189 7665 12192
rect 7699 12189 7711 12223
rect 7653 12183 7711 12189
rect 9766 12180 9772 12232
rect 9824 12180 9830 12232
rect 10873 12223 10931 12229
rect 10873 12189 10885 12223
rect 10919 12220 10931 12223
rect 11330 12220 11336 12232
rect 10919 12192 11336 12220
rect 10919 12189 10931 12192
rect 10873 12183 10931 12189
rect 11330 12180 11336 12192
rect 11388 12180 11394 12232
rect 11422 12180 11428 12232
rect 11480 12220 11486 12232
rect 11977 12223 12035 12229
rect 11977 12220 11989 12223
rect 11480 12192 11989 12220
rect 11480 12180 11486 12192
rect 11977 12189 11989 12192
rect 12023 12189 12035 12223
rect 12176 12220 12204 12260
rect 12253 12257 12265 12291
rect 12299 12288 12311 12291
rect 13280 12288 13308 12328
rect 14826 12316 14832 12328
rect 14884 12316 14890 12368
rect 17037 12359 17095 12365
rect 17037 12325 17049 12359
rect 17083 12356 17095 12359
rect 24688 12356 24716 12396
rect 17083 12328 24716 12356
rect 27448 12356 27476 12396
rect 27890 12384 27896 12436
rect 27948 12384 27954 12436
rect 28074 12384 28080 12436
rect 28132 12424 28138 12436
rect 28258 12424 28264 12436
rect 28132 12396 28264 12424
rect 28132 12384 28138 12396
rect 28258 12384 28264 12396
rect 28316 12384 28322 12436
rect 28629 12427 28687 12433
rect 28629 12393 28641 12427
rect 28675 12424 28687 12427
rect 28718 12424 28724 12436
rect 28675 12396 28724 12424
rect 28675 12393 28687 12396
rect 28629 12387 28687 12393
rect 28718 12384 28724 12396
rect 28776 12384 28782 12436
rect 30282 12384 30288 12436
rect 30340 12384 30346 12436
rect 33318 12384 33324 12436
rect 33376 12424 33382 12436
rect 33413 12427 33471 12433
rect 33413 12424 33425 12427
rect 33376 12396 33425 12424
rect 33376 12384 33382 12396
rect 33413 12393 33425 12396
rect 33459 12393 33471 12427
rect 33413 12387 33471 12393
rect 38654 12384 38660 12436
rect 38712 12424 38718 12436
rect 38933 12427 38991 12433
rect 38933 12424 38945 12427
rect 38712 12396 38945 12424
rect 38712 12384 38718 12396
rect 38933 12393 38945 12396
rect 38979 12393 38991 12427
rect 38933 12387 38991 12393
rect 40034 12384 40040 12436
rect 40092 12384 40098 12436
rect 28350 12356 28356 12368
rect 27448 12328 28356 12356
rect 17083 12325 17095 12328
rect 17037 12319 17095 12325
rect 28350 12316 28356 12328
rect 28408 12316 28414 12368
rect 28534 12316 28540 12368
rect 28592 12356 28598 12368
rect 28813 12359 28871 12365
rect 28813 12356 28825 12359
rect 28592 12328 28825 12356
rect 28592 12316 28598 12328
rect 28813 12325 28825 12328
rect 28859 12325 28871 12359
rect 28813 12319 28871 12325
rect 12299 12260 13308 12288
rect 13357 12291 13415 12297
rect 12299 12257 12311 12260
rect 12253 12251 12311 12257
rect 13357 12257 13369 12291
rect 13403 12288 13415 12291
rect 13446 12288 13452 12300
rect 13403 12260 13452 12288
rect 13403 12257 13415 12260
rect 13357 12251 13415 12257
rect 13446 12248 13452 12260
rect 13504 12248 13510 12300
rect 13725 12291 13783 12297
rect 13725 12257 13737 12291
rect 13771 12288 13783 12291
rect 13771 12260 16896 12288
rect 13771 12257 13783 12260
rect 13725 12251 13783 12257
rect 12618 12220 12624 12232
rect 12176 12192 12624 12220
rect 11977 12183 12035 12189
rect 5776 12124 5856 12152
rect 5776 12112 5782 12124
rect 5902 12112 5908 12164
rect 5960 12152 5966 12164
rect 11146 12152 11152 12164
rect 5960 12124 11152 12152
rect 5960 12112 5966 12124
rect 11146 12112 11152 12124
rect 11204 12112 11210 12164
rect 11241 12155 11299 12161
rect 11241 12121 11253 12155
rect 11287 12152 11299 12155
rect 11514 12152 11520 12164
rect 11287 12124 11520 12152
rect 11287 12121 11299 12124
rect 11241 12115 11299 12121
rect 4111 12056 5212 12084
rect 4111 12053 4123 12056
rect 4065 12047 4123 12053
rect 7742 12044 7748 12096
rect 7800 12044 7806 12096
rect 11054 12044 11060 12096
rect 11112 12084 11118 12096
rect 11256 12084 11284 12115
rect 11514 12112 11520 12124
rect 11572 12112 11578 12164
rect 11992 12152 12020 12183
rect 12618 12180 12624 12192
rect 12676 12180 12682 12232
rect 12710 12180 12716 12232
rect 12768 12220 12774 12232
rect 12805 12223 12863 12229
rect 12805 12220 12817 12223
rect 12768 12192 12817 12220
rect 12768 12180 12774 12192
rect 12805 12189 12817 12192
rect 12851 12189 12863 12223
rect 12805 12183 12863 12189
rect 13280 12192 13492 12220
rect 12250 12152 12256 12164
rect 11992 12124 12256 12152
rect 12250 12112 12256 12124
rect 12308 12112 12314 12164
rect 12345 12155 12403 12161
rect 12345 12121 12357 12155
rect 12391 12152 12403 12155
rect 13280 12152 13308 12192
rect 12391 12124 13308 12152
rect 12391 12121 12403 12124
rect 12345 12115 12403 12121
rect 11112 12056 11284 12084
rect 11112 12044 11118 12056
rect 11790 12044 11796 12096
rect 11848 12084 11854 12096
rect 13354 12084 13360 12096
rect 11848 12056 13360 12084
rect 11848 12044 11854 12056
rect 13354 12044 13360 12056
rect 13412 12044 13418 12096
rect 13464 12084 13492 12192
rect 13630 12180 13636 12232
rect 13688 12220 13694 12232
rect 16868 12229 16896 12260
rect 23842 12248 23848 12300
rect 23900 12248 23906 12300
rect 25317 12291 25375 12297
rect 25317 12288 25329 12291
rect 24780 12260 25329 12288
rect 14402 12223 14460 12229
rect 14402 12220 14414 12223
rect 13688 12192 14414 12220
rect 13688 12180 13694 12192
rect 14402 12189 14414 12192
rect 14448 12189 14460 12223
rect 14402 12183 14460 12189
rect 14921 12223 14979 12229
rect 14921 12189 14933 12223
rect 14967 12189 14979 12223
rect 14921 12183 14979 12189
rect 16853 12223 16911 12229
rect 16853 12189 16865 12223
rect 16899 12220 16911 12223
rect 16942 12220 16948 12232
rect 16899 12192 16948 12220
rect 16899 12189 16911 12192
rect 16853 12183 16911 12189
rect 14936 12152 14964 12183
rect 16942 12180 16948 12192
rect 17000 12180 17006 12232
rect 17129 12223 17187 12229
rect 17129 12189 17141 12223
rect 17175 12189 17187 12223
rect 17129 12183 17187 12189
rect 14384 12124 14964 12152
rect 17144 12152 17172 12183
rect 17770 12180 17776 12232
rect 17828 12220 17834 12232
rect 18049 12223 18107 12229
rect 18049 12220 18061 12223
rect 17828 12192 18061 12220
rect 17828 12180 17834 12192
rect 18049 12189 18061 12192
rect 18095 12189 18107 12223
rect 18049 12183 18107 12189
rect 20993 12223 21051 12229
rect 20993 12189 21005 12223
rect 21039 12220 21051 12223
rect 21358 12220 21364 12232
rect 21039 12192 21364 12220
rect 21039 12189 21051 12192
rect 20993 12183 21051 12189
rect 21358 12180 21364 12192
rect 21416 12180 21422 12232
rect 21450 12180 21456 12232
rect 21508 12180 21514 12232
rect 24780 12229 24808 12260
rect 25317 12257 25329 12260
rect 25363 12257 25375 12291
rect 25317 12251 25375 12257
rect 26142 12248 26148 12300
rect 26200 12248 26206 12300
rect 27430 12248 27436 12300
rect 27488 12288 27494 12300
rect 30558 12288 30564 12300
rect 27488 12260 28396 12288
rect 27488 12248 27494 12260
rect 21729 12223 21787 12229
rect 21729 12189 21741 12223
rect 21775 12220 21787 12223
rect 22373 12223 22431 12229
rect 22373 12220 22385 12223
rect 21775 12192 22385 12220
rect 21775 12189 21787 12192
rect 21729 12183 21787 12189
rect 22373 12189 22385 12192
rect 22419 12189 22431 12223
rect 22373 12183 22431 12189
rect 24765 12223 24823 12229
rect 24765 12189 24777 12223
rect 24811 12189 24823 12223
rect 24765 12183 24823 12189
rect 25222 12180 25228 12232
rect 25280 12180 25286 12232
rect 28368 12229 28396 12260
rect 29748 12260 30564 12288
rect 28353 12223 28411 12229
rect 28353 12189 28365 12223
rect 28399 12189 28411 12223
rect 28353 12183 28411 12189
rect 23661 12155 23719 12161
rect 17144 12124 23612 12152
rect 14384 12084 14412 12124
rect 13464 12056 14412 12084
rect 14458 12044 14464 12096
rect 14516 12044 14522 12096
rect 14936 12084 14964 12124
rect 19518 12084 19524 12096
rect 14936 12056 19524 12084
rect 19518 12044 19524 12056
rect 19576 12044 19582 12096
rect 20809 12087 20867 12093
rect 20809 12053 20821 12087
rect 20855 12084 20867 12087
rect 20990 12084 20996 12096
rect 20855 12056 20996 12084
rect 20855 12053 20867 12056
rect 20809 12047 20867 12053
rect 20990 12044 20996 12056
rect 21048 12044 21054 12096
rect 22094 12044 22100 12096
rect 22152 12084 22158 12096
rect 22189 12087 22247 12093
rect 22189 12084 22201 12087
rect 22152 12056 22201 12084
rect 22152 12044 22158 12056
rect 22189 12053 22201 12056
rect 22235 12053 22247 12087
rect 23584 12084 23612 12124
rect 23661 12121 23673 12155
rect 23707 12152 23719 12155
rect 23707 12124 26372 12152
rect 23707 12121 23719 12124
rect 23661 12115 23719 12121
rect 23753 12087 23811 12093
rect 23753 12084 23765 12087
rect 23584 12056 23765 12084
rect 22189 12047 22247 12053
rect 23753 12053 23765 12056
rect 23799 12084 23811 12087
rect 24946 12084 24952 12096
rect 23799 12056 24952 12084
rect 23799 12053 23811 12056
rect 23753 12047 23811 12053
rect 24946 12044 24952 12056
rect 25004 12044 25010 12096
rect 26344 12084 26372 12124
rect 26418 12112 26424 12164
rect 26476 12112 26482 12164
rect 26878 12112 26884 12164
rect 26936 12112 26942 12164
rect 28368 12152 28396 12183
rect 28534 12180 28540 12232
rect 28592 12180 28598 12232
rect 28626 12180 28632 12232
rect 28684 12180 28690 12232
rect 29748 12220 29776 12260
rect 30558 12248 30564 12260
rect 30616 12248 30622 12300
rect 31846 12288 31852 12300
rect 30760 12260 31852 12288
rect 28808 12192 29776 12220
rect 28808 12152 28836 12192
rect 30466 12180 30472 12232
rect 30524 12180 30530 12232
rect 30760 12229 30788 12260
rect 31846 12248 31852 12260
rect 31904 12248 31910 12300
rect 37185 12291 37243 12297
rect 37185 12288 37197 12291
rect 34900 12260 37197 12288
rect 34900 12232 34928 12260
rect 37185 12257 37197 12260
rect 37231 12288 37243 12291
rect 38194 12288 38200 12300
rect 37231 12260 38200 12288
rect 37231 12257 37243 12260
rect 37185 12251 37243 12257
rect 38194 12248 38200 12260
rect 38252 12248 38258 12300
rect 41506 12248 41512 12300
rect 41564 12248 41570 12300
rect 30745 12223 30803 12229
rect 30745 12220 30757 12223
rect 30576 12192 30757 12220
rect 28368 12124 28836 12152
rect 28902 12112 28908 12164
rect 28960 12152 28966 12164
rect 30576 12152 30604 12192
rect 30745 12189 30757 12192
rect 30791 12189 30803 12223
rect 30745 12183 30803 12189
rect 30926 12180 30932 12232
rect 30984 12220 30990 12232
rect 31205 12223 31263 12229
rect 31205 12220 31217 12223
rect 30984 12192 31217 12220
rect 30984 12180 30990 12192
rect 31205 12189 31217 12192
rect 31251 12189 31263 12223
rect 31205 12183 31263 12189
rect 33594 12180 33600 12232
rect 33652 12180 33658 12232
rect 34330 12180 34336 12232
rect 34388 12180 34394 12232
rect 34882 12180 34888 12232
rect 34940 12180 34946 12232
rect 40218 12180 40224 12232
rect 40276 12180 40282 12232
rect 41233 12223 41291 12229
rect 41233 12189 41245 12223
rect 41279 12220 41291 12223
rect 41414 12220 41420 12232
rect 41279 12192 41420 12220
rect 41279 12189 41291 12192
rect 41233 12183 41291 12189
rect 41414 12180 41420 12192
rect 41472 12180 41478 12232
rect 28960 12124 30604 12152
rect 30653 12155 30711 12161
rect 28960 12112 28966 12124
rect 30653 12121 30665 12155
rect 30699 12121 30711 12155
rect 30653 12115 30711 12121
rect 28626 12084 28632 12096
rect 26344 12056 28632 12084
rect 28626 12044 28632 12056
rect 28684 12084 28690 12096
rect 30668 12084 30696 12115
rect 31386 12112 31392 12164
rect 31444 12152 31450 12164
rect 31481 12155 31539 12161
rect 31481 12152 31493 12155
rect 31444 12124 31493 12152
rect 31444 12112 31450 12124
rect 31481 12121 31493 12124
rect 31527 12121 31539 12155
rect 33134 12152 33140 12164
rect 32706 12124 33140 12152
rect 31481 12115 31539 12121
rect 33134 12112 33140 12124
rect 33192 12112 33198 12164
rect 35161 12155 35219 12161
rect 35161 12121 35173 12155
rect 35207 12121 35219 12155
rect 36538 12152 36544 12164
rect 36386 12124 36544 12152
rect 35161 12115 35219 12121
rect 32490 12084 32496 12096
rect 28684 12056 32496 12084
rect 28684 12044 28690 12056
rect 32490 12044 32496 12056
rect 32548 12084 32554 12096
rect 32953 12087 33011 12093
rect 32953 12084 32965 12087
rect 32548 12056 32965 12084
rect 32548 12044 32554 12056
rect 32953 12053 32965 12056
rect 32999 12053 33011 12087
rect 32953 12047 33011 12053
rect 34149 12087 34207 12093
rect 34149 12053 34161 12087
rect 34195 12084 34207 12087
rect 35176 12084 35204 12115
rect 36538 12112 36544 12124
rect 36596 12112 36602 12164
rect 37458 12112 37464 12164
rect 37516 12112 37522 12164
rect 38102 12112 38108 12164
rect 38160 12112 38166 12164
rect 34195 12056 35204 12084
rect 34195 12053 34207 12056
rect 34149 12047 34207 12053
rect 36630 12044 36636 12096
rect 36688 12084 36694 12096
rect 39114 12084 39120 12096
rect 36688 12056 39120 12084
rect 36688 12044 36694 12056
rect 39114 12044 39120 12056
rect 39172 12044 39178 12096
rect 1104 11994 45051 12016
rect 1104 11942 11896 11994
rect 11948 11942 11960 11994
rect 12012 11942 12024 11994
rect 12076 11942 12088 11994
rect 12140 11942 12152 11994
rect 12204 11942 22843 11994
rect 22895 11942 22907 11994
rect 22959 11942 22971 11994
rect 23023 11942 23035 11994
rect 23087 11942 23099 11994
rect 23151 11942 33790 11994
rect 33842 11942 33854 11994
rect 33906 11942 33918 11994
rect 33970 11942 33982 11994
rect 34034 11942 34046 11994
rect 34098 11942 44737 11994
rect 44789 11942 44801 11994
rect 44853 11942 44865 11994
rect 44917 11942 44929 11994
rect 44981 11942 44993 11994
rect 45045 11942 45051 11994
rect 1104 11920 45051 11942
rect 4062 11840 4068 11892
rect 4120 11840 4126 11892
rect 4982 11840 4988 11892
rect 5040 11880 5046 11892
rect 5997 11883 6055 11889
rect 5997 11880 6009 11883
rect 5040 11852 6009 11880
rect 5040 11840 5046 11852
rect 5997 11849 6009 11852
rect 6043 11849 6055 11883
rect 5997 11843 6055 11849
rect 11149 11883 11207 11889
rect 11149 11849 11161 11883
rect 11195 11880 11207 11883
rect 11238 11880 11244 11892
rect 11195 11852 11244 11880
rect 11195 11849 11207 11852
rect 11149 11843 11207 11849
rect 11238 11840 11244 11852
rect 11296 11840 11302 11892
rect 12710 11840 12716 11892
rect 12768 11840 12774 11892
rect 14458 11840 14464 11892
rect 14516 11880 14522 11892
rect 16853 11883 16911 11889
rect 16853 11880 16865 11883
rect 14516 11852 16865 11880
rect 14516 11840 14522 11852
rect 16853 11849 16865 11852
rect 16899 11849 16911 11883
rect 16853 11843 16911 11849
rect 18046 11840 18052 11892
rect 18104 11840 18110 11892
rect 18693 11883 18751 11889
rect 18693 11849 18705 11883
rect 18739 11880 18751 11883
rect 19426 11880 19432 11892
rect 18739 11852 19432 11880
rect 18739 11849 18751 11852
rect 18693 11843 18751 11849
rect 19426 11840 19432 11852
rect 19484 11840 19490 11892
rect 19518 11840 19524 11892
rect 19576 11880 19582 11892
rect 20717 11883 20775 11889
rect 20717 11880 20729 11883
rect 19576 11852 20729 11880
rect 19576 11840 19582 11852
rect 20717 11849 20729 11852
rect 20763 11849 20775 11883
rect 20717 11843 20775 11849
rect 20898 11840 20904 11892
rect 20956 11880 20962 11892
rect 21082 11880 21088 11892
rect 20956 11852 21088 11880
rect 20956 11840 20962 11852
rect 21082 11840 21088 11852
rect 21140 11840 21146 11892
rect 21358 11840 21364 11892
rect 21416 11880 21422 11892
rect 22005 11883 22063 11889
rect 22005 11880 22017 11883
rect 21416 11852 22017 11880
rect 21416 11840 21422 11852
rect 22005 11849 22017 11852
rect 22051 11849 22063 11883
rect 22005 11843 22063 11849
rect 22462 11840 22468 11892
rect 22520 11840 22526 11892
rect 26418 11840 26424 11892
rect 26476 11840 26482 11892
rect 32677 11883 32735 11889
rect 26528 11852 30972 11880
rect 4080 11812 4108 11840
rect 5902 11812 5908 11824
rect 3804 11784 4108 11812
rect 5736 11784 5908 11812
rect 2130 11704 2136 11756
rect 2188 11704 2194 11756
rect 3326 11704 3332 11756
rect 3384 11744 3390 11756
rect 3804 11753 3832 11784
rect 3789 11747 3847 11753
rect 3789 11744 3801 11747
rect 3384 11716 3801 11744
rect 3384 11704 3390 11716
rect 3789 11713 3801 11716
rect 3835 11713 3847 11747
rect 3789 11707 3847 11713
rect 3878 11704 3884 11756
rect 3936 11744 3942 11756
rect 4045 11747 4103 11753
rect 4045 11744 4057 11747
rect 3936 11716 4057 11744
rect 3936 11704 3942 11716
rect 4045 11713 4057 11716
rect 4091 11713 4103 11747
rect 4045 11707 4103 11713
rect 4338 11704 4344 11756
rect 4396 11744 4402 11756
rect 5736 11753 5764 11784
rect 5902 11772 5908 11784
rect 5960 11772 5966 11824
rect 10781 11815 10839 11821
rect 10781 11781 10793 11815
rect 10827 11812 10839 11815
rect 10827 11784 12112 11812
rect 10827 11781 10839 11784
rect 10781 11775 10839 11781
rect 12084 11756 12112 11784
rect 16942 11772 16948 11824
rect 17000 11812 17006 11824
rect 23842 11812 23848 11824
rect 17000 11784 23848 11812
rect 17000 11772 17006 11784
rect 23842 11772 23848 11784
rect 23900 11772 23906 11824
rect 24946 11772 24952 11824
rect 25004 11812 25010 11824
rect 26528 11812 26556 11852
rect 27801 11815 27859 11821
rect 27801 11812 27813 11815
rect 25004 11784 26556 11812
rect 26712 11784 27813 11812
rect 25004 11772 25010 11784
rect 5721 11747 5779 11753
rect 4396 11716 5212 11744
rect 4396 11704 4402 11716
rect 2774 11636 2780 11688
rect 2832 11636 2838 11688
rect 5184 11617 5212 11716
rect 5721 11713 5733 11747
rect 5767 11713 5779 11747
rect 5721 11707 5779 11713
rect 5169 11611 5227 11617
rect 5169 11577 5181 11611
rect 5215 11608 5227 11611
rect 5736 11608 5764 11707
rect 5810 11704 5816 11756
rect 5868 11704 5874 11756
rect 6914 11704 6920 11756
rect 6972 11704 6978 11756
rect 7009 11747 7067 11753
rect 7009 11713 7021 11747
rect 7055 11744 7067 11747
rect 7650 11744 7656 11756
rect 7055 11716 7656 11744
rect 7055 11713 7067 11716
rect 7009 11707 7067 11713
rect 7650 11704 7656 11716
rect 7708 11704 7714 11756
rect 7742 11704 7748 11756
rect 7800 11744 7806 11756
rect 10597 11747 10655 11753
rect 10597 11744 10609 11747
rect 7800 11716 10609 11744
rect 7800 11704 7806 11716
rect 10597 11713 10609 11716
rect 10643 11713 10655 11747
rect 10597 11707 10655 11713
rect 7098 11636 7104 11688
rect 7156 11636 7162 11688
rect 10612 11676 10640 11707
rect 10870 11704 10876 11756
rect 10928 11704 10934 11756
rect 10965 11747 11023 11753
rect 10965 11713 10977 11747
rect 11011 11744 11023 11747
rect 11422 11744 11428 11756
rect 11011 11716 11428 11744
rect 11011 11713 11023 11716
rect 10965 11707 11023 11713
rect 11422 11704 11428 11716
rect 11480 11704 11486 11756
rect 11790 11704 11796 11756
rect 11848 11744 11854 11756
rect 11977 11747 12035 11753
rect 11848 11742 11928 11744
rect 11977 11742 11989 11747
rect 11848 11716 11989 11742
rect 11848 11704 11854 11716
rect 11900 11714 11989 11716
rect 11977 11713 11989 11714
rect 12023 11713 12035 11747
rect 11977 11707 12035 11713
rect 12066 11704 12072 11756
rect 12124 11744 12130 11756
rect 12161 11747 12219 11753
rect 12161 11744 12173 11747
rect 12124 11716 12173 11744
rect 12124 11704 12130 11716
rect 12161 11713 12173 11716
rect 12207 11713 12219 11747
rect 12161 11707 12219 11713
rect 12342 11704 12348 11756
rect 12400 11704 12406 11756
rect 12434 11704 12440 11756
rect 12492 11744 12498 11756
rect 12529 11747 12587 11753
rect 12529 11744 12541 11747
rect 12492 11716 12541 11744
rect 12492 11704 12498 11716
rect 12529 11713 12541 11716
rect 12575 11713 12587 11747
rect 12529 11707 12587 11713
rect 13541 11747 13599 11753
rect 13541 11713 13553 11747
rect 13587 11713 13599 11747
rect 13541 11707 13599 11713
rect 13633 11747 13691 11753
rect 13633 11713 13645 11747
rect 13679 11744 13691 11747
rect 17218 11744 17224 11756
rect 13679 11716 17224 11744
rect 13679 11713 13691 11716
rect 13633 11707 13691 11713
rect 12253 11679 12311 11685
rect 12253 11676 12265 11679
rect 10612 11648 12265 11676
rect 12253 11645 12265 11648
rect 12299 11645 12311 11679
rect 12253 11639 12311 11645
rect 5215 11580 5764 11608
rect 12360 11608 12388 11704
rect 13173 11611 13231 11617
rect 13173 11608 13185 11611
rect 12360 11580 13185 11608
rect 5215 11577 5227 11580
rect 5169 11571 5227 11577
rect 13173 11577 13185 11580
rect 13219 11577 13231 11611
rect 13173 11571 13231 11577
rect 6549 11543 6607 11549
rect 6549 11509 6561 11543
rect 6595 11540 6607 11543
rect 7926 11540 7932 11552
rect 6595 11512 7932 11540
rect 6595 11509 6607 11512
rect 6549 11503 6607 11509
rect 7926 11500 7932 11512
rect 7984 11500 7990 11552
rect 11238 11500 11244 11552
rect 11296 11540 11302 11552
rect 13556 11540 13584 11707
rect 17218 11704 17224 11716
rect 17276 11704 17282 11756
rect 17313 11747 17371 11753
rect 17313 11713 17325 11747
rect 17359 11744 17371 11747
rect 17359 11716 18184 11744
rect 17359 11713 17371 11716
rect 17313 11707 17371 11713
rect 13722 11636 13728 11688
rect 13780 11676 13786 11688
rect 17497 11679 17555 11685
rect 17497 11676 17509 11679
rect 13780 11648 17509 11676
rect 13780 11636 13786 11648
rect 17497 11645 17509 11648
rect 17543 11645 17555 11679
rect 18156 11676 18184 11716
rect 18230 11704 18236 11756
rect 18288 11704 18294 11756
rect 18874 11704 18880 11756
rect 18932 11704 18938 11756
rect 22002 11744 22008 11756
rect 21192 11716 22008 11744
rect 21192 11688 21220 11716
rect 22002 11704 22008 11716
rect 22060 11744 22066 11756
rect 22373 11747 22431 11753
rect 22373 11744 22385 11747
rect 22060 11716 22385 11744
rect 22060 11704 22066 11716
rect 22373 11713 22385 11716
rect 22419 11713 22431 11747
rect 22373 11707 22431 11713
rect 20898 11676 20904 11688
rect 18156 11648 20904 11676
rect 17497 11639 17555 11645
rect 17512 11608 17540 11639
rect 20898 11636 20904 11648
rect 20956 11636 20962 11688
rect 21174 11636 21180 11688
rect 21232 11636 21238 11688
rect 21361 11679 21419 11685
rect 21361 11645 21373 11679
rect 21407 11645 21419 11679
rect 21361 11639 21419 11645
rect 22649 11679 22707 11685
rect 22649 11645 22661 11679
rect 22695 11676 22707 11679
rect 22738 11676 22744 11688
rect 22695 11648 22744 11676
rect 22695 11645 22707 11648
rect 22649 11639 22707 11645
rect 21376 11608 21404 11639
rect 22738 11636 22744 11648
rect 22796 11636 22802 11688
rect 23860 11676 23888 11772
rect 26605 11747 26663 11753
rect 26605 11713 26617 11747
rect 26651 11742 26663 11747
rect 26712 11742 26740 11784
rect 27801 11781 27813 11784
rect 27847 11781 27859 11815
rect 27801 11775 27859 11781
rect 29181 11815 29239 11821
rect 29181 11781 29193 11815
rect 29227 11812 29239 11815
rect 30374 11812 30380 11824
rect 29227 11784 30380 11812
rect 29227 11781 29239 11784
rect 29181 11775 29239 11781
rect 30374 11772 30380 11784
rect 30432 11772 30438 11824
rect 30944 11821 30972 11852
rect 32677 11849 32689 11883
rect 32723 11880 32735 11883
rect 32766 11880 32772 11892
rect 32723 11852 32772 11880
rect 32723 11849 32735 11852
rect 32677 11843 32735 11849
rect 32766 11840 32772 11852
rect 32824 11840 32830 11892
rect 36541 11883 36599 11889
rect 36541 11849 36553 11883
rect 36587 11880 36599 11883
rect 37642 11880 37648 11892
rect 36587 11852 37648 11880
rect 36587 11849 36599 11852
rect 36541 11843 36599 11849
rect 37642 11840 37648 11852
rect 37700 11840 37706 11892
rect 30929 11815 30987 11821
rect 30929 11781 30941 11815
rect 30975 11781 30987 11815
rect 30929 11775 30987 11781
rect 35713 11815 35771 11821
rect 35713 11781 35725 11815
rect 35759 11812 35771 11815
rect 37090 11812 37096 11824
rect 35759 11784 37096 11812
rect 35759 11781 35771 11784
rect 35713 11775 35771 11781
rect 37090 11772 37096 11784
rect 37148 11772 37154 11824
rect 37182 11772 37188 11824
rect 37240 11812 37246 11824
rect 40954 11821 40960 11824
rect 40948 11812 40960 11821
rect 37240 11784 37504 11812
rect 37240 11772 37246 11784
rect 26651 11714 26740 11742
rect 26651 11713 26663 11714
rect 26605 11707 26663 11713
rect 27430 11704 27436 11756
rect 27488 11704 27494 11756
rect 27614 11704 27620 11756
rect 27672 11704 27678 11756
rect 28994 11704 29000 11756
rect 29052 11704 29058 11756
rect 30009 11747 30067 11753
rect 30009 11713 30021 11747
rect 30055 11713 30067 11747
rect 30009 11707 30067 11713
rect 28166 11676 28172 11688
rect 23860 11648 28172 11676
rect 28166 11636 28172 11648
rect 28224 11676 28230 11688
rect 28902 11676 28908 11688
rect 28224 11648 28908 11676
rect 28224 11636 28230 11648
rect 28902 11636 28908 11648
rect 28960 11676 28966 11688
rect 30024 11676 30052 11707
rect 30650 11704 30656 11756
rect 30708 11704 30714 11756
rect 30834 11704 30840 11756
rect 30892 11704 30898 11756
rect 31018 11704 31024 11756
rect 31076 11744 31082 11756
rect 31202 11744 31208 11756
rect 31076 11716 31208 11744
rect 31076 11704 31082 11716
rect 31202 11704 31208 11716
rect 31260 11704 31266 11756
rect 32306 11704 32312 11756
rect 32364 11704 32370 11756
rect 32490 11704 32496 11756
rect 32548 11704 32554 11756
rect 33594 11704 33600 11756
rect 33652 11744 33658 11756
rect 35621 11747 35679 11753
rect 35621 11744 35633 11747
rect 33652 11716 35633 11744
rect 33652 11704 33658 11716
rect 35621 11713 35633 11716
rect 35667 11713 35679 11747
rect 35621 11707 35679 11713
rect 35894 11704 35900 11756
rect 35952 11744 35958 11756
rect 36265 11747 36323 11753
rect 36265 11744 36277 11747
rect 35952 11716 36277 11744
rect 35952 11704 35958 11716
rect 36265 11713 36277 11716
rect 36311 11713 36323 11747
rect 36265 11707 36323 11713
rect 36354 11704 36360 11756
rect 36412 11704 36418 11756
rect 36633 11747 36691 11753
rect 36633 11713 36645 11747
rect 36679 11744 36691 11747
rect 37274 11744 37280 11756
rect 36679 11716 37280 11744
rect 36679 11713 36691 11716
rect 36633 11707 36691 11713
rect 37274 11704 37280 11716
rect 37332 11704 37338 11756
rect 37476 11753 37504 11784
rect 38396 11784 40724 11812
rect 40915 11784 40960 11812
rect 37461 11747 37519 11753
rect 37461 11713 37473 11747
rect 37507 11713 37519 11747
rect 37461 11707 37519 11713
rect 38194 11704 38200 11756
rect 38252 11744 38258 11756
rect 38396 11753 38424 11784
rect 40696 11756 40724 11784
rect 40948 11775 40960 11784
rect 40954 11772 40960 11775
rect 41012 11772 41018 11824
rect 38654 11753 38660 11756
rect 38381 11747 38439 11753
rect 38381 11744 38393 11747
rect 38252 11716 38393 11744
rect 38252 11704 38258 11716
rect 38381 11713 38393 11716
rect 38427 11713 38439 11747
rect 38381 11707 38439 11713
rect 38648 11707 38660 11753
rect 38654 11704 38660 11707
rect 38712 11704 38718 11756
rect 40678 11704 40684 11756
rect 40736 11704 40742 11756
rect 28960 11648 30052 11676
rect 30668 11676 30696 11704
rect 35986 11676 35992 11688
rect 30668 11648 35992 11676
rect 28960 11636 28966 11648
rect 35986 11636 35992 11648
rect 36044 11636 36050 11688
rect 36446 11636 36452 11688
rect 36504 11676 36510 11688
rect 37553 11679 37611 11685
rect 37553 11676 37565 11679
rect 36504 11648 37565 11676
rect 36504 11636 36510 11648
rect 37553 11645 37565 11648
rect 37599 11645 37611 11679
rect 37553 11639 37611 11645
rect 25590 11608 25596 11620
rect 17512 11580 25596 11608
rect 25590 11568 25596 11580
rect 25648 11568 25654 11620
rect 27614 11568 27620 11620
rect 27672 11608 27678 11620
rect 27672 11580 30144 11608
rect 27672 11568 27678 11580
rect 11296 11512 13584 11540
rect 11296 11500 11302 11512
rect 20070 11500 20076 11552
rect 20128 11540 20134 11552
rect 20806 11540 20812 11552
rect 20128 11512 20812 11540
rect 20128 11500 20134 11512
rect 20806 11500 20812 11512
rect 20864 11500 20870 11552
rect 20898 11500 20904 11552
rect 20956 11540 20962 11552
rect 21450 11540 21456 11552
rect 20956 11512 21456 11540
rect 20956 11500 20962 11512
rect 21450 11500 21456 11512
rect 21508 11540 21514 11552
rect 22278 11540 22284 11552
rect 21508 11512 22284 11540
rect 21508 11500 21514 11512
rect 22278 11500 22284 11512
rect 22336 11540 22342 11552
rect 23382 11540 23388 11552
rect 22336 11512 23388 11540
rect 22336 11500 22342 11512
rect 23382 11500 23388 11512
rect 23440 11540 23446 11552
rect 27154 11540 27160 11552
rect 23440 11512 27160 11540
rect 23440 11500 23446 11512
rect 27154 11500 27160 11512
rect 27212 11500 27218 11552
rect 30116 11549 30144 11580
rect 30466 11568 30472 11620
rect 30524 11608 30530 11620
rect 30524 11580 32536 11608
rect 30524 11568 30530 11580
rect 30101 11543 30159 11549
rect 30101 11509 30113 11543
rect 30147 11540 30159 11543
rect 31018 11540 31024 11552
rect 30147 11512 31024 11540
rect 30147 11509 30159 11512
rect 30101 11503 30159 11509
rect 31018 11500 31024 11512
rect 31076 11500 31082 11552
rect 31205 11543 31263 11549
rect 31205 11509 31217 11543
rect 31251 11540 31263 11543
rect 32214 11540 32220 11552
rect 31251 11512 32220 11540
rect 31251 11509 31263 11512
rect 31205 11503 31263 11509
rect 32214 11500 32220 11512
rect 32272 11500 32278 11552
rect 32508 11549 32536 11580
rect 32493 11543 32551 11549
rect 32493 11509 32505 11543
rect 32539 11540 32551 11543
rect 36630 11540 36636 11552
rect 32539 11512 36636 11540
rect 32539 11509 32551 11512
rect 32493 11503 32551 11509
rect 36630 11500 36636 11512
rect 36688 11500 36694 11552
rect 37458 11500 37464 11552
rect 37516 11540 37522 11552
rect 37918 11540 37924 11552
rect 37516 11512 37924 11540
rect 37516 11500 37522 11512
rect 37918 11500 37924 11512
rect 37976 11540 37982 11552
rect 39761 11543 39819 11549
rect 39761 11540 39773 11543
rect 37976 11512 39773 11540
rect 37976 11500 37982 11512
rect 39761 11509 39773 11512
rect 39807 11509 39819 11543
rect 39761 11503 39819 11509
rect 41874 11500 41880 11552
rect 41932 11540 41938 11552
rect 42061 11543 42119 11549
rect 42061 11540 42073 11543
rect 41932 11512 42073 11540
rect 41932 11500 41938 11512
rect 42061 11509 42073 11512
rect 42107 11509 42119 11543
rect 42061 11503 42119 11509
rect 1104 11450 44896 11472
rect 1104 11398 6423 11450
rect 6475 11398 6487 11450
rect 6539 11398 6551 11450
rect 6603 11398 6615 11450
rect 6667 11398 6679 11450
rect 6731 11398 17370 11450
rect 17422 11398 17434 11450
rect 17486 11398 17498 11450
rect 17550 11398 17562 11450
rect 17614 11398 17626 11450
rect 17678 11398 28317 11450
rect 28369 11398 28381 11450
rect 28433 11398 28445 11450
rect 28497 11398 28509 11450
rect 28561 11398 28573 11450
rect 28625 11398 39264 11450
rect 39316 11398 39328 11450
rect 39380 11398 39392 11450
rect 39444 11398 39456 11450
rect 39508 11398 39520 11450
rect 39572 11398 44896 11450
rect 1104 11376 44896 11398
rect 3418 11296 3424 11348
rect 3476 11296 3482 11348
rect 4430 11296 4436 11348
rect 4488 11336 4494 11348
rect 5350 11336 5356 11348
rect 4488 11308 5356 11336
rect 4488 11296 4494 11308
rect 5350 11296 5356 11308
rect 5408 11296 5414 11348
rect 6914 11296 6920 11348
rect 6972 11336 6978 11348
rect 7285 11339 7343 11345
rect 7285 11336 7297 11339
rect 6972 11308 7297 11336
rect 6972 11296 6978 11308
rect 7285 11305 7297 11308
rect 7331 11305 7343 11339
rect 7285 11299 7343 11305
rect 9858 11296 9864 11348
rect 9916 11336 9922 11348
rect 10781 11339 10839 11345
rect 10781 11336 10793 11339
rect 9916 11308 10793 11336
rect 9916 11296 9922 11308
rect 10781 11305 10793 11308
rect 10827 11305 10839 11339
rect 10781 11299 10839 11305
rect 11977 11339 12035 11345
rect 11977 11305 11989 11339
rect 12023 11336 12035 11339
rect 12066 11336 12072 11348
rect 12023 11308 12072 11336
rect 12023 11305 12035 11308
rect 11977 11299 12035 11305
rect 12066 11296 12072 11308
rect 12124 11296 12130 11348
rect 13446 11296 13452 11348
rect 13504 11296 13510 11348
rect 17681 11339 17739 11345
rect 17681 11305 17693 11339
rect 17727 11336 17739 11339
rect 17770 11336 17776 11348
rect 17727 11308 17776 11336
rect 17727 11305 17739 11308
rect 17681 11299 17739 11305
rect 17770 11296 17776 11308
rect 17828 11296 17834 11348
rect 20070 11296 20076 11348
rect 20128 11296 20134 11348
rect 23201 11339 23259 11345
rect 23201 11336 23213 11339
rect 20824 11308 23213 11336
rect 7745 11271 7803 11277
rect 7745 11237 7757 11271
rect 7791 11237 7803 11271
rect 13722 11268 13728 11280
rect 7745 11231 7803 11237
rect 12636 11240 13728 11268
rect 4614 11160 4620 11212
rect 4672 11160 4678 11212
rect 2041 11135 2099 11141
rect 2041 11101 2053 11135
rect 2087 11132 2099 11135
rect 3326 11132 3332 11144
rect 2087 11104 3332 11132
rect 2087 11101 2099 11104
rect 2041 11095 2099 11101
rect 3326 11092 3332 11104
rect 3384 11092 3390 11144
rect 3418 11092 3424 11144
rect 3476 11132 3482 11144
rect 4341 11135 4399 11141
rect 4341 11132 4353 11135
rect 3476 11104 4353 11132
rect 3476 11092 3482 11104
rect 4341 11101 4353 11104
rect 4387 11101 4399 11135
rect 4341 11095 4399 11101
rect 5166 11092 5172 11144
rect 5224 11092 5230 11144
rect 5534 11092 5540 11144
rect 5592 11132 5598 11144
rect 5905 11135 5963 11141
rect 5905 11132 5917 11135
rect 5592 11104 5917 11132
rect 5592 11092 5598 11104
rect 5905 11101 5917 11104
rect 5951 11101 5963 11135
rect 5905 11095 5963 11101
rect 6172 11135 6230 11141
rect 6172 11101 6184 11135
rect 6218 11132 6230 11135
rect 7760 11132 7788 11231
rect 11238 11160 11244 11212
rect 11296 11160 11302 11212
rect 11425 11203 11483 11209
rect 11425 11169 11437 11203
rect 11471 11200 11483 11203
rect 12434 11200 12440 11212
rect 11471 11172 12440 11200
rect 11471 11169 11483 11172
rect 11425 11163 11483 11169
rect 12434 11160 12440 11172
rect 12492 11200 12498 11212
rect 12636 11209 12664 11240
rect 13722 11228 13728 11240
rect 13780 11228 13786 11280
rect 16853 11271 16911 11277
rect 16853 11237 16865 11271
rect 16899 11268 16911 11271
rect 18230 11268 18236 11280
rect 16899 11240 18236 11268
rect 16899 11237 16911 11240
rect 16853 11231 16911 11237
rect 18230 11228 18236 11240
rect 18288 11228 18294 11280
rect 20254 11228 20260 11280
rect 20312 11268 20318 11280
rect 20824 11268 20852 11308
rect 23201 11305 23213 11308
rect 23247 11305 23259 11339
rect 23201 11299 23259 11305
rect 25590 11296 25596 11348
rect 25648 11336 25654 11348
rect 30374 11336 30380 11348
rect 25648 11308 27016 11336
rect 25648 11296 25654 11308
rect 20312 11240 20852 11268
rect 20312 11228 20318 11240
rect 22002 11228 22008 11280
rect 22060 11268 22066 11280
rect 22465 11271 22523 11277
rect 22465 11268 22477 11271
rect 22060 11240 22477 11268
rect 22060 11228 22066 11240
rect 22465 11237 22477 11240
rect 22511 11237 22523 11271
rect 22465 11231 22523 11237
rect 12621 11203 12679 11209
rect 12621 11200 12633 11203
rect 12492 11172 12633 11200
rect 12492 11160 12498 11172
rect 12621 11169 12633 11172
rect 12667 11169 12679 11203
rect 14458 11200 14464 11212
rect 12621 11163 12679 11169
rect 13464 11172 14464 11200
rect 6218 11104 7788 11132
rect 6218 11101 6230 11104
rect 6172 11095 6230 11101
rect 7926 11092 7932 11144
rect 7984 11092 7990 11144
rect 9950 11092 9956 11144
rect 10008 11092 10014 11144
rect 13464 11141 13492 11172
rect 14458 11160 14464 11172
rect 14516 11160 14522 11212
rect 17126 11200 17132 11212
rect 16500 11172 17132 11200
rect 13449 11135 13507 11141
rect 13449 11101 13461 11135
rect 13495 11101 13507 11135
rect 13449 11095 13507 11101
rect 13630 11092 13636 11144
rect 13688 11092 13694 11144
rect 15378 11092 15384 11144
rect 15436 11132 15442 11144
rect 16500 11141 16528 11172
rect 17126 11160 17132 11172
rect 17184 11200 17190 11212
rect 17313 11203 17371 11209
rect 17313 11200 17325 11203
rect 17184 11172 17325 11200
rect 17184 11160 17190 11172
rect 17313 11169 17325 11172
rect 17359 11200 17371 11203
rect 18322 11200 18328 11212
rect 17359 11172 18328 11200
rect 17359 11169 17371 11172
rect 17313 11163 17371 11169
rect 18322 11160 18328 11172
rect 18380 11160 18386 11212
rect 19978 11160 19984 11212
rect 20036 11200 20042 11212
rect 20622 11200 20628 11212
rect 20036 11172 20628 11200
rect 20036 11160 20042 11172
rect 20622 11160 20628 11172
rect 20680 11160 20686 11212
rect 20714 11160 20720 11212
rect 20772 11160 20778 11212
rect 20990 11160 20996 11212
rect 21048 11160 21054 11212
rect 24854 11160 24860 11212
rect 24912 11200 24918 11212
rect 25133 11203 25191 11209
rect 25133 11200 25145 11203
rect 24912 11172 25145 11200
rect 24912 11160 24918 11172
rect 25133 11169 25145 11172
rect 25179 11169 25191 11203
rect 25133 11163 25191 11169
rect 25409 11203 25467 11209
rect 25409 11169 25421 11203
rect 25455 11200 25467 11203
rect 26786 11200 26792 11212
rect 25455 11172 26792 11200
rect 25455 11169 25467 11172
rect 25409 11163 25467 11169
rect 26786 11160 26792 11172
rect 26844 11160 26850 11212
rect 26878 11160 26884 11212
rect 26936 11160 26942 11212
rect 26988 11200 27016 11308
rect 28644 11308 30380 11336
rect 27154 11228 27160 11280
rect 27212 11268 27218 11280
rect 27890 11268 27896 11280
rect 27212 11240 27896 11268
rect 27212 11228 27218 11240
rect 27890 11228 27896 11240
rect 27948 11228 27954 11280
rect 27341 11203 27399 11209
rect 27341 11200 27353 11203
rect 26988 11172 27353 11200
rect 27341 11169 27353 11172
rect 27387 11200 27399 11203
rect 28534 11200 28540 11212
rect 27387 11172 28540 11200
rect 27387 11169 27399 11172
rect 27341 11163 27399 11169
rect 28534 11160 28540 11172
rect 28592 11160 28598 11212
rect 16485 11135 16543 11141
rect 16485 11132 16497 11135
rect 15436 11104 16497 11132
rect 15436 11092 15442 11104
rect 16485 11101 16497 11104
rect 16531 11101 16543 11135
rect 16485 11095 16543 11101
rect 16669 11135 16727 11141
rect 16669 11101 16681 11135
rect 16715 11101 16727 11135
rect 16669 11095 16727 11101
rect 17497 11135 17555 11141
rect 17497 11101 17509 11135
rect 17543 11132 17555 11135
rect 18230 11132 18236 11144
rect 17543 11104 18236 11132
rect 17543 11101 17555 11104
rect 17497 11095 17555 11101
rect 2308 11067 2366 11073
rect 2308 11033 2320 11067
rect 2354 11064 2366 11067
rect 2866 11064 2872 11076
rect 2354 11036 2872 11064
rect 2354 11033 2366 11036
rect 2308 11027 2366 11033
rect 2866 11024 2872 11036
rect 2924 11024 2930 11076
rect 3878 11024 3884 11076
rect 3936 11064 3942 11076
rect 4433 11067 4491 11073
rect 4433 11064 4445 11067
rect 3936 11036 4445 11064
rect 3936 11024 3942 11036
rect 4433 11033 4445 11036
rect 4479 11033 4491 11067
rect 4433 11027 4491 11033
rect 12345 11067 12403 11073
rect 12345 11033 12357 11067
rect 12391 11064 12403 11067
rect 13170 11064 13176 11076
rect 12391 11036 13176 11064
rect 12391 11033 12403 11036
rect 12345 11027 12403 11033
rect 13170 11024 13176 11036
rect 13228 11024 13234 11076
rect 16298 11024 16304 11076
rect 16356 11064 16362 11076
rect 16684 11064 16712 11095
rect 18230 11092 18236 11104
rect 18288 11092 18294 11144
rect 20257 11135 20315 11141
rect 20257 11101 20269 11135
rect 20303 11101 20315 11135
rect 20257 11095 20315 11101
rect 16356 11036 16712 11064
rect 20272 11064 20300 11095
rect 22094 11092 22100 11144
rect 22152 11092 22158 11144
rect 23382 11092 23388 11144
rect 23440 11092 23446 11144
rect 27525 11135 27583 11141
rect 27525 11101 27537 11135
rect 27571 11132 27583 11135
rect 27614 11132 27620 11144
rect 27571 11104 27620 11132
rect 27571 11101 27583 11104
rect 27525 11095 27583 11101
rect 27614 11092 27620 11104
rect 27672 11092 27678 11144
rect 28644 11141 28672 11308
rect 30374 11296 30380 11308
rect 30432 11296 30438 11348
rect 30558 11296 30564 11348
rect 30616 11336 30622 11348
rect 31570 11336 31576 11348
rect 30616 11308 31576 11336
rect 30616 11296 30622 11308
rect 31570 11296 31576 11308
rect 31628 11336 31634 11348
rect 32677 11339 32735 11345
rect 32677 11336 32689 11339
rect 31628 11308 32689 11336
rect 31628 11296 31634 11308
rect 32677 11305 32689 11308
rect 32723 11305 32735 11339
rect 32677 11299 32735 11305
rect 38654 11296 38660 11348
rect 38712 11336 38718 11348
rect 38841 11339 38899 11345
rect 38841 11336 38853 11339
rect 38712 11308 38853 11336
rect 38712 11296 38718 11308
rect 38841 11305 38853 11308
rect 38887 11305 38899 11339
rect 38841 11299 38899 11305
rect 40405 11339 40463 11345
rect 40405 11305 40417 11339
rect 40451 11336 40463 11339
rect 41046 11336 41052 11348
rect 40451 11308 41052 11336
rect 40451 11305 40463 11308
rect 40405 11299 40463 11305
rect 41046 11296 41052 11308
rect 41104 11296 41110 11348
rect 41414 11296 41420 11348
rect 41472 11296 41478 11348
rect 28718 11228 28724 11280
rect 28776 11268 28782 11280
rect 30285 11271 30343 11277
rect 28776 11240 29132 11268
rect 28776 11228 28782 11240
rect 29104 11209 29132 11240
rect 30285 11237 30297 11271
rect 30331 11237 30343 11271
rect 30285 11231 30343 11237
rect 29089 11203 29147 11209
rect 29089 11169 29101 11203
rect 29135 11169 29147 11203
rect 30300 11200 30328 11231
rect 35802 11228 35808 11280
rect 35860 11268 35866 11280
rect 37550 11268 37556 11280
rect 35860 11240 37556 11268
rect 35860 11228 35866 11240
rect 37550 11228 37556 11240
rect 37608 11228 37614 11280
rect 37737 11271 37795 11277
rect 37737 11237 37749 11271
rect 37783 11237 37795 11271
rect 37737 11231 37795 11237
rect 38289 11271 38347 11277
rect 38289 11237 38301 11271
rect 38335 11268 38347 11271
rect 40218 11268 40224 11280
rect 38335 11240 40224 11268
rect 38335 11237 38347 11240
rect 38289 11231 38347 11237
rect 31205 11203 31263 11209
rect 31205 11200 31217 11203
rect 30300 11172 31217 11200
rect 29089 11163 29147 11169
rect 31205 11169 31217 11172
rect 31251 11169 31263 11203
rect 31205 11163 31263 11169
rect 32214 11160 32220 11212
rect 32272 11200 32278 11212
rect 36078 11200 36084 11212
rect 32272 11172 33364 11200
rect 32272 11160 32278 11172
rect 28629 11135 28687 11141
rect 28629 11101 28641 11135
rect 28675 11101 28687 11135
rect 28813 11135 28871 11141
rect 28813 11132 28825 11135
rect 28629 11095 28687 11101
rect 28808 11101 28825 11132
rect 28859 11101 28871 11135
rect 28808 11095 28871 11101
rect 20714 11064 20720 11076
rect 20272 11036 20720 11064
rect 16356 11024 16362 11036
rect 20714 11024 20720 11036
rect 20772 11024 20778 11076
rect 26418 11024 26424 11076
rect 26476 11024 26482 11076
rect 27430 11024 27436 11076
rect 27488 11064 27494 11076
rect 27709 11067 27767 11073
rect 27709 11064 27721 11067
rect 27488 11036 27721 11064
rect 27488 11024 27494 11036
rect 27709 11033 27721 11036
rect 27755 11033 27767 11067
rect 27709 11027 27767 11033
rect 28721 11067 28779 11073
rect 28721 11033 28733 11067
rect 28767 11033 28779 11067
rect 28808 11064 28836 11095
rect 28902 11092 28908 11144
rect 28960 11141 28966 11144
rect 28960 11135 28989 11141
rect 28977 11101 28989 11135
rect 28960 11095 28989 11101
rect 28960 11092 28966 11095
rect 30466 11092 30472 11144
rect 30524 11092 30530 11144
rect 30926 11092 30932 11144
rect 30984 11092 30990 11144
rect 32306 11092 32312 11144
rect 32364 11092 32370 11144
rect 33336 11141 33364 11172
rect 35084 11172 36084 11200
rect 35084 11144 35112 11172
rect 36078 11160 36084 11172
rect 36136 11200 36142 11212
rect 37752 11200 37780 11231
rect 40218 11228 40224 11240
rect 40276 11228 40282 11280
rect 36136 11172 37688 11200
rect 37752 11172 39068 11200
rect 36136 11160 36142 11172
rect 33321 11135 33379 11141
rect 33321 11101 33333 11135
rect 33367 11101 33379 11135
rect 33321 11095 33379 11101
rect 33594 11092 33600 11144
rect 33652 11132 33658 11144
rect 33965 11135 34023 11141
rect 33965 11132 33977 11135
rect 33652 11104 33977 11132
rect 33652 11092 33658 11104
rect 33965 11101 33977 11104
rect 34011 11101 34023 11135
rect 33965 11095 34023 11101
rect 35066 11092 35072 11144
rect 35124 11092 35130 11144
rect 35986 11092 35992 11144
rect 36044 11092 36050 11144
rect 36170 11092 36176 11144
rect 36228 11132 36234 11144
rect 37182 11132 37188 11144
rect 36228 11104 37188 11132
rect 36228 11092 36234 11104
rect 37182 11092 37188 11104
rect 37240 11092 37246 11144
rect 37274 11092 37280 11144
rect 37332 11132 37338 11144
rect 37553 11135 37611 11141
rect 37553 11132 37565 11135
rect 37332 11104 37565 11132
rect 37332 11092 37338 11104
rect 37553 11101 37565 11104
rect 37599 11101 37611 11135
rect 37660 11132 37688 11172
rect 39040 11141 39068 11172
rect 41874 11160 41880 11212
rect 41932 11160 41938 11212
rect 41966 11160 41972 11212
rect 42024 11160 42030 11212
rect 38197 11135 38255 11141
rect 38197 11132 38209 11135
rect 37660 11104 38209 11132
rect 37553 11095 37611 11101
rect 38197 11101 38209 11104
rect 38243 11101 38255 11135
rect 38197 11095 38255 11101
rect 39025 11135 39083 11141
rect 39025 11101 39037 11135
rect 39071 11101 39083 11135
rect 39025 11095 39083 11101
rect 39114 11092 39120 11144
rect 39172 11132 39178 11144
rect 40221 11135 40279 11141
rect 40221 11132 40233 11135
rect 39172 11104 40233 11132
rect 39172 11092 39178 11104
rect 40221 11101 40233 11104
rect 40267 11101 40279 11135
rect 40221 11095 40279 11101
rect 44361 11135 44419 11141
rect 44361 11101 44373 11135
rect 44407 11132 44419 11135
rect 45002 11132 45008 11144
rect 44407 11104 45008 11132
rect 44407 11101 44419 11104
rect 44361 11095 44419 11101
rect 45002 11092 45008 11104
rect 45060 11092 45066 11144
rect 30650 11064 30656 11076
rect 28808 11036 30656 11064
rect 28721 11027 28779 11033
rect 3970 10956 3976 11008
rect 4028 10956 4034 11008
rect 9769 10999 9827 11005
rect 9769 10965 9781 10999
rect 9815 10996 9827 10999
rect 10686 10996 10692 11008
rect 9815 10968 10692 10996
rect 9815 10965 9827 10968
rect 9769 10959 9827 10965
rect 10686 10956 10692 10968
rect 10744 10956 10750 11008
rect 11146 10956 11152 11008
rect 11204 10956 11210 11008
rect 12250 10956 12256 11008
rect 12308 10996 12314 11008
rect 12437 10999 12495 11005
rect 12437 10996 12449 10999
rect 12308 10968 12449 10996
rect 12308 10956 12314 10968
rect 12437 10965 12449 10968
rect 12483 10965 12495 10999
rect 12437 10959 12495 10965
rect 16022 10956 16028 11008
rect 16080 10996 16086 11008
rect 20898 10996 20904 11008
rect 16080 10968 20904 10996
rect 16080 10956 16086 10968
rect 20898 10956 20904 10968
rect 20956 10956 20962 11008
rect 20990 10956 20996 11008
rect 21048 10996 21054 11008
rect 26694 10996 26700 11008
rect 21048 10968 26700 10996
rect 21048 10956 21054 10968
rect 26694 10956 26700 10968
rect 26752 10956 26758 11008
rect 27614 10956 27620 11008
rect 27672 10996 27678 11008
rect 28445 10999 28503 11005
rect 28445 10996 28457 10999
rect 27672 10968 28457 10996
rect 27672 10956 27678 10968
rect 28445 10965 28457 10968
rect 28491 10965 28503 10999
rect 28736 10996 28764 11027
rect 30650 11024 30656 11036
rect 30708 11024 30714 11076
rect 34790 11024 34796 11076
rect 34848 11064 34854 11076
rect 35802 11064 35808 11076
rect 34848 11036 35808 11064
rect 34848 11024 34854 11036
rect 35802 11024 35808 11036
rect 35860 11024 35866 11076
rect 37366 11024 37372 11076
rect 37424 11024 37430 11076
rect 37458 11024 37464 11076
rect 37516 11024 37522 11076
rect 39758 11024 39764 11076
rect 39816 11064 39822 11076
rect 40037 11067 40095 11073
rect 40037 11064 40049 11067
rect 39816 11036 40049 11064
rect 39816 11024 39822 11036
rect 40037 11033 40049 11036
rect 40083 11033 40095 11067
rect 40037 11027 40095 11033
rect 41782 11024 41788 11076
rect 41840 11024 41846 11076
rect 30282 10996 30288 11008
rect 28736 10968 30288 10996
rect 28445 10959 28503 10965
rect 30282 10956 30288 10968
rect 30340 10956 30346 11008
rect 33134 10956 33140 11008
rect 33192 10956 33198 11008
rect 33502 10956 33508 11008
rect 33560 10996 33566 11008
rect 33781 10999 33839 11005
rect 33781 10996 33793 10999
rect 33560 10968 33793 10996
rect 33560 10956 33566 10968
rect 33781 10965 33793 10968
rect 33827 10965 33839 10999
rect 33781 10959 33839 10965
rect 34514 10956 34520 11008
rect 34572 10996 34578 11008
rect 35253 10999 35311 11005
rect 35253 10996 35265 10999
rect 34572 10968 35265 10996
rect 34572 10956 34578 10968
rect 35253 10965 35265 10968
rect 35299 10965 35311 10999
rect 35253 10959 35311 10965
rect 36173 10999 36231 11005
rect 36173 10965 36185 10999
rect 36219 10996 36231 10999
rect 36814 10996 36820 11008
rect 36219 10968 36820 10996
rect 36219 10965 36231 10968
rect 36173 10959 36231 10965
rect 36814 10956 36820 10968
rect 36872 10996 36878 11008
rect 38102 10996 38108 11008
rect 36872 10968 38108 10996
rect 36872 10956 36878 10968
rect 38102 10956 38108 10968
rect 38160 10956 38166 11008
rect 1104 10906 45051 10928
rect 1104 10854 11896 10906
rect 11948 10854 11960 10906
rect 12012 10854 12024 10906
rect 12076 10854 12088 10906
rect 12140 10854 12152 10906
rect 12204 10854 22843 10906
rect 22895 10854 22907 10906
rect 22959 10854 22971 10906
rect 23023 10854 23035 10906
rect 23087 10854 23099 10906
rect 23151 10854 33790 10906
rect 33842 10854 33854 10906
rect 33906 10854 33918 10906
rect 33970 10854 33982 10906
rect 34034 10854 34046 10906
rect 34098 10854 44737 10906
rect 44789 10854 44801 10906
rect 44853 10854 44865 10906
rect 44917 10854 44929 10906
rect 44981 10854 44993 10906
rect 45045 10854 45051 10906
rect 1104 10832 45051 10854
rect 2685 10795 2743 10801
rect 2685 10761 2697 10795
rect 2731 10761 2743 10795
rect 2685 10755 2743 10761
rect 5721 10795 5779 10801
rect 5721 10761 5733 10795
rect 5767 10792 5779 10795
rect 7006 10792 7012 10804
rect 5767 10764 7012 10792
rect 5767 10761 5779 10764
rect 5721 10755 5779 10761
rect 2700 10724 2728 10755
rect 7006 10752 7012 10764
rect 7064 10752 7070 10804
rect 9950 10752 9956 10804
rect 10008 10792 10014 10804
rect 10413 10795 10471 10801
rect 10413 10792 10425 10795
rect 10008 10764 10425 10792
rect 10008 10752 10014 10764
rect 10413 10761 10425 10764
rect 10459 10761 10471 10795
rect 10413 10755 10471 10761
rect 10781 10795 10839 10801
rect 10781 10761 10793 10795
rect 10827 10792 10839 10795
rect 11238 10792 11244 10804
rect 10827 10764 11244 10792
rect 10827 10761 10839 10764
rect 10781 10755 10839 10761
rect 11238 10752 11244 10764
rect 11296 10752 11302 10804
rect 11330 10752 11336 10804
rect 11388 10792 11394 10804
rect 11793 10795 11851 10801
rect 11793 10792 11805 10795
rect 11388 10764 11805 10792
rect 11388 10752 11394 10764
rect 11793 10761 11805 10764
rect 11839 10761 11851 10795
rect 11793 10755 11851 10761
rect 12161 10795 12219 10801
rect 12161 10761 12173 10795
rect 12207 10792 12219 10795
rect 12250 10792 12256 10804
rect 12207 10764 12256 10792
rect 12207 10761 12219 10764
rect 12161 10755 12219 10761
rect 12250 10752 12256 10764
rect 12308 10752 12314 10804
rect 13814 10752 13820 10804
rect 13872 10792 13878 10804
rect 14277 10795 14335 10801
rect 14277 10792 14289 10795
rect 13872 10764 14289 10792
rect 13872 10752 13878 10764
rect 14277 10761 14289 10764
rect 14323 10761 14335 10795
rect 14277 10755 14335 10761
rect 15381 10795 15439 10801
rect 15381 10761 15393 10795
rect 15427 10792 15439 10795
rect 15427 10764 16988 10792
rect 15427 10761 15439 10764
rect 15381 10755 15439 10761
rect 3574 10727 3632 10733
rect 3574 10724 3586 10727
rect 2700 10696 3586 10724
rect 3574 10693 3586 10696
rect 3620 10693 3632 10727
rect 3574 10687 3632 10693
rect 5166 10684 5172 10736
rect 5224 10724 5230 10736
rect 7837 10727 7895 10733
rect 5224 10696 6914 10724
rect 5224 10684 5230 10696
rect 2869 10659 2927 10665
rect 2869 10625 2881 10659
rect 2915 10656 2927 10659
rect 3234 10656 3240 10668
rect 2915 10628 3240 10656
rect 2915 10625 2927 10628
rect 2869 10619 2927 10625
rect 3234 10616 3240 10628
rect 3292 10616 3298 10668
rect 3326 10616 3332 10668
rect 3384 10616 3390 10668
rect 4982 10616 4988 10668
rect 5040 10656 5046 10668
rect 5350 10656 5356 10668
rect 5040 10628 5356 10656
rect 5040 10616 5046 10628
rect 5350 10616 5356 10628
rect 5408 10616 5414 10668
rect 5537 10659 5595 10665
rect 5537 10625 5549 10659
rect 5583 10625 5595 10659
rect 5537 10619 5595 10625
rect 4338 10480 4344 10532
rect 4396 10520 4402 10532
rect 4709 10523 4767 10529
rect 4709 10520 4721 10523
rect 4396 10492 4721 10520
rect 4396 10480 4402 10492
rect 4709 10489 4721 10492
rect 4755 10520 4767 10523
rect 5552 10520 5580 10619
rect 4755 10492 5580 10520
rect 6886 10520 6914 10696
rect 7837 10693 7849 10727
rect 7883 10724 7895 10727
rect 14292 10724 14320 10755
rect 16960 10724 16988 10764
rect 17218 10752 17224 10804
rect 17276 10792 17282 10804
rect 18601 10795 18659 10801
rect 18601 10792 18613 10795
rect 17276 10764 18613 10792
rect 17276 10752 17282 10764
rect 18601 10761 18613 10764
rect 18647 10761 18659 10795
rect 18601 10755 18659 10761
rect 19242 10752 19248 10804
rect 19300 10792 19306 10804
rect 20990 10792 20996 10804
rect 19300 10764 20996 10792
rect 19300 10752 19306 10764
rect 20990 10752 20996 10764
rect 21048 10752 21054 10804
rect 21085 10795 21143 10801
rect 21085 10761 21097 10795
rect 21131 10792 21143 10795
rect 21174 10792 21180 10804
rect 21131 10764 21180 10792
rect 21131 10761 21143 10764
rect 21085 10755 21143 10761
rect 21174 10752 21180 10764
rect 21232 10752 21238 10804
rect 25590 10752 25596 10804
rect 25648 10752 25654 10804
rect 26694 10752 26700 10804
rect 26752 10792 26758 10804
rect 26752 10764 28764 10792
rect 26752 10752 26758 10764
rect 23198 10724 23204 10736
rect 7883 10696 13032 10724
rect 14292 10696 16896 10724
rect 16960 10696 17618 10724
rect 22066 10696 23204 10724
rect 7883 10693 7895 10696
rect 7837 10687 7895 10693
rect 11146 10616 11152 10668
rect 11204 10656 11210 10668
rect 12253 10659 12311 10665
rect 12253 10656 12265 10659
rect 11204 10628 12265 10656
rect 11204 10616 11210 10628
rect 12253 10625 12265 10628
rect 12299 10656 12311 10659
rect 12894 10656 12900 10668
rect 12299 10628 12900 10656
rect 12299 10625 12311 10628
rect 12253 10619 12311 10625
rect 12894 10616 12900 10628
rect 12952 10616 12958 10668
rect 13004 10665 13032 10696
rect 12989 10659 13047 10665
rect 12989 10625 13001 10659
rect 13035 10656 13047 10659
rect 13262 10656 13268 10668
rect 13035 10628 13268 10656
rect 13035 10625 13047 10628
rect 12989 10619 13047 10625
rect 13262 10616 13268 10628
rect 13320 10616 13326 10668
rect 15565 10660 15623 10665
rect 15565 10659 15700 10660
rect 15565 10625 15577 10659
rect 15611 10632 15700 10659
rect 15611 10625 15623 10632
rect 15565 10619 15623 10625
rect 10870 10548 10876 10600
rect 10928 10548 10934 10600
rect 10962 10548 10968 10600
rect 11020 10548 11026 10600
rect 12434 10548 12440 10600
rect 12492 10548 12498 10600
rect 15672 10588 15700 10632
rect 16022 10616 16028 10668
rect 16080 10616 16086 10668
rect 16868 10665 16896 10696
rect 16853 10659 16911 10665
rect 16853 10625 16865 10659
rect 16899 10625 16911 10659
rect 16853 10619 16911 10625
rect 20254 10616 20260 10668
rect 20312 10616 20318 10668
rect 21177 10659 21235 10665
rect 21177 10625 21189 10659
rect 21223 10656 21235 10659
rect 22066 10656 22094 10696
rect 23198 10684 23204 10696
rect 23256 10684 23262 10736
rect 25501 10727 25559 10733
rect 25501 10724 25513 10727
rect 23584 10696 25513 10724
rect 22554 10665 22560 10668
rect 21223 10628 22094 10656
rect 21223 10625 21235 10628
rect 21177 10619 21235 10625
rect 22548 10619 22560 10665
rect 22612 10656 22618 10668
rect 22612 10628 22648 10656
rect 22554 10616 22560 10619
rect 22612 10616 22618 10628
rect 15672 10560 16068 10588
rect 16040 10529 16068 10560
rect 16482 10548 16488 10600
rect 16540 10588 16546 10600
rect 17129 10591 17187 10597
rect 17129 10588 17141 10591
rect 16540 10560 17141 10588
rect 16540 10548 16546 10560
rect 17129 10557 17141 10560
rect 17175 10557 17187 10591
rect 17129 10551 17187 10557
rect 21361 10591 21419 10597
rect 21361 10557 21373 10591
rect 21407 10588 21419 10591
rect 21407 10560 22094 10588
rect 21407 10557 21419 10560
rect 21361 10551 21419 10557
rect 16025 10523 16083 10529
rect 6886 10492 15976 10520
rect 4755 10489 4767 10492
rect 4709 10483 4767 10489
rect 934 10412 940 10464
rect 992 10452 998 10464
rect 2774 10452 2780 10464
rect 992 10424 2780 10452
rect 992 10412 998 10424
rect 2774 10412 2780 10424
rect 2832 10412 2838 10464
rect 5534 10412 5540 10464
rect 5592 10452 5598 10464
rect 9125 10455 9183 10461
rect 9125 10452 9137 10455
rect 5592 10424 9137 10452
rect 5592 10412 5598 10424
rect 9125 10421 9137 10424
rect 9171 10452 9183 10455
rect 10134 10452 10140 10464
rect 9171 10424 10140 10452
rect 9171 10421 9183 10424
rect 9125 10415 9183 10421
rect 10134 10412 10140 10424
rect 10192 10452 10198 10464
rect 10318 10452 10324 10464
rect 10192 10424 10324 10452
rect 10192 10412 10198 10424
rect 10318 10412 10324 10424
rect 10376 10412 10382 10464
rect 10870 10412 10876 10464
rect 10928 10452 10934 10464
rect 15194 10452 15200 10464
rect 10928 10424 15200 10452
rect 10928 10412 10934 10424
rect 15194 10412 15200 10424
rect 15252 10452 15258 10464
rect 15654 10452 15660 10464
rect 15252 10424 15660 10452
rect 15252 10412 15258 10424
rect 15654 10412 15660 10424
rect 15712 10412 15718 10464
rect 15948 10452 15976 10492
rect 16025 10489 16037 10523
rect 16071 10489 16083 10523
rect 19702 10520 19708 10532
rect 16025 10483 16083 10489
rect 18524 10492 19708 10520
rect 18524 10452 18552 10492
rect 19702 10480 19708 10492
rect 19760 10480 19766 10532
rect 20073 10523 20131 10529
rect 20073 10489 20085 10523
rect 20119 10520 20131 10523
rect 21266 10520 21272 10532
rect 20119 10492 21272 10520
rect 20119 10489 20131 10492
rect 20073 10483 20131 10489
rect 21266 10480 21272 10492
rect 21324 10480 21330 10532
rect 15948 10424 18552 10452
rect 18598 10412 18604 10464
rect 18656 10452 18662 10464
rect 20717 10455 20775 10461
rect 20717 10452 20729 10455
rect 18656 10424 20729 10452
rect 18656 10412 18662 10424
rect 20717 10421 20729 10424
rect 20763 10421 20775 10455
rect 22066 10452 22094 10560
rect 22186 10548 22192 10600
rect 22244 10588 22250 10600
rect 22281 10591 22339 10597
rect 22281 10588 22293 10591
rect 22244 10560 22293 10588
rect 22244 10548 22250 10560
rect 22281 10557 22293 10560
rect 22327 10557 22339 10591
rect 22281 10551 22339 10557
rect 23584 10452 23612 10696
rect 25501 10693 25513 10696
rect 25547 10724 25559 10727
rect 26878 10724 26884 10736
rect 25547 10696 26884 10724
rect 25547 10693 25559 10696
rect 25501 10687 25559 10693
rect 26878 10684 26884 10696
rect 26936 10684 26942 10736
rect 28166 10684 28172 10736
rect 28224 10684 28230 10736
rect 28736 10724 28764 10764
rect 30926 10752 30932 10804
rect 30984 10752 30990 10804
rect 31726 10764 34744 10792
rect 31478 10724 31484 10736
rect 28736 10696 31484 10724
rect 31478 10684 31484 10696
rect 31536 10684 31542 10736
rect 25222 10616 25228 10668
rect 25280 10656 25286 10668
rect 26050 10656 26056 10668
rect 25280 10628 26056 10656
rect 25280 10616 25286 10628
rect 26050 10616 26056 10628
rect 26108 10656 26114 10668
rect 26329 10659 26387 10665
rect 26329 10656 26341 10659
rect 26108 10628 26341 10656
rect 26108 10616 26114 10628
rect 26329 10625 26341 10628
rect 26375 10625 26387 10659
rect 26329 10619 26387 10625
rect 26344 10520 26372 10619
rect 29638 10616 29644 10668
rect 29696 10656 29702 10668
rect 31726 10656 31754 10764
rect 33502 10684 33508 10736
rect 33560 10684 33566 10736
rect 34716 10733 34744 10764
rect 37274 10752 37280 10804
rect 37332 10792 37338 10804
rect 37553 10795 37611 10801
rect 37553 10792 37565 10795
rect 37332 10764 37565 10792
rect 37332 10752 37338 10764
rect 37553 10761 37565 10764
rect 37599 10761 37611 10795
rect 37553 10755 37611 10761
rect 38102 10752 38108 10804
rect 38160 10792 38166 10804
rect 40053 10795 40111 10801
rect 40053 10792 40065 10795
rect 38160 10764 40065 10792
rect 38160 10752 38166 10764
rect 40053 10761 40065 10764
rect 40099 10761 40111 10795
rect 42061 10795 42119 10801
rect 42061 10792 42073 10795
rect 40053 10755 40111 10761
rect 40328 10764 42073 10792
rect 34701 10727 34759 10733
rect 34701 10693 34713 10727
rect 34747 10693 34759 10727
rect 34701 10687 34759 10693
rect 39666 10684 39672 10736
rect 39724 10724 39730 10736
rect 39853 10727 39911 10733
rect 39853 10724 39865 10727
rect 39724 10696 39865 10724
rect 39724 10684 39730 10696
rect 39853 10693 39865 10696
rect 39899 10724 39911 10727
rect 40328 10724 40356 10764
rect 42061 10761 42073 10764
rect 42107 10761 42119 10795
rect 42061 10755 42119 10761
rect 42613 10795 42671 10801
rect 42613 10761 42625 10795
rect 42659 10761 42671 10795
rect 42613 10755 42671 10761
rect 39899 10696 40356 10724
rect 40948 10727 41006 10733
rect 39899 10693 39911 10696
rect 39853 10687 39911 10693
rect 40948 10693 40960 10727
rect 40994 10724 41006 10727
rect 42628 10724 42656 10755
rect 40994 10696 42656 10724
rect 40994 10693 41006 10696
rect 40948 10687 41006 10693
rect 29696 10628 31754 10656
rect 37461 10659 37519 10665
rect 29696 10616 29702 10628
rect 37461 10625 37473 10659
rect 37507 10656 37519 10659
rect 37550 10656 37556 10668
rect 37507 10628 37556 10656
rect 37507 10625 37519 10628
rect 37461 10619 37519 10625
rect 37550 10616 37556 10628
rect 37608 10616 37614 10668
rect 37645 10659 37703 10665
rect 37645 10625 37657 10659
rect 37691 10625 37703 10659
rect 37645 10619 37703 10625
rect 39393 10659 39451 10665
rect 39393 10625 39405 10659
rect 39439 10656 39451 10659
rect 39942 10656 39948 10668
rect 39439 10628 39948 10656
rect 39439 10625 39451 10628
rect 39393 10619 39451 10625
rect 27154 10548 27160 10600
rect 27212 10548 27218 10600
rect 27430 10548 27436 10600
rect 27488 10548 27494 10600
rect 29086 10548 29092 10600
rect 29144 10588 29150 10600
rect 29181 10591 29239 10597
rect 29181 10588 29193 10591
rect 29144 10560 29193 10588
rect 29144 10548 29150 10560
rect 29181 10557 29193 10560
rect 29227 10557 29239 10591
rect 29181 10551 29239 10557
rect 32493 10591 32551 10597
rect 32493 10557 32505 10591
rect 32539 10557 32551 10591
rect 32493 10551 32551 10557
rect 32769 10591 32827 10597
rect 32769 10557 32781 10591
rect 32815 10588 32827 10591
rect 33134 10588 33140 10600
rect 32815 10560 33140 10588
rect 32815 10557 32827 10560
rect 32769 10551 32827 10557
rect 26344 10492 26648 10520
rect 22066 10424 23612 10452
rect 20717 10415 20775 10421
rect 23658 10412 23664 10464
rect 23716 10412 23722 10464
rect 26326 10412 26332 10464
rect 26384 10412 26390 10464
rect 26620 10452 26648 10492
rect 28994 10452 29000 10464
rect 26620 10424 29000 10452
rect 28994 10412 29000 10424
rect 29052 10452 29058 10464
rect 32398 10452 32404 10464
rect 29052 10424 32404 10452
rect 29052 10412 29058 10424
rect 32398 10412 32404 10424
rect 32456 10412 32462 10464
rect 32508 10452 32536 10551
rect 33134 10548 33140 10560
rect 33192 10548 33198 10600
rect 37274 10548 37280 10600
rect 37332 10588 37338 10600
rect 37660 10588 37688 10619
rect 39942 10616 39948 10628
rect 40000 10616 40006 10668
rect 40678 10616 40684 10668
rect 40736 10616 40742 10668
rect 42794 10616 42800 10668
rect 42852 10616 42858 10668
rect 37332 10560 37688 10588
rect 37332 10548 37338 10560
rect 34882 10520 34888 10532
rect 34164 10492 34888 10520
rect 34164 10452 34192 10492
rect 34882 10480 34888 10492
rect 34940 10520 34946 10532
rect 35989 10523 36047 10529
rect 35989 10520 36001 10523
rect 34940 10492 36001 10520
rect 34940 10480 34946 10492
rect 35989 10489 36001 10492
rect 36035 10489 36047 10523
rect 40586 10520 40592 10532
rect 35989 10483 36047 10489
rect 40052 10492 40592 10520
rect 32508 10424 34192 10452
rect 34241 10455 34299 10461
rect 34241 10421 34253 10455
rect 34287 10452 34299 10455
rect 35158 10452 35164 10464
rect 34287 10424 35164 10452
rect 34287 10421 34299 10424
rect 34241 10415 34299 10421
rect 35158 10412 35164 10424
rect 35216 10412 35222 10464
rect 39209 10455 39267 10461
rect 39209 10421 39221 10455
rect 39255 10452 39267 10455
rect 39850 10452 39856 10464
rect 39255 10424 39856 10452
rect 39255 10421 39267 10424
rect 39209 10415 39267 10421
rect 39850 10412 39856 10424
rect 39908 10412 39914 10464
rect 40052 10461 40080 10492
rect 40586 10480 40592 10492
rect 40644 10480 40650 10532
rect 40037 10455 40095 10461
rect 40037 10421 40049 10455
rect 40083 10421 40095 10455
rect 40037 10415 40095 10421
rect 40221 10455 40279 10461
rect 40221 10421 40233 10455
rect 40267 10452 40279 10455
rect 40402 10452 40408 10464
rect 40267 10424 40408 10452
rect 40267 10421 40279 10424
rect 40221 10415 40279 10421
rect 40402 10412 40408 10424
rect 40460 10412 40466 10464
rect 1104 10362 44896 10384
rect 1104 10310 6423 10362
rect 6475 10310 6487 10362
rect 6539 10310 6551 10362
rect 6603 10310 6615 10362
rect 6667 10310 6679 10362
rect 6731 10310 17370 10362
rect 17422 10310 17434 10362
rect 17486 10310 17498 10362
rect 17550 10310 17562 10362
rect 17614 10310 17626 10362
rect 17678 10310 28317 10362
rect 28369 10310 28381 10362
rect 28433 10310 28445 10362
rect 28497 10310 28509 10362
rect 28561 10310 28573 10362
rect 28625 10310 39264 10362
rect 39316 10310 39328 10362
rect 39380 10310 39392 10362
rect 39444 10310 39456 10362
rect 39508 10310 39520 10362
rect 39572 10310 44896 10362
rect 1104 10288 44896 10310
rect 2866 10208 2872 10260
rect 2924 10208 2930 10260
rect 3234 10208 3240 10260
rect 3292 10248 3298 10260
rect 3973 10251 4031 10257
rect 3973 10248 3985 10251
rect 3292 10220 3985 10248
rect 3292 10208 3298 10220
rect 3973 10217 3985 10220
rect 4019 10217 4031 10251
rect 3973 10211 4031 10217
rect 11238 10208 11244 10260
rect 11296 10248 11302 10260
rect 12115 10251 12173 10257
rect 12115 10248 12127 10251
rect 11296 10220 12127 10248
rect 11296 10208 11302 10220
rect 12115 10217 12127 10220
rect 12161 10217 12173 10251
rect 12115 10211 12173 10217
rect 14274 10208 14280 10260
rect 14332 10248 14338 10260
rect 16022 10248 16028 10260
rect 14332 10220 16028 10248
rect 14332 10208 14338 10220
rect 16022 10208 16028 10220
rect 16080 10208 16086 10260
rect 16482 10208 16488 10260
rect 16540 10208 16546 10260
rect 18693 10251 18751 10257
rect 18693 10217 18705 10251
rect 18739 10248 18751 10251
rect 18874 10248 18880 10260
rect 18739 10220 18880 10248
rect 18739 10217 18751 10220
rect 18693 10211 18751 10217
rect 18874 10208 18880 10220
rect 18932 10208 18938 10260
rect 20898 10208 20904 10260
rect 20956 10248 20962 10260
rect 22833 10251 22891 10257
rect 22833 10248 22845 10251
rect 20956 10220 22845 10248
rect 20956 10208 20962 10220
rect 22833 10217 22845 10220
rect 22879 10217 22891 10251
rect 22833 10211 22891 10217
rect 26145 10251 26203 10257
rect 26145 10217 26157 10251
rect 26191 10248 26203 10251
rect 26418 10248 26424 10260
rect 26191 10220 26424 10248
rect 26191 10217 26203 10220
rect 26145 10211 26203 10217
rect 26418 10208 26424 10220
rect 26476 10208 26482 10260
rect 26786 10208 26792 10260
rect 26844 10208 26850 10260
rect 28166 10208 28172 10260
rect 28224 10248 28230 10260
rect 28261 10251 28319 10257
rect 28261 10248 28273 10251
rect 28224 10220 28273 10248
rect 28224 10208 28230 10220
rect 28261 10217 28273 10220
rect 28307 10217 28319 10251
rect 28261 10211 28319 10217
rect 30561 10251 30619 10257
rect 30561 10217 30573 10251
rect 30607 10248 30619 10251
rect 30834 10248 30840 10260
rect 30607 10220 30840 10248
rect 30607 10217 30619 10220
rect 30561 10211 30619 10217
rect 30834 10208 30840 10220
rect 30892 10208 30898 10260
rect 31404 10220 33548 10248
rect 11514 10140 11520 10192
rect 11572 10180 11578 10192
rect 13081 10183 13139 10189
rect 13081 10180 13093 10183
rect 11572 10152 13093 10180
rect 11572 10140 11578 10152
rect 13081 10149 13093 10152
rect 13127 10149 13139 10183
rect 13081 10143 13139 10149
rect 14200 10152 14504 10180
rect 4614 10072 4620 10124
rect 4672 10112 4678 10124
rect 5810 10112 5816 10124
rect 4672 10084 5816 10112
rect 4672 10072 4678 10084
rect 5810 10072 5816 10084
rect 5868 10072 5874 10124
rect 10318 10072 10324 10124
rect 10376 10072 10382 10124
rect 10686 10072 10692 10124
rect 10744 10072 10750 10124
rect 14200 10112 14228 10152
rect 10796 10084 14228 10112
rect 14476 10112 14504 10152
rect 14826 10140 14832 10192
rect 14884 10180 14890 10192
rect 18598 10180 18604 10192
rect 14884 10152 18604 10180
rect 14884 10140 14890 10152
rect 18598 10140 18604 10152
rect 18656 10140 18662 10192
rect 21726 10140 21732 10192
rect 21784 10180 21790 10192
rect 22738 10180 22744 10192
rect 21784 10152 22744 10180
rect 21784 10140 21790 10152
rect 22738 10140 22744 10152
rect 22796 10180 22802 10192
rect 22796 10152 23428 10180
rect 22796 10140 22802 10152
rect 16574 10112 16580 10124
rect 14476 10084 16580 10112
rect 3053 10047 3111 10053
rect 3053 10013 3065 10047
rect 3099 10044 3111 10047
rect 3970 10044 3976 10056
rect 3099 10016 3976 10044
rect 3099 10013 3111 10016
rect 3053 10007 3111 10013
rect 3970 10004 3976 10016
rect 4028 10004 4034 10056
rect 4338 10004 4344 10056
rect 4396 10004 4402 10056
rect 6270 10004 6276 10056
rect 6328 10044 6334 10056
rect 6549 10047 6607 10053
rect 6549 10044 6561 10047
rect 6328 10016 6561 10044
rect 6328 10004 6334 10016
rect 6549 10013 6561 10016
rect 6595 10013 6607 10047
rect 6549 10007 6607 10013
rect 6816 10047 6874 10053
rect 6816 10013 6828 10047
rect 6862 10044 6874 10047
rect 10796 10044 10824 10084
rect 16574 10072 16580 10084
rect 16632 10072 16638 10124
rect 17770 10072 17776 10124
rect 17828 10112 17834 10124
rect 20533 10115 20591 10121
rect 17828 10084 19932 10112
rect 17828 10072 17834 10084
rect 6862 10016 10824 10044
rect 6862 10013 6874 10016
rect 6816 10007 6874 10013
rect 12434 10004 12440 10056
rect 12492 10044 12498 10056
rect 12989 10047 13047 10053
rect 12989 10044 13001 10047
rect 12492 10016 13001 10044
rect 12492 10004 12498 10016
rect 12989 10013 13001 10016
rect 13035 10013 13047 10047
rect 12989 10007 13047 10013
rect 13170 10004 13176 10056
rect 13228 10044 13234 10056
rect 13446 10044 13452 10056
rect 13228 10016 13452 10044
rect 13228 10004 13234 10016
rect 13446 10004 13452 10016
rect 13504 10004 13510 10056
rect 14274 10004 14280 10056
rect 14332 10004 14338 10056
rect 14369 10047 14427 10053
rect 14369 10013 14381 10047
rect 14415 10044 14427 10047
rect 15105 10047 15163 10053
rect 15105 10044 15117 10047
rect 14415 10016 15117 10044
rect 14415 10013 14427 10016
rect 14369 10007 14427 10013
rect 15105 10013 15117 10016
rect 15151 10013 15163 10047
rect 15105 10007 15163 10013
rect 16669 10047 16727 10053
rect 16669 10013 16681 10047
rect 16715 10044 16727 10047
rect 16715 10016 17172 10044
rect 16715 10013 16727 10016
rect 16669 10007 16727 10013
rect 11730 9948 14964 9976
rect 4430 9868 4436 9920
rect 4488 9868 4494 9920
rect 7926 9868 7932 9920
rect 7984 9868 7990 9920
rect 12342 9868 12348 9920
rect 12400 9908 12406 9920
rect 14826 9908 14832 9920
rect 12400 9880 14832 9908
rect 12400 9868 12406 9880
rect 14826 9868 14832 9880
rect 14884 9868 14890 9920
rect 14936 9917 14964 9948
rect 17144 9917 17172 10016
rect 17218 10004 17224 10056
rect 17276 10044 17282 10056
rect 17497 10047 17555 10053
rect 17497 10044 17509 10047
rect 17276 10016 17509 10044
rect 17276 10004 17282 10016
rect 17497 10013 17509 10016
rect 17543 10013 17555 10047
rect 17497 10007 17555 10013
rect 17589 10047 17647 10053
rect 17589 10013 17601 10047
rect 17635 10044 17647 10047
rect 17954 10044 17960 10056
rect 17635 10016 17960 10044
rect 17635 10013 17647 10016
rect 17589 10007 17647 10013
rect 17954 10004 17960 10016
rect 18012 10004 18018 10056
rect 18322 10004 18328 10056
rect 18380 10004 18386 10056
rect 18506 10004 18512 10056
rect 18564 10004 18570 10056
rect 19702 10004 19708 10056
rect 19760 10004 19766 10056
rect 14921 9911 14979 9917
rect 14921 9877 14933 9911
rect 14967 9877 14979 9911
rect 14921 9871 14979 9877
rect 17129 9911 17187 9917
rect 17129 9877 17141 9911
rect 17175 9877 17187 9911
rect 18340 9908 18368 10004
rect 19242 9908 19248 9920
rect 18340 9880 19248 9908
rect 17129 9871 17187 9877
rect 19242 9868 19248 9880
rect 19300 9908 19306 9920
rect 19797 9911 19855 9917
rect 19797 9908 19809 9911
rect 19300 9880 19809 9908
rect 19300 9868 19306 9880
rect 19797 9877 19809 9880
rect 19843 9877 19855 9911
rect 19904 9908 19932 10084
rect 20533 10081 20545 10115
rect 20579 10112 20591 10115
rect 22186 10112 22192 10124
rect 20579 10084 22192 10112
rect 20579 10081 20591 10084
rect 20533 10075 20591 10081
rect 22186 10072 22192 10084
rect 22244 10072 22250 10124
rect 23400 10121 23428 10152
rect 30466 10140 30472 10192
rect 30524 10180 30530 10192
rect 31113 10183 31171 10189
rect 31113 10180 31125 10183
rect 30524 10152 31125 10180
rect 30524 10140 30530 10152
rect 31113 10149 31125 10152
rect 31159 10149 31171 10183
rect 31113 10143 31171 10149
rect 23385 10115 23443 10121
rect 23385 10081 23397 10115
rect 23431 10081 23443 10115
rect 27614 10112 27620 10124
rect 23385 10075 23443 10081
rect 26988 10084 27620 10112
rect 20806 10004 20812 10056
rect 20864 10044 20870 10056
rect 20901 10047 20959 10053
rect 20901 10044 20913 10047
rect 20864 10016 20913 10044
rect 20864 10004 20870 10016
rect 20901 10013 20913 10016
rect 20947 10013 20959 10047
rect 20901 10007 20959 10013
rect 23198 10004 23204 10056
rect 23256 10004 23262 10056
rect 26326 10004 26332 10056
rect 26384 10004 26390 10056
rect 26988 10053 27016 10084
rect 27614 10072 27620 10084
rect 27672 10072 27678 10124
rect 27890 10112 27896 10124
rect 27724 10084 27896 10112
rect 27724 10053 27752 10084
rect 27890 10072 27896 10084
rect 27948 10112 27954 10124
rect 28166 10112 28172 10124
rect 27948 10084 28172 10112
rect 27948 10072 27954 10084
rect 28166 10072 28172 10084
rect 28224 10072 28230 10124
rect 30484 10084 31340 10112
rect 26973 10047 27031 10053
rect 26973 10013 26985 10047
rect 27019 10013 27031 10047
rect 26973 10007 27031 10013
rect 27709 10047 27767 10053
rect 27709 10013 27721 10047
rect 27755 10013 27767 10047
rect 27709 10007 27767 10013
rect 27801 10047 27859 10053
rect 27801 10013 27813 10047
rect 27847 10044 27859 10047
rect 28445 10047 28503 10053
rect 28445 10044 28457 10047
rect 27847 10016 28457 10044
rect 27847 10013 27859 10016
rect 27801 10007 27859 10013
rect 28445 10013 28457 10016
rect 28491 10013 28503 10047
rect 28445 10007 28503 10013
rect 28994 10004 29000 10056
rect 29052 10044 29058 10056
rect 29917 10047 29975 10053
rect 29917 10044 29929 10047
rect 29052 10016 29929 10044
rect 29052 10004 29058 10016
rect 29917 10013 29929 10016
rect 29963 10013 29975 10047
rect 29917 10007 29975 10013
rect 30374 10004 30380 10056
rect 30432 10044 30438 10056
rect 30484 10053 30512 10084
rect 31312 10056 31340 10084
rect 30469 10047 30527 10053
rect 30469 10044 30481 10047
rect 30432 10016 30481 10044
rect 30432 10004 30438 10016
rect 30469 10013 30481 10016
rect 30515 10013 30527 10047
rect 30653 10047 30711 10053
rect 30653 10046 30665 10047
rect 30469 10007 30527 10013
rect 30576 10018 30665 10046
rect 21266 9936 21272 9988
rect 21324 9936 21330 9988
rect 30282 9936 30288 9988
rect 30340 9976 30346 9988
rect 30576 9976 30604 10018
rect 30653 10013 30665 10018
rect 30699 10013 30711 10047
rect 30653 10007 30711 10013
rect 31294 10004 31300 10056
rect 31352 10004 31358 10056
rect 31404 10053 31432 10220
rect 33520 10180 33548 10220
rect 33594 10208 33600 10260
rect 33652 10208 33658 10260
rect 36354 10248 36360 10260
rect 34992 10220 36360 10248
rect 34992 10180 35020 10220
rect 36354 10208 36360 10220
rect 36412 10208 36418 10260
rect 38289 10251 38347 10257
rect 38289 10217 38301 10251
rect 38335 10248 38347 10251
rect 39758 10248 39764 10260
rect 38335 10220 39764 10248
rect 38335 10217 38347 10220
rect 38289 10211 38347 10217
rect 39758 10208 39764 10220
rect 39816 10208 39822 10260
rect 39942 10208 39948 10260
rect 40000 10248 40006 10260
rect 40037 10251 40095 10257
rect 40037 10248 40049 10251
rect 40000 10220 40049 10248
rect 40000 10208 40006 10220
rect 40037 10217 40049 10220
rect 40083 10217 40095 10251
rect 40037 10211 40095 10217
rect 40310 10208 40316 10260
rect 40368 10248 40374 10260
rect 40368 10220 41920 10248
rect 40368 10208 40374 10220
rect 40494 10180 40500 10192
rect 33520 10152 35020 10180
rect 39132 10152 40500 10180
rect 31757 10115 31815 10121
rect 31757 10081 31769 10115
rect 31803 10112 31815 10115
rect 31846 10112 31852 10124
rect 31803 10084 31852 10112
rect 31803 10081 31815 10084
rect 31757 10075 31815 10081
rect 31846 10072 31852 10084
rect 31904 10072 31910 10124
rect 32214 10072 32220 10124
rect 32272 10112 32278 10124
rect 32493 10115 32551 10121
rect 32493 10112 32505 10115
rect 32272 10084 32505 10112
rect 32272 10072 32278 10084
rect 32493 10081 32505 10084
rect 32539 10081 32551 10115
rect 32493 10075 32551 10081
rect 34882 10072 34888 10124
rect 34940 10072 34946 10124
rect 35158 10072 35164 10124
rect 35216 10072 35222 10124
rect 35894 10072 35900 10124
rect 35952 10112 35958 10124
rect 37182 10112 37188 10124
rect 35952 10084 37188 10112
rect 35952 10072 35958 10084
rect 37182 10072 37188 10084
rect 37240 10072 37246 10124
rect 37550 10072 37556 10124
rect 37608 10072 37614 10124
rect 39132 10121 39160 10152
rect 40494 10140 40500 10152
rect 40552 10140 40558 10192
rect 41892 10180 41920 10220
rect 42794 10208 42800 10260
rect 42852 10208 42858 10260
rect 41892 10152 43116 10180
rect 39117 10115 39175 10121
rect 39117 10081 39129 10115
rect 39163 10081 39175 10115
rect 39117 10075 39175 10081
rect 39850 10072 39856 10124
rect 39908 10112 39914 10124
rect 39908 10084 40632 10112
rect 39908 10072 39914 10084
rect 31389 10047 31447 10053
rect 31389 10013 31401 10047
rect 31435 10013 31447 10047
rect 31389 10007 31447 10013
rect 31496 10016 31754 10044
rect 30340 9948 30604 9976
rect 30340 9936 30346 9948
rect 20990 9908 20996 9920
rect 19904 9880 20996 9908
rect 19797 9871 19855 9877
rect 20990 9868 20996 9880
rect 21048 9868 21054 9920
rect 21174 9868 21180 9920
rect 21232 9908 21238 9920
rect 22327 9911 22385 9917
rect 22327 9908 22339 9911
rect 21232 9880 22339 9908
rect 21232 9868 21238 9880
rect 22327 9877 22339 9880
rect 22373 9877 22385 9911
rect 22327 9871 22385 9877
rect 23293 9911 23351 9917
rect 23293 9877 23305 9911
rect 23339 9908 23351 9911
rect 23474 9908 23480 9920
rect 23339 9880 23480 9908
rect 23339 9877 23351 9880
rect 23293 9871 23351 9877
rect 23474 9868 23480 9880
rect 23532 9868 23538 9920
rect 29546 9868 29552 9920
rect 29604 9908 29610 9920
rect 29733 9911 29791 9917
rect 29733 9908 29745 9911
rect 29604 9880 29745 9908
rect 29604 9868 29610 9880
rect 29733 9877 29745 9880
rect 29779 9877 29791 9911
rect 30576 9908 30604 9948
rect 31110 9936 31116 9988
rect 31168 9976 31174 9988
rect 31496 9985 31524 10016
rect 31481 9979 31539 9985
rect 31481 9976 31493 9979
rect 31168 9948 31493 9976
rect 31168 9936 31174 9948
rect 31481 9945 31493 9948
rect 31527 9945 31539 9979
rect 31481 9939 31539 9945
rect 31570 9936 31576 9988
rect 31628 9985 31634 9988
rect 31628 9979 31657 9985
rect 31645 9945 31657 9979
rect 31726 9976 31754 10016
rect 32398 10004 32404 10056
rect 32456 10044 32462 10056
rect 33597 10047 33655 10053
rect 33597 10044 33609 10047
rect 32456 10016 33609 10044
rect 32456 10004 32462 10016
rect 33597 10013 33609 10016
rect 33643 10044 33655 10047
rect 33686 10044 33692 10056
rect 33643 10016 33692 10044
rect 33643 10013 33655 10016
rect 33597 10007 33655 10013
rect 33686 10004 33692 10016
rect 33744 10004 33750 10056
rect 34333 10047 34391 10053
rect 34333 10013 34345 10047
rect 34379 10044 34391 10047
rect 34514 10044 34520 10056
rect 34379 10016 34520 10044
rect 34379 10013 34391 10016
rect 34333 10007 34391 10013
rect 34514 10004 34520 10016
rect 34572 10004 34578 10056
rect 36722 10004 36728 10056
rect 36780 10044 36786 10056
rect 37369 10047 37427 10053
rect 37369 10044 37381 10047
rect 36780 10016 37381 10044
rect 36780 10004 36786 10016
rect 37369 10013 37381 10016
rect 37415 10013 37427 10047
rect 37369 10007 37427 10013
rect 37642 10004 37648 10056
rect 37700 10004 37706 10056
rect 38102 10004 38108 10056
rect 38160 10004 38166 10056
rect 39301 10047 39359 10053
rect 39301 10013 39313 10047
rect 39347 10013 39359 10047
rect 39301 10007 39359 10013
rect 34790 9976 34796 9988
rect 31726 9948 34796 9976
rect 31628 9939 31657 9945
rect 31628 9936 31634 9939
rect 34790 9936 34796 9948
rect 34848 9936 34854 9988
rect 39316 9976 39344 10007
rect 40218 10004 40224 10056
rect 40276 10004 40282 10056
rect 40402 10004 40408 10056
rect 40460 10004 40466 10056
rect 40494 10004 40500 10056
rect 40552 10004 40558 10056
rect 40604 10044 40632 10084
rect 40678 10072 40684 10124
rect 40736 10112 40742 10124
rect 43088 10121 43116 10152
rect 40957 10115 41015 10121
rect 40957 10112 40969 10115
rect 40736 10084 40969 10112
rect 40736 10072 40742 10084
rect 40957 10081 40969 10084
rect 41003 10081 41015 10115
rect 40957 10075 41015 10081
rect 43073 10115 43131 10121
rect 43073 10081 43085 10115
rect 43119 10081 43131 10115
rect 43073 10075 43131 10081
rect 41213 10047 41271 10053
rect 41213 10044 41225 10047
rect 40604 10016 41225 10044
rect 41213 10013 41225 10016
rect 41259 10013 41271 10047
rect 41213 10007 41271 10013
rect 42797 10047 42855 10053
rect 42797 10013 42809 10047
rect 42843 10013 42855 10047
rect 42797 10007 42855 10013
rect 40420 9976 40448 10004
rect 42812 9976 42840 10007
rect 42886 10004 42892 10056
rect 42944 10004 42950 10056
rect 35268 9948 35650 9976
rect 39316 9948 42840 9976
rect 32950 9908 32956 9920
rect 30576 9880 32956 9908
rect 29733 9871 29791 9877
rect 32950 9868 32956 9880
rect 33008 9868 33014 9920
rect 34149 9911 34207 9917
rect 34149 9877 34161 9911
rect 34195 9908 34207 9911
rect 35268 9908 35296 9948
rect 34195 9880 35296 9908
rect 34195 9877 34207 9880
rect 34149 9871 34207 9877
rect 35986 9868 35992 9920
rect 36044 9908 36050 9920
rect 36633 9911 36691 9917
rect 36633 9908 36645 9911
rect 36044 9880 36645 9908
rect 36044 9868 36050 9880
rect 36633 9877 36645 9880
rect 36679 9877 36691 9911
rect 36633 9871 36691 9877
rect 39485 9911 39543 9917
rect 39485 9877 39497 9911
rect 39531 9908 39543 9911
rect 40034 9908 40040 9920
rect 39531 9880 40040 9908
rect 39531 9877 39543 9880
rect 39485 9871 39543 9877
rect 40034 9868 40040 9880
rect 40092 9868 40098 9920
rect 40494 9868 40500 9920
rect 40552 9908 40558 9920
rect 40954 9908 40960 9920
rect 40552 9880 40960 9908
rect 40552 9868 40558 9880
rect 40954 9868 40960 9880
rect 41012 9908 41018 9920
rect 42337 9911 42395 9917
rect 42337 9908 42349 9911
rect 41012 9880 42349 9908
rect 41012 9868 41018 9880
rect 42337 9877 42349 9880
rect 42383 9877 42395 9911
rect 42337 9871 42395 9877
rect 1104 9818 45051 9840
rect 1104 9766 11896 9818
rect 11948 9766 11960 9818
rect 12012 9766 12024 9818
rect 12076 9766 12088 9818
rect 12140 9766 12152 9818
rect 12204 9766 22843 9818
rect 22895 9766 22907 9818
rect 22959 9766 22971 9818
rect 23023 9766 23035 9818
rect 23087 9766 23099 9818
rect 23151 9766 33790 9818
rect 33842 9766 33854 9818
rect 33906 9766 33918 9818
rect 33970 9766 33982 9818
rect 34034 9766 34046 9818
rect 34098 9766 44737 9818
rect 44789 9766 44801 9818
rect 44853 9766 44865 9818
rect 44917 9766 44929 9818
rect 44981 9766 44993 9818
rect 45045 9766 45051 9818
rect 1104 9744 45051 9766
rect 13446 9664 13452 9716
rect 13504 9664 13510 9716
rect 13538 9664 13544 9716
rect 13596 9704 13602 9716
rect 17770 9704 17776 9716
rect 13596 9676 17776 9704
rect 13596 9664 13602 9676
rect 17770 9664 17776 9676
rect 17828 9664 17834 9716
rect 22002 9704 22008 9716
rect 20180 9676 22008 9704
rect 2498 9596 2504 9648
rect 2556 9636 2562 9648
rect 5721 9639 5779 9645
rect 2556 9608 3556 9636
rect 2556 9596 2562 9608
rect 2768 9571 2826 9577
rect 2768 9537 2780 9571
rect 2814 9568 2826 9571
rect 3142 9568 3148 9580
rect 2814 9540 3148 9568
rect 2814 9537 2826 9540
rect 2768 9531 2826 9537
rect 3142 9528 3148 9540
rect 3200 9528 3206 9580
rect 2501 9503 2559 9509
rect 2501 9469 2513 9503
rect 2547 9469 2559 9503
rect 3528 9500 3556 9608
rect 5721 9605 5733 9639
rect 5767 9636 5779 9639
rect 6794 9639 6852 9645
rect 6794 9636 6806 9639
rect 5767 9608 6806 9636
rect 5767 9605 5779 9608
rect 5721 9599 5779 9605
rect 6794 9605 6806 9608
rect 6840 9636 6852 9639
rect 7926 9636 7932 9648
rect 6840 9608 7932 9636
rect 6840 9605 6852 9608
rect 6794 9599 6852 9605
rect 7926 9596 7932 9608
rect 7984 9596 7990 9648
rect 10781 9639 10839 9645
rect 10781 9605 10793 9639
rect 10827 9636 10839 9639
rect 12250 9636 12256 9648
rect 10827 9608 12256 9636
rect 10827 9605 10839 9608
rect 10781 9599 10839 9605
rect 12250 9596 12256 9608
rect 12308 9596 12314 9648
rect 13262 9596 13268 9648
rect 13320 9636 13326 9648
rect 13320 9608 17908 9636
rect 13320 9596 13326 9608
rect 5626 9528 5632 9580
rect 5684 9528 5690 9580
rect 10686 9568 10692 9580
rect 5736 9540 10692 9568
rect 5736 9500 5764 9540
rect 10686 9528 10692 9540
rect 10744 9528 10750 9580
rect 13078 9528 13084 9580
rect 13136 9528 13142 9580
rect 13354 9528 13360 9580
rect 13412 9568 13418 9580
rect 13412 9540 14044 9568
rect 13412 9528 13418 9540
rect 3528 9472 5764 9500
rect 2501 9463 2559 9469
rect 2516 9364 2544 9463
rect 5810 9460 5816 9512
rect 5868 9460 5874 9512
rect 6270 9460 6276 9512
rect 6328 9500 6334 9512
rect 6549 9503 6607 9509
rect 6549 9500 6561 9503
rect 6328 9472 6561 9500
rect 6328 9460 6334 9472
rect 6549 9469 6561 9472
rect 6595 9469 6607 9503
rect 6549 9463 6607 9469
rect 10870 9460 10876 9512
rect 10928 9460 10934 9512
rect 10962 9460 10968 9512
rect 11020 9460 11026 9512
rect 11701 9503 11759 9509
rect 11701 9469 11713 9503
rect 11747 9469 11759 9503
rect 11701 9463 11759 9469
rect 11977 9503 12035 9509
rect 11977 9469 11989 9503
rect 12023 9500 12035 9503
rect 14016 9500 14044 9540
rect 14090 9528 14096 9580
rect 14148 9528 14154 9580
rect 17126 9577 17132 9580
rect 15177 9571 15235 9577
rect 15177 9568 15189 9571
rect 14200 9540 15189 9568
rect 14200 9500 14228 9540
rect 15177 9537 15189 9540
rect 15223 9537 15235 9571
rect 17120 9568 17132 9577
rect 17087 9540 17132 9568
rect 15177 9531 15235 9537
rect 17120 9531 17132 9540
rect 17126 9528 17132 9531
rect 17184 9528 17190 9580
rect 12023 9472 13952 9500
rect 14016 9472 14228 9500
rect 12023 9469 12035 9472
rect 11977 9463 12035 9469
rect 3878 9392 3884 9444
rect 3936 9392 3942 9444
rect 7650 9392 7656 9444
rect 7708 9432 7714 9444
rect 7929 9435 7987 9441
rect 7929 9432 7941 9435
rect 7708 9404 7941 9432
rect 7708 9392 7714 9404
rect 7929 9401 7941 9404
rect 7975 9401 7987 9435
rect 7929 9395 7987 9401
rect 2774 9364 2780 9376
rect 2516 9336 2780 9364
rect 2774 9324 2780 9336
rect 2832 9324 2838 9376
rect 5261 9367 5319 9373
rect 5261 9333 5273 9367
rect 5307 9364 5319 9367
rect 6178 9364 6184 9376
rect 5307 9336 6184 9364
rect 5307 9333 5319 9336
rect 5261 9327 5319 9333
rect 6178 9324 6184 9336
rect 6236 9324 6242 9376
rect 10413 9367 10471 9373
rect 10413 9333 10425 9367
rect 10459 9364 10471 9367
rect 11146 9364 11152 9376
rect 10459 9336 11152 9364
rect 10459 9333 10471 9336
rect 10413 9327 10471 9333
rect 11146 9324 11152 9336
rect 11204 9324 11210 9376
rect 11716 9364 11744 9463
rect 12986 9392 12992 9444
rect 13044 9432 13050 9444
rect 13354 9432 13360 9444
rect 13044 9404 13360 9432
rect 13044 9392 13050 9404
rect 13354 9392 13360 9404
rect 13412 9392 13418 9444
rect 13814 9364 13820 9376
rect 11716 9336 13820 9364
rect 13814 9324 13820 9336
rect 13872 9324 13878 9376
rect 13924 9373 13952 9472
rect 14918 9460 14924 9512
rect 14976 9460 14982 9512
rect 16850 9460 16856 9512
rect 16908 9460 16914 9512
rect 13998 9392 14004 9444
rect 14056 9432 14062 9444
rect 14936 9432 14964 9460
rect 14056 9404 14964 9432
rect 14056 9392 14062 9404
rect 16298 9392 16304 9444
rect 16356 9392 16362 9444
rect 17880 9432 17908 9608
rect 20180 9577 20208 9676
rect 22002 9664 22008 9676
rect 22060 9664 22066 9716
rect 27157 9707 27215 9713
rect 23768 9676 23980 9704
rect 20806 9596 20812 9648
rect 20864 9636 20870 9648
rect 23768 9636 23796 9676
rect 20864 9608 23796 9636
rect 20864 9596 20870 9608
rect 23842 9596 23848 9648
rect 23900 9636 23906 9648
rect 23952 9636 23980 9676
rect 27157 9673 27169 9707
rect 27203 9704 27215 9707
rect 27430 9704 27436 9716
rect 27203 9676 27436 9704
rect 27203 9673 27215 9676
rect 27157 9667 27215 9673
rect 27430 9664 27436 9676
rect 27488 9664 27494 9716
rect 31294 9664 31300 9716
rect 31352 9704 31358 9716
rect 31662 9704 31668 9716
rect 31352 9676 31668 9704
rect 31352 9664 31358 9676
rect 31662 9664 31668 9676
rect 31720 9704 31726 9716
rect 35894 9704 35900 9716
rect 31720 9676 35900 9704
rect 31720 9664 31726 9676
rect 35894 9664 35900 9676
rect 35952 9664 35958 9716
rect 36354 9664 36360 9716
rect 36412 9704 36418 9716
rect 39666 9704 39672 9716
rect 36412 9676 37596 9704
rect 36412 9664 36418 9676
rect 29638 9636 29644 9648
rect 23900 9608 23980 9636
rect 24136 9608 29644 9636
rect 23900 9596 23906 9608
rect 19521 9571 19579 9577
rect 19521 9537 19533 9571
rect 19567 9537 19579 9571
rect 19521 9531 19579 9537
rect 20165 9571 20223 9577
rect 20165 9537 20177 9571
rect 20211 9537 20223 9571
rect 20165 9531 20223 9537
rect 19536 9500 19564 9531
rect 21082 9528 21088 9580
rect 21140 9528 21146 9580
rect 21174 9528 21180 9580
rect 21232 9568 21238 9580
rect 22094 9568 22100 9580
rect 21232 9540 22100 9568
rect 21232 9528 21238 9540
rect 22094 9528 22100 9540
rect 22152 9528 22158 9580
rect 22189 9571 22247 9577
rect 22189 9537 22201 9571
rect 22235 9568 22247 9571
rect 23290 9568 23296 9580
rect 22235 9540 23296 9568
rect 22235 9537 22247 9540
rect 22189 9531 22247 9537
rect 23290 9528 23296 9540
rect 23348 9528 23354 9580
rect 20898 9500 20904 9512
rect 19536 9472 20904 9500
rect 20898 9460 20904 9472
rect 20956 9460 20962 9512
rect 20990 9460 20996 9512
rect 21048 9500 21054 9512
rect 21361 9503 21419 9509
rect 21361 9500 21373 9503
rect 21048 9472 21373 9500
rect 21048 9460 21054 9472
rect 21361 9469 21373 9472
rect 21407 9500 21419 9503
rect 21726 9500 21732 9512
rect 21407 9472 21732 9500
rect 21407 9469 21419 9472
rect 21361 9463 21419 9469
rect 21726 9460 21732 9472
rect 21784 9460 21790 9512
rect 23845 9503 23903 9509
rect 23845 9500 23857 9503
rect 22204 9472 23857 9500
rect 22204 9432 22232 9472
rect 23845 9469 23857 9472
rect 23891 9500 23903 9503
rect 24136 9500 24164 9608
rect 29638 9596 29644 9608
rect 29696 9596 29702 9648
rect 32858 9596 32864 9648
rect 32916 9636 32922 9648
rect 35158 9636 35164 9648
rect 32916 9608 33456 9636
rect 32916 9596 32922 9608
rect 33428 9580 33456 9608
rect 34716 9608 35164 9636
rect 25222 9528 25228 9580
rect 25280 9528 25286 9580
rect 26326 9528 26332 9580
rect 26384 9568 26390 9580
rect 26421 9571 26479 9577
rect 26421 9568 26433 9571
rect 26384 9540 26433 9568
rect 26384 9528 26390 9540
rect 26421 9537 26433 9540
rect 26467 9537 26479 9571
rect 26421 9531 26479 9537
rect 27338 9528 27344 9580
rect 27396 9528 27402 9580
rect 27982 9528 27988 9580
rect 28040 9528 28046 9580
rect 28074 9528 28080 9580
rect 28132 9568 28138 9580
rect 28445 9571 28503 9577
rect 28445 9568 28457 9571
rect 28132 9540 28457 9568
rect 28132 9528 28138 9540
rect 28445 9537 28457 9540
rect 28491 9537 28503 9571
rect 28445 9531 28503 9537
rect 28629 9571 28687 9577
rect 28629 9537 28641 9571
rect 28675 9568 28687 9571
rect 29178 9568 29184 9580
rect 28675 9540 29184 9568
rect 28675 9537 28687 9540
rect 28629 9531 28687 9537
rect 29178 9528 29184 9540
rect 29236 9528 29242 9580
rect 29546 9577 29552 9580
rect 29540 9568 29552 9577
rect 29507 9540 29552 9568
rect 29540 9531 29552 9540
rect 29546 9528 29552 9531
rect 29604 9528 29610 9580
rect 31110 9528 31116 9580
rect 31168 9528 31174 9580
rect 31294 9528 31300 9580
rect 31352 9528 31358 9580
rect 32214 9528 32220 9580
rect 32272 9568 32278 9580
rect 32585 9571 32643 9577
rect 32585 9568 32597 9571
rect 32272 9540 32597 9568
rect 32272 9528 32278 9540
rect 32585 9537 32597 9540
rect 32631 9537 32643 9571
rect 32585 9531 32643 9537
rect 32950 9528 32956 9580
rect 33008 9568 33014 9580
rect 33229 9571 33287 9577
rect 33229 9568 33241 9571
rect 33008 9540 33241 9568
rect 33008 9528 33014 9540
rect 33229 9537 33241 9540
rect 33275 9537 33287 9571
rect 33229 9531 33287 9537
rect 33410 9528 33416 9580
rect 33468 9528 33474 9580
rect 34716 9577 34744 9608
rect 35158 9596 35164 9608
rect 35216 9636 35222 9648
rect 37568 9645 37596 9676
rect 39408 9676 39672 9704
rect 39408 9645 39436 9676
rect 39666 9664 39672 9676
rect 39724 9704 39730 9716
rect 39942 9704 39948 9716
rect 39724 9676 39948 9704
rect 39724 9664 39730 9676
rect 39942 9664 39948 9676
rect 40000 9664 40006 9716
rect 40405 9707 40463 9713
rect 40405 9673 40417 9707
rect 40451 9704 40463 9707
rect 40494 9704 40500 9716
rect 40451 9676 40500 9704
rect 40451 9673 40463 9676
rect 40405 9667 40463 9673
rect 40494 9664 40500 9676
rect 40552 9664 40558 9716
rect 35989 9639 36047 9645
rect 35216 9608 35848 9636
rect 35216 9596 35222 9608
rect 35820 9577 35848 9608
rect 35989 9605 36001 9639
rect 36035 9636 36047 9639
rect 37553 9639 37611 9645
rect 36035 9608 36768 9636
rect 36035 9605 36047 9608
rect 35989 9599 36047 9605
rect 36740 9580 36768 9608
rect 37553 9605 37565 9639
rect 37599 9605 37611 9639
rect 37553 9599 37611 9605
rect 39393 9639 39451 9645
rect 39393 9605 39405 9639
rect 39439 9605 39451 9639
rect 42886 9636 42892 9648
rect 39393 9599 39451 9605
rect 39500 9608 42892 9636
rect 34701 9571 34759 9577
rect 34701 9537 34713 9571
rect 34747 9537 34759 9571
rect 34701 9531 34759 9537
rect 34885 9571 34943 9577
rect 34885 9537 34897 9571
rect 34931 9568 34943 9571
rect 35713 9571 35771 9577
rect 35713 9568 35725 9571
rect 34931 9540 35725 9568
rect 34931 9537 34943 9540
rect 34885 9531 34943 9537
rect 35713 9537 35725 9540
rect 35759 9537 35771 9571
rect 35713 9531 35771 9537
rect 35805 9571 35863 9577
rect 35805 9537 35817 9571
rect 35851 9537 35863 9571
rect 35805 9531 35863 9537
rect 36449 9571 36507 9577
rect 36449 9537 36461 9571
rect 36495 9537 36507 9571
rect 36449 9531 36507 9537
rect 23891 9472 24164 9500
rect 28813 9503 28871 9509
rect 23891 9469 23903 9472
rect 23845 9463 23903 9469
rect 28813 9469 28825 9503
rect 28859 9500 28871 9503
rect 28994 9500 29000 9512
rect 28859 9472 29000 9500
rect 28859 9469 28871 9472
rect 28813 9463 28871 9469
rect 28994 9460 29000 9472
rect 29052 9460 29058 9512
rect 29270 9460 29276 9512
rect 29328 9460 29334 9512
rect 33321 9503 33379 9509
rect 33321 9469 33333 9503
rect 33367 9500 33379 9503
rect 34900 9500 34928 9531
rect 33367 9472 34928 9500
rect 35345 9503 35403 9509
rect 33367 9469 33379 9472
rect 33321 9463 33379 9469
rect 35345 9469 35357 9503
rect 35391 9500 35403 9503
rect 36354 9500 36360 9512
rect 35391 9472 36360 9500
rect 35391 9469 35403 9472
rect 35345 9463 35403 9469
rect 36354 9460 36360 9472
rect 36412 9460 36418 9512
rect 27706 9432 27712 9444
rect 17880 9404 22232 9432
rect 22296 9404 27712 9432
rect 13909 9367 13967 9373
rect 13909 9333 13921 9367
rect 13955 9333 13967 9367
rect 13909 9327 13967 9333
rect 18230 9324 18236 9376
rect 18288 9324 18294 9376
rect 19334 9324 19340 9376
rect 19392 9324 19398 9376
rect 20165 9367 20223 9373
rect 20165 9333 20177 9367
rect 20211 9364 20223 9367
rect 20346 9364 20352 9376
rect 20211 9336 20352 9364
rect 20211 9333 20223 9336
rect 20165 9327 20223 9333
rect 20346 9324 20352 9336
rect 20404 9324 20410 9376
rect 20714 9324 20720 9376
rect 20772 9324 20778 9376
rect 22094 9324 22100 9376
rect 22152 9364 22158 9376
rect 22296 9364 22324 9404
rect 27706 9392 27712 9404
rect 27764 9392 27770 9444
rect 32214 9432 32220 9444
rect 30208 9404 32220 9432
rect 22152 9336 22324 9364
rect 25041 9367 25099 9373
rect 22152 9324 22158 9336
rect 25041 9333 25053 9367
rect 25087 9364 25099 9367
rect 25314 9364 25320 9376
rect 25087 9336 25320 9364
rect 25087 9333 25099 9336
rect 25041 9327 25099 9333
rect 25314 9324 25320 9336
rect 25372 9324 25378 9376
rect 26513 9367 26571 9373
rect 26513 9333 26525 9367
rect 26559 9364 26571 9367
rect 27062 9364 27068 9376
rect 26559 9336 27068 9364
rect 26559 9333 26571 9336
rect 26513 9327 26571 9333
rect 27062 9324 27068 9336
rect 27120 9324 27126 9376
rect 27798 9324 27804 9376
rect 27856 9324 27862 9376
rect 27890 9324 27896 9376
rect 27948 9364 27954 9376
rect 30208 9364 30236 9404
rect 32214 9392 32220 9404
rect 32272 9392 32278 9444
rect 32306 9392 32312 9444
rect 32364 9432 32370 9444
rect 32401 9435 32459 9441
rect 32401 9432 32413 9435
rect 32364 9404 32413 9432
rect 32364 9392 32370 9404
rect 32401 9401 32413 9404
rect 32447 9401 32459 9435
rect 32401 9395 32459 9401
rect 34793 9435 34851 9441
rect 34793 9401 34805 9435
rect 34839 9432 34851 9435
rect 36464 9432 36492 9531
rect 36722 9528 36728 9580
rect 36780 9528 36786 9580
rect 36814 9528 36820 9580
rect 36872 9528 36878 9580
rect 37458 9528 37464 9580
rect 37516 9528 37522 9580
rect 36541 9503 36599 9509
rect 36541 9469 36553 9503
rect 36587 9500 36599 9503
rect 37550 9500 37556 9512
rect 36587 9472 37556 9500
rect 36587 9469 36599 9472
rect 36541 9463 36599 9469
rect 37550 9460 37556 9472
rect 37608 9460 37614 9512
rect 37642 9432 37648 9444
rect 34839 9404 37648 9432
rect 34839 9401 34851 9404
rect 34793 9395 34851 9401
rect 37642 9392 37648 9404
rect 37700 9392 37706 9444
rect 39393 9435 39451 9441
rect 39393 9401 39405 9435
rect 39439 9432 39451 9435
rect 39500 9432 39528 9608
rect 42886 9596 42892 9608
rect 42944 9596 42950 9648
rect 39577 9571 39635 9577
rect 39577 9537 39589 9571
rect 39623 9537 39635 9571
rect 39577 9531 39635 9537
rect 39669 9571 39727 9577
rect 39669 9537 39681 9571
rect 39715 9568 39727 9571
rect 39758 9568 39764 9580
rect 39715 9540 39764 9568
rect 39715 9537 39727 9540
rect 39669 9531 39727 9537
rect 39439 9404 39528 9432
rect 39592 9432 39620 9531
rect 39758 9528 39764 9540
rect 39816 9528 39822 9580
rect 39942 9528 39948 9580
rect 40000 9568 40006 9580
rect 40402 9568 40408 9580
rect 40000 9540 40408 9568
rect 40000 9528 40006 9540
rect 40402 9528 40408 9540
rect 40460 9568 40466 9580
rect 40460 9540 40540 9568
rect 40460 9528 40466 9540
rect 40126 9460 40132 9512
rect 40184 9460 40190 9512
rect 40512 9509 40540 9540
rect 41598 9528 41604 9580
rect 41656 9528 41662 9580
rect 41693 9571 41751 9577
rect 41693 9537 41705 9571
rect 41739 9568 41751 9571
rect 41739 9540 42564 9568
rect 41739 9537 41751 9540
rect 41693 9531 41751 9537
rect 40497 9503 40555 9509
rect 40497 9469 40509 9503
rect 40543 9469 40555 9503
rect 40497 9463 40555 9469
rect 40586 9460 40592 9512
rect 40644 9509 40650 9512
rect 40644 9503 40672 9509
rect 40660 9500 40672 9503
rect 41046 9500 41052 9512
rect 40660 9472 41052 9500
rect 40660 9469 40672 9472
rect 40644 9463 40672 9469
rect 40644 9460 40650 9463
rect 41046 9460 41052 9472
rect 41104 9460 41110 9512
rect 41877 9503 41935 9509
rect 41877 9469 41889 9503
rect 41923 9500 41935 9503
rect 41966 9500 41972 9512
rect 41923 9472 41972 9500
rect 41923 9469 41935 9472
rect 41877 9463 41935 9469
rect 41966 9460 41972 9472
rect 42024 9460 42030 9512
rect 39666 9432 39672 9444
rect 39592 9404 39672 9432
rect 39439 9401 39451 9404
rect 39393 9395 39451 9401
rect 39666 9392 39672 9404
rect 39724 9392 39730 9444
rect 40034 9392 40040 9444
rect 40092 9432 40098 9444
rect 41233 9435 41291 9441
rect 40092 9404 40908 9432
rect 40092 9392 40098 9404
rect 27948 9336 30236 9364
rect 27948 9324 27954 9336
rect 30558 9324 30564 9376
rect 30616 9364 30622 9376
rect 30653 9367 30711 9373
rect 30653 9364 30665 9367
rect 30616 9336 30665 9364
rect 30616 9324 30622 9336
rect 30653 9333 30665 9336
rect 30699 9333 30711 9367
rect 30653 9327 30711 9333
rect 30742 9324 30748 9376
rect 30800 9364 30806 9376
rect 31113 9367 31171 9373
rect 31113 9364 31125 9367
rect 30800 9336 31125 9364
rect 30800 9324 30806 9336
rect 31113 9333 31125 9336
rect 31159 9333 31171 9367
rect 31113 9327 31171 9333
rect 36909 9367 36967 9373
rect 36909 9333 36921 9367
rect 36955 9364 36967 9367
rect 36998 9364 37004 9376
rect 36955 9336 37004 9364
rect 36955 9333 36967 9336
rect 36909 9327 36967 9333
rect 36998 9324 37004 9336
rect 37056 9324 37062 9376
rect 37550 9324 37556 9376
rect 37608 9364 37614 9376
rect 40773 9367 40831 9373
rect 40773 9364 40785 9367
rect 37608 9336 40785 9364
rect 37608 9324 37614 9336
rect 40773 9333 40785 9336
rect 40819 9333 40831 9367
rect 40880 9364 40908 9404
rect 41233 9401 41245 9435
rect 41279 9432 41291 9435
rect 41782 9432 41788 9444
rect 41279 9404 41788 9432
rect 41279 9401 41291 9404
rect 41233 9395 41291 9401
rect 41782 9392 41788 9404
rect 41840 9392 41846 9444
rect 42536 9432 42564 9540
rect 42610 9528 42616 9580
rect 42668 9528 42674 9580
rect 42702 9528 42708 9580
rect 42760 9568 42766 9580
rect 42797 9571 42855 9577
rect 42797 9568 42809 9571
rect 42760 9540 42809 9568
rect 42760 9528 42766 9540
rect 42797 9537 42809 9540
rect 42843 9537 42855 9571
rect 42797 9531 42855 9537
rect 44174 9432 44180 9444
rect 42536 9404 44180 9432
rect 44174 9392 44180 9404
rect 44232 9392 44238 9444
rect 41322 9364 41328 9376
rect 40880 9336 41328 9364
rect 40773 9327 40831 9333
rect 41322 9324 41328 9336
rect 41380 9364 41386 9376
rect 42610 9364 42616 9376
rect 41380 9336 42616 9364
rect 41380 9324 41386 9336
rect 42610 9324 42616 9336
rect 42668 9324 42674 9376
rect 42705 9367 42763 9373
rect 42705 9333 42717 9367
rect 42751 9364 42763 9367
rect 42886 9364 42892 9376
rect 42751 9336 42892 9364
rect 42751 9333 42763 9336
rect 42705 9327 42763 9333
rect 42886 9324 42892 9336
rect 42944 9324 42950 9376
rect 1104 9274 44896 9296
rect 1104 9222 6423 9274
rect 6475 9222 6487 9274
rect 6539 9222 6551 9274
rect 6603 9222 6615 9274
rect 6667 9222 6679 9274
rect 6731 9222 17370 9274
rect 17422 9222 17434 9274
rect 17486 9222 17498 9274
rect 17550 9222 17562 9274
rect 17614 9222 17626 9274
rect 17678 9222 28317 9274
rect 28369 9222 28381 9274
rect 28433 9222 28445 9274
rect 28497 9222 28509 9274
rect 28561 9222 28573 9274
rect 28625 9222 39264 9274
rect 39316 9222 39328 9274
rect 39380 9222 39392 9274
rect 39444 9222 39456 9274
rect 39508 9222 39520 9274
rect 39572 9222 44896 9274
rect 1104 9200 44896 9222
rect 5810 9120 5816 9172
rect 5868 9160 5874 9172
rect 7098 9160 7104 9172
rect 5868 9132 7104 9160
rect 5868 9120 5874 9132
rect 7098 9120 7104 9132
rect 7156 9120 7162 9172
rect 10870 9120 10876 9172
rect 10928 9160 10934 9172
rect 12161 9163 12219 9169
rect 10928 9132 12112 9160
rect 10928 9120 10934 9132
rect 7558 9052 7564 9104
rect 7616 9052 7622 9104
rect 12084 9092 12112 9132
rect 12161 9129 12173 9163
rect 12207 9160 12219 9163
rect 12250 9160 12256 9172
rect 12207 9132 12256 9160
rect 12207 9129 12219 9132
rect 12161 9123 12219 9129
rect 12250 9120 12256 9132
rect 12308 9120 12314 9172
rect 12986 9160 12992 9172
rect 12406 9132 12992 9160
rect 12406 9092 12434 9132
rect 12986 9120 12992 9132
rect 13044 9120 13050 9172
rect 13078 9120 13084 9172
rect 13136 9160 13142 9172
rect 14277 9163 14335 9169
rect 14277 9160 14289 9163
rect 13136 9132 14289 9160
rect 13136 9120 13142 9132
rect 14277 9129 14289 9132
rect 14323 9129 14335 9163
rect 17218 9160 17224 9172
rect 14277 9123 14335 9129
rect 16224 9132 17224 9160
rect 12084 9064 12434 9092
rect 12621 9095 12679 9101
rect 12621 9061 12633 9095
rect 12667 9092 12679 9095
rect 14090 9092 14096 9104
rect 12667 9064 14096 9092
rect 12667 9061 12679 9064
rect 12621 9055 12679 9061
rect 14090 9052 14096 9064
rect 14148 9052 14154 9104
rect 10686 8984 10692 9036
rect 10744 9024 10750 9036
rect 13081 9027 13139 9033
rect 13081 9024 13093 9027
rect 10744 8996 12296 9024
rect 10744 8984 10750 8996
rect 4154 8916 4160 8968
rect 4212 8956 4218 8968
rect 5261 8959 5319 8965
rect 5261 8956 5273 8959
rect 4212 8928 5273 8956
rect 4212 8916 4218 8928
rect 5261 8925 5273 8928
rect 5307 8925 5319 8959
rect 5261 8919 5319 8925
rect 5626 8916 5632 8968
rect 5684 8956 5690 8968
rect 5684 8928 8064 8956
rect 5684 8916 5690 8928
rect 6270 8848 6276 8900
rect 6328 8888 6334 8900
rect 7837 8891 7895 8897
rect 7837 8888 7849 8891
rect 6328 8860 7849 8888
rect 6328 8848 6334 8860
rect 7837 8857 7849 8860
rect 7883 8857 7895 8891
rect 7837 8851 7895 8857
rect 8036 8832 8064 8928
rect 9950 8916 9956 8968
rect 10008 8916 10014 8968
rect 10413 8959 10471 8965
rect 10413 8925 10425 8959
rect 10459 8925 10471 8959
rect 10413 8919 10471 8925
rect 8113 8891 8171 8897
rect 8113 8857 8125 8891
rect 8159 8888 8171 8891
rect 10226 8888 10232 8900
rect 8159 8860 10232 8888
rect 8159 8857 8171 8860
rect 8113 8851 8171 8857
rect 10226 8848 10232 8860
rect 10284 8848 10290 8900
rect 10428 8888 10456 8919
rect 10594 8888 10600 8900
rect 10428 8860 10600 8888
rect 10594 8848 10600 8860
rect 10652 8848 10658 8900
rect 10689 8891 10747 8897
rect 10689 8857 10701 8891
rect 10735 8888 10747 8891
rect 10962 8888 10968 8900
rect 10735 8860 10968 8888
rect 10735 8857 10747 8860
rect 10689 8851 10747 8857
rect 10962 8848 10968 8860
rect 11020 8848 11026 8900
rect 11072 8860 11178 8888
rect 5534 8780 5540 8832
rect 5592 8820 5598 8832
rect 6549 8823 6607 8829
rect 6549 8820 6561 8823
rect 5592 8792 6561 8820
rect 5592 8780 5598 8792
rect 6549 8789 6561 8792
rect 6595 8789 6607 8823
rect 6549 8783 6607 8789
rect 8018 8780 8024 8832
rect 8076 8780 8082 8832
rect 9766 8780 9772 8832
rect 9824 8780 9830 8832
rect 10318 8780 10324 8832
rect 10376 8820 10382 8832
rect 11072 8820 11100 8860
rect 10376 8792 11100 8820
rect 12268 8820 12296 8996
rect 12912 8996 13093 9024
rect 12912 8888 12940 8996
rect 13081 8993 13093 8996
rect 13127 8993 13139 9027
rect 13081 8987 13139 8993
rect 13265 9027 13323 9033
rect 13265 8993 13277 9027
rect 13311 9024 13323 9027
rect 13538 9024 13544 9036
rect 13311 8996 13544 9024
rect 13311 8993 13323 8996
rect 13265 8987 13323 8993
rect 13538 8984 13544 8996
rect 13596 8984 13602 9036
rect 16224 9024 16252 9132
rect 17218 9120 17224 9132
rect 17276 9120 17282 9172
rect 17589 9163 17647 9169
rect 17589 9129 17601 9163
rect 17635 9160 17647 9163
rect 18506 9160 18512 9172
rect 17635 9132 18512 9160
rect 17635 9129 17647 9132
rect 17589 9123 17647 9129
rect 18506 9120 18512 9132
rect 18564 9120 18570 9172
rect 23474 9120 23480 9172
rect 23532 9160 23538 9172
rect 23750 9160 23756 9172
rect 23532 9132 23756 9160
rect 23532 9120 23538 9132
rect 23750 9120 23756 9132
rect 23808 9160 23814 9172
rect 23808 9132 25912 9160
rect 23808 9120 23814 9132
rect 19334 9052 19340 9104
rect 19392 9092 19398 9104
rect 19392 9064 20944 9092
rect 19392 9052 19398 9064
rect 14844 8996 16252 9024
rect 12989 8959 13047 8965
rect 12989 8925 13001 8959
rect 13035 8956 13047 8959
rect 13446 8956 13452 8968
rect 13035 8928 13452 8956
rect 13035 8925 13047 8928
rect 12989 8919 13047 8925
rect 13446 8916 13452 8928
rect 13504 8916 13510 8968
rect 14458 8916 14464 8968
rect 14516 8916 14522 8968
rect 14844 8888 14872 8996
rect 19886 8984 19892 9036
rect 19944 9024 19950 9036
rect 20809 9027 20867 9033
rect 20809 9024 20821 9027
rect 19944 8996 20821 9024
rect 19944 8984 19950 8996
rect 20809 8993 20821 8996
rect 20855 8993 20867 9027
rect 20916 9024 20944 9064
rect 22554 9052 22560 9104
rect 22612 9092 22618 9104
rect 23293 9095 23351 9101
rect 23293 9092 23305 9095
rect 22612 9064 23305 9092
rect 22612 9052 22618 9064
rect 23293 9061 23305 9064
rect 23339 9061 23351 9095
rect 25884 9092 25912 9132
rect 26326 9120 26332 9172
rect 26384 9120 26390 9172
rect 28074 9160 28080 9172
rect 26436 9132 28080 9160
rect 26436 9092 26464 9132
rect 28074 9120 28080 9132
rect 28132 9120 28138 9172
rect 29178 9120 29184 9172
rect 29236 9120 29242 9172
rect 35158 9120 35164 9172
rect 35216 9120 35222 9172
rect 40037 9163 40095 9169
rect 40037 9129 40049 9163
rect 40083 9160 40095 9163
rect 40218 9160 40224 9172
rect 40083 9132 40224 9160
rect 40083 9129 40095 9132
rect 40037 9123 40095 9129
rect 40218 9120 40224 9132
rect 40276 9120 40282 9172
rect 41598 9160 41604 9172
rect 40328 9132 41604 9160
rect 25884 9064 26464 9092
rect 23293 9055 23351 9061
rect 31386 9052 31392 9104
rect 31444 9092 31450 9104
rect 32033 9095 32091 9101
rect 31444 9064 31616 9092
rect 31444 9052 31450 9064
rect 21085 9027 21143 9033
rect 21085 9024 21097 9027
rect 20916 8996 21097 9024
rect 20809 8987 20867 8993
rect 21085 8993 21097 8996
rect 21131 8993 21143 9027
rect 21085 8987 21143 8993
rect 23017 9027 23075 9033
rect 23017 8993 23029 9027
rect 23063 9024 23075 9027
rect 23658 9024 23664 9036
rect 23063 8996 23664 9024
rect 23063 8993 23075 8996
rect 23017 8987 23075 8993
rect 23658 8984 23664 8996
rect 23716 9024 23722 9036
rect 31588 9033 31616 9064
rect 32033 9061 32045 9095
rect 32079 9092 32091 9095
rect 35802 9092 35808 9104
rect 32079 9064 35808 9092
rect 32079 9061 32091 9064
rect 32033 9055 32091 9061
rect 30745 9027 30803 9033
rect 30745 9024 30757 9027
rect 23716 8996 27936 9024
rect 23716 8984 23722 8996
rect 14918 8916 14924 8968
rect 14976 8956 14982 8968
rect 16209 8959 16267 8965
rect 16209 8956 16221 8959
rect 14976 8928 16221 8956
rect 14976 8916 14982 8928
rect 16209 8925 16221 8928
rect 16255 8956 16267 8959
rect 16850 8956 16856 8968
rect 16255 8928 16856 8956
rect 16255 8925 16267 8928
rect 16209 8919 16267 8925
rect 16850 8916 16856 8928
rect 16908 8916 16914 8968
rect 18230 8916 18236 8968
rect 18288 8916 18294 8968
rect 19705 8959 19763 8965
rect 19705 8925 19717 8959
rect 19751 8956 19763 8959
rect 20162 8956 20168 8968
rect 19751 8928 20168 8956
rect 19751 8925 19763 8928
rect 19705 8919 19763 8925
rect 20162 8916 20168 8928
rect 20220 8916 20226 8968
rect 20346 8916 20352 8968
rect 20404 8916 20410 8968
rect 24486 8916 24492 8968
rect 24544 8956 24550 8968
rect 24581 8959 24639 8965
rect 24581 8956 24593 8959
rect 24544 8928 24593 8956
rect 24544 8916 24550 8928
rect 24581 8925 24593 8928
rect 24627 8925 24639 8959
rect 26973 8959 27031 8965
rect 26973 8956 26985 8959
rect 24581 8919 24639 8925
rect 26160 8928 26985 8956
rect 12912 8860 14872 8888
rect 15562 8848 15568 8900
rect 15620 8888 15626 8900
rect 16454 8891 16512 8897
rect 16454 8888 16466 8891
rect 15620 8860 16466 8888
rect 15620 8848 15626 8860
rect 16454 8857 16466 8860
rect 16500 8857 16512 8891
rect 20806 8888 20812 8900
rect 16454 8851 16512 8857
rect 17236 8860 20812 8888
rect 17236 8820 17264 8860
rect 20806 8848 20812 8860
rect 20864 8848 20870 8900
rect 21192 8860 21574 8888
rect 12268 8792 17264 8820
rect 10376 8780 10382 8792
rect 18046 8780 18052 8832
rect 18104 8780 18110 8832
rect 19518 8780 19524 8832
rect 19576 8780 19582 8832
rect 20165 8823 20223 8829
rect 20165 8789 20177 8823
rect 20211 8820 20223 8823
rect 21192 8820 21220 8860
rect 24854 8848 24860 8900
rect 24912 8848 24918 8900
rect 25314 8848 25320 8900
rect 25372 8848 25378 8900
rect 20211 8792 21220 8820
rect 22557 8823 22615 8829
rect 20211 8789 20223 8792
rect 20165 8783 20223 8789
rect 22557 8789 22569 8823
rect 22603 8820 22615 8823
rect 23198 8820 23204 8832
rect 22603 8792 23204 8820
rect 22603 8789 22615 8792
rect 22557 8783 22615 8789
rect 23198 8780 23204 8792
rect 23256 8780 23262 8832
rect 23474 8780 23480 8832
rect 23532 8780 23538 8832
rect 25130 8780 25136 8832
rect 25188 8820 25194 8832
rect 26160 8820 26188 8928
rect 26973 8925 26985 8928
rect 27019 8925 27031 8959
rect 26973 8919 27031 8925
rect 26988 8888 27016 8919
rect 27062 8916 27068 8968
rect 27120 8956 27126 8968
rect 27249 8959 27307 8965
rect 27249 8956 27261 8959
rect 27120 8928 27261 8956
rect 27120 8916 27126 8928
rect 27249 8925 27261 8928
rect 27295 8925 27307 8959
rect 27249 8919 27307 8925
rect 27522 8916 27528 8968
rect 27580 8956 27586 8968
rect 27801 8959 27859 8965
rect 27801 8956 27813 8959
rect 27580 8928 27813 8956
rect 27580 8916 27586 8928
rect 27801 8925 27813 8928
rect 27847 8925 27859 8959
rect 27908 8956 27936 8996
rect 29840 8996 30757 9024
rect 29840 8956 29868 8996
rect 30745 8993 30757 8996
rect 30791 8993 30803 9027
rect 30745 8987 30803 8993
rect 31573 9027 31631 9033
rect 31573 8993 31585 9027
rect 31619 8993 31631 9027
rect 31573 8987 31631 8993
rect 32214 8984 32220 9036
rect 32272 9024 32278 9036
rect 33873 9027 33931 9033
rect 33873 9024 33885 9027
rect 32272 8996 33885 9024
rect 32272 8984 32278 8996
rect 33873 8993 33885 8996
rect 33919 8993 33931 9027
rect 33873 8987 33931 8993
rect 35250 8984 35256 9036
rect 35308 9024 35314 9036
rect 35452 9033 35480 9064
rect 35802 9052 35808 9064
rect 35860 9052 35866 9104
rect 39209 9095 39267 9101
rect 39209 9061 39221 9095
rect 39255 9092 39267 9095
rect 39850 9092 39856 9104
rect 39255 9064 39856 9092
rect 39255 9061 39267 9064
rect 39209 9055 39267 9061
rect 39850 9052 39856 9064
rect 39908 9052 39914 9104
rect 40328 9092 40356 9132
rect 41598 9120 41604 9132
rect 41656 9120 41662 9172
rect 40144 9064 40356 9092
rect 35345 9027 35403 9033
rect 35345 9024 35357 9027
rect 35308 8996 35357 9024
rect 35308 8984 35314 8996
rect 35345 8993 35357 8996
rect 35391 8993 35403 9027
rect 35345 8987 35403 8993
rect 35437 9027 35495 9033
rect 35437 8993 35449 9027
rect 35483 8993 35495 9027
rect 37274 9024 37280 9036
rect 35437 8987 35495 8993
rect 35544 8996 37280 9024
rect 27908 8928 29868 8956
rect 27801 8919 27859 8925
rect 30558 8916 30564 8968
rect 30616 8916 30622 8968
rect 31478 8916 31484 8968
rect 31536 8956 31542 8968
rect 31665 8959 31723 8965
rect 31665 8956 31677 8959
rect 31536 8928 31677 8956
rect 31536 8916 31542 8928
rect 31665 8925 31677 8928
rect 31711 8925 31723 8959
rect 31665 8919 31723 8925
rect 33965 8959 34023 8965
rect 33965 8925 33977 8959
rect 34011 8956 34023 8959
rect 34146 8956 34152 8968
rect 34011 8928 34152 8956
rect 34011 8925 34023 8928
rect 33965 8919 34023 8925
rect 34146 8916 34152 8928
rect 34204 8916 34210 8968
rect 35544 8956 35572 8996
rect 37274 8984 37280 8996
rect 37332 8984 37338 9036
rect 37366 8984 37372 9036
rect 37424 9024 37430 9036
rect 40144 9024 40172 9064
rect 37424 8996 40172 9024
rect 37424 8984 37430 8996
rect 34256 8952 35388 8956
rect 35452 8952 35572 8956
rect 34256 8928 35572 8952
rect 28074 8897 28080 8900
rect 26988 8860 28028 8888
rect 25188 8792 26188 8820
rect 25188 8780 25194 8792
rect 26234 8780 26240 8832
rect 26292 8820 26298 8832
rect 26789 8823 26847 8829
rect 26789 8820 26801 8823
rect 26292 8792 26801 8820
rect 26292 8780 26298 8792
rect 26789 8789 26801 8792
rect 26835 8789 26847 8823
rect 26789 8783 26847 8789
rect 27157 8823 27215 8829
rect 27157 8789 27169 8823
rect 27203 8820 27215 8823
rect 27890 8820 27896 8832
rect 27203 8792 27896 8820
rect 27203 8789 27215 8792
rect 27157 8783 27215 8789
rect 27890 8780 27896 8792
rect 27948 8780 27954 8832
rect 28000 8820 28028 8860
rect 28068 8851 28080 8897
rect 28132 8888 28138 8900
rect 30098 8888 30104 8900
rect 28132 8860 30104 8888
rect 28074 8848 28080 8851
rect 28132 8848 28138 8860
rect 30098 8848 30104 8860
rect 30156 8848 30162 8900
rect 34256 8888 34284 8928
rect 35360 8924 35480 8928
rect 35618 8916 35624 8968
rect 35676 8956 35682 8968
rect 35805 8959 35863 8965
rect 35805 8956 35817 8959
rect 35676 8928 35817 8956
rect 35676 8916 35682 8928
rect 35805 8925 35817 8928
rect 35851 8956 35863 8959
rect 36265 8959 36323 8965
rect 35851 8928 35940 8956
rect 35851 8925 35863 8928
rect 35805 8919 35863 8925
rect 30208 8860 34284 8888
rect 29086 8820 29092 8832
rect 28000 8792 29092 8820
rect 29086 8780 29092 8792
rect 29144 8780 29150 8832
rect 30208 8829 30236 8860
rect 35066 8848 35072 8900
rect 35124 8888 35130 8900
rect 35912 8888 35940 8928
rect 36265 8925 36277 8959
rect 36311 8956 36323 8959
rect 36998 8956 37004 8968
rect 36311 8928 37004 8956
rect 36311 8925 36323 8928
rect 36265 8919 36323 8925
rect 36998 8916 37004 8928
rect 37056 8916 37062 8968
rect 38749 8959 38807 8965
rect 38749 8925 38761 8959
rect 38795 8956 38807 8959
rect 39390 8956 39396 8968
rect 38795 8928 39396 8956
rect 38795 8925 38807 8928
rect 38749 8919 38807 8925
rect 39390 8916 39396 8928
rect 39448 8916 39454 8968
rect 39485 8959 39543 8965
rect 39485 8925 39497 8959
rect 39531 8956 39543 8959
rect 39758 8956 39764 8968
rect 39531 8928 39764 8956
rect 39531 8925 39543 8928
rect 39485 8919 39543 8925
rect 39758 8916 39764 8928
rect 39816 8916 39822 8968
rect 40034 8916 40040 8968
rect 40092 8916 40098 8968
rect 40221 8959 40279 8965
rect 40221 8925 40233 8959
rect 40267 8956 40279 8959
rect 40310 8956 40316 8968
rect 40267 8928 40316 8956
rect 40267 8925 40279 8928
rect 40221 8919 40279 8925
rect 40310 8916 40316 8928
rect 40368 8916 40374 8968
rect 40494 8916 40500 8968
rect 40552 8956 40558 8968
rect 40681 8959 40739 8965
rect 40681 8956 40693 8959
rect 40552 8928 40693 8956
rect 40552 8916 40558 8928
rect 40681 8925 40693 8928
rect 40727 8956 40739 8959
rect 42521 8959 42579 8965
rect 42521 8956 42533 8959
rect 40727 8928 42533 8956
rect 40727 8925 40739 8928
rect 40681 8919 40739 8925
rect 42521 8925 42533 8928
rect 42567 8925 42579 8959
rect 42521 8919 42579 8925
rect 38930 8888 38936 8900
rect 35124 8860 35848 8888
rect 35912 8860 38936 8888
rect 35124 8848 35130 8860
rect 30193 8823 30251 8829
rect 30193 8789 30205 8823
rect 30239 8789 30251 8823
rect 30193 8783 30251 8789
rect 30653 8823 30711 8829
rect 30653 8789 30665 8823
rect 30699 8820 30711 8823
rect 31202 8820 31208 8832
rect 30699 8792 31208 8820
rect 30699 8789 30711 8792
rect 30653 8783 30711 8789
rect 31202 8780 31208 8792
rect 31260 8780 31266 8832
rect 34333 8823 34391 8829
rect 34333 8789 34345 8823
rect 34379 8820 34391 8823
rect 35529 8823 35587 8829
rect 35529 8820 35541 8823
rect 34379 8792 35541 8820
rect 34379 8789 34391 8792
rect 34333 8783 34391 8789
rect 35529 8789 35541 8792
rect 35575 8820 35587 8823
rect 35618 8820 35624 8832
rect 35575 8792 35624 8820
rect 35575 8789 35587 8792
rect 35529 8783 35587 8789
rect 35618 8780 35624 8792
rect 35676 8780 35682 8832
rect 35710 8780 35716 8832
rect 35768 8780 35774 8832
rect 35820 8820 35848 8860
rect 38930 8848 38936 8860
rect 38988 8848 38994 8900
rect 39206 8848 39212 8900
rect 39264 8848 39270 8900
rect 42794 8897 42800 8900
rect 40926 8891 40984 8897
rect 40926 8888 40938 8891
rect 39316 8860 40938 8888
rect 36449 8823 36507 8829
rect 36449 8820 36461 8823
rect 35820 8792 36461 8820
rect 36449 8789 36461 8792
rect 36495 8820 36507 8823
rect 38470 8820 38476 8832
rect 36495 8792 38476 8820
rect 36495 8789 36507 8792
rect 36449 8783 36507 8789
rect 38470 8780 38476 8792
rect 38528 8780 38534 8832
rect 38565 8823 38623 8829
rect 38565 8789 38577 8823
rect 38611 8820 38623 8823
rect 39316 8820 39344 8860
rect 40926 8857 40938 8860
rect 40972 8857 40984 8891
rect 40926 8851 40984 8857
rect 42788 8851 42800 8897
rect 42794 8848 42800 8851
rect 42852 8848 42858 8900
rect 38611 8792 39344 8820
rect 39393 8823 39451 8829
rect 38611 8789 38623 8792
rect 38565 8783 38623 8789
rect 39393 8789 39405 8823
rect 39439 8820 39451 8823
rect 39666 8820 39672 8832
rect 39439 8792 39672 8820
rect 39439 8789 39451 8792
rect 39393 8783 39451 8789
rect 39666 8780 39672 8792
rect 39724 8820 39730 8832
rect 41046 8820 41052 8832
rect 39724 8792 41052 8820
rect 39724 8780 39730 8792
rect 41046 8780 41052 8792
rect 41104 8820 41110 8832
rect 42061 8823 42119 8829
rect 42061 8820 42073 8823
rect 41104 8792 42073 8820
rect 41104 8780 41110 8792
rect 42061 8789 42073 8792
rect 42107 8789 42119 8823
rect 42061 8783 42119 8789
rect 42702 8780 42708 8832
rect 42760 8820 42766 8832
rect 43901 8823 43959 8829
rect 43901 8820 43913 8823
rect 42760 8792 43913 8820
rect 42760 8780 42766 8792
rect 43901 8789 43913 8792
rect 43947 8789 43959 8823
rect 43901 8783 43959 8789
rect 1104 8730 45051 8752
rect 1104 8678 11896 8730
rect 11948 8678 11960 8730
rect 12012 8678 12024 8730
rect 12076 8678 12088 8730
rect 12140 8678 12152 8730
rect 12204 8678 22843 8730
rect 22895 8678 22907 8730
rect 22959 8678 22971 8730
rect 23023 8678 23035 8730
rect 23087 8678 23099 8730
rect 23151 8678 33790 8730
rect 33842 8678 33854 8730
rect 33906 8678 33918 8730
rect 33970 8678 33982 8730
rect 34034 8678 34046 8730
rect 34098 8678 44737 8730
rect 44789 8678 44801 8730
rect 44853 8678 44865 8730
rect 44917 8678 44929 8730
rect 44981 8678 44993 8730
rect 45045 8678 45051 8730
rect 1104 8656 45051 8678
rect 2774 8616 2780 8628
rect 2148 8588 2780 8616
rect 2148 8489 2176 8588
rect 2774 8576 2780 8588
rect 2832 8616 2838 8628
rect 3786 8616 3792 8628
rect 2832 8588 3792 8616
rect 2832 8576 2838 8588
rect 3786 8576 3792 8588
rect 3844 8576 3850 8628
rect 7650 8616 7656 8628
rect 3896 8588 4660 8616
rect 2133 8483 2191 8489
rect 2133 8449 2145 8483
rect 2179 8449 2191 8483
rect 2133 8443 2191 8449
rect 2400 8483 2458 8489
rect 2400 8449 2412 8483
rect 2446 8480 2458 8483
rect 3896 8480 3924 8588
rect 4240 8551 4298 8557
rect 4240 8517 4252 8551
rect 4286 8548 4298 8551
rect 4430 8548 4436 8560
rect 4286 8520 4436 8548
rect 4286 8517 4298 8520
rect 4240 8511 4298 8517
rect 2446 8452 3924 8480
rect 2446 8449 2458 8452
rect 2400 8443 2458 8449
rect 3970 8440 3976 8492
rect 4028 8440 4034 8492
rect 4255 8480 4283 8511
rect 4430 8508 4436 8520
rect 4488 8508 4494 8560
rect 4080 8452 4283 8480
rect 4632 8480 4660 8588
rect 6932 8588 7656 8616
rect 6816 8551 6874 8557
rect 6816 8517 6828 8551
rect 6862 8548 6874 8551
rect 6932 8548 6960 8588
rect 7650 8576 7656 8588
rect 7708 8576 7714 8628
rect 8018 8576 8024 8628
rect 8076 8616 8082 8628
rect 9769 8619 9827 8625
rect 9769 8616 9781 8619
rect 8076 8588 9781 8616
rect 8076 8576 8082 8588
rect 9769 8585 9781 8588
rect 9815 8585 9827 8619
rect 9769 8579 9827 8585
rect 10318 8576 10324 8628
rect 10376 8576 10382 8628
rect 10962 8576 10968 8628
rect 11020 8576 11026 8628
rect 11606 8576 11612 8628
rect 11664 8616 11670 8628
rect 11664 8588 12112 8616
rect 11664 8576 11670 8588
rect 6862 8520 6960 8548
rect 6862 8517 6874 8520
rect 6816 8511 6874 8517
rect 7006 8508 7012 8560
rect 7064 8548 7070 8560
rect 8634 8551 8692 8557
rect 8634 8548 8646 8551
rect 7064 8520 8646 8548
rect 7064 8508 7070 8520
rect 8634 8517 8646 8520
rect 8680 8517 8692 8551
rect 8634 8511 8692 8517
rect 10226 8508 10232 8560
rect 10284 8548 10290 8560
rect 11514 8548 11520 8560
rect 10284 8520 11520 8548
rect 10284 8508 10290 8520
rect 11514 8508 11520 8520
rect 11572 8508 11578 8560
rect 11882 8508 11888 8560
rect 11940 8548 11946 8560
rect 11977 8551 12035 8557
rect 11977 8548 11989 8551
rect 11940 8520 11989 8548
rect 11940 8508 11946 8520
rect 11977 8517 11989 8520
rect 12023 8517 12035 8551
rect 12084 8548 12112 8588
rect 12894 8576 12900 8628
rect 12952 8616 12958 8628
rect 13449 8619 13507 8625
rect 13449 8616 13461 8619
rect 12952 8588 13461 8616
rect 12952 8576 12958 8588
rect 13449 8585 13461 8588
rect 13495 8585 13507 8619
rect 13449 8579 13507 8585
rect 14936 8588 19932 8616
rect 12084 8520 12466 8548
rect 11977 8511 12035 8517
rect 4632 8452 7972 8480
rect 4080 8412 4108 8452
rect 3528 8384 4108 8412
rect 3528 8353 3556 8384
rect 6270 8372 6276 8424
rect 6328 8412 6334 8424
rect 6549 8415 6607 8421
rect 6549 8412 6561 8415
rect 6328 8384 6561 8412
rect 6328 8372 6334 8384
rect 6549 8381 6561 8384
rect 6595 8381 6607 8415
rect 6549 8375 6607 8381
rect 7944 8356 7972 8452
rect 8202 8440 8208 8492
rect 8260 8480 8266 8492
rect 8260 8452 9444 8480
rect 8260 8440 8266 8452
rect 8389 8415 8447 8421
rect 8389 8381 8401 8415
rect 8435 8381 8447 8415
rect 8389 8375 8447 8381
rect 3513 8347 3571 8353
rect 3513 8313 3525 8347
rect 3559 8313 3571 8347
rect 3513 8307 3571 8313
rect 7926 8304 7932 8356
rect 7984 8304 7990 8356
rect 8404 8344 8432 8375
rect 8312 8316 8432 8344
rect 9416 8344 9444 8452
rect 10502 8440 10508 8492
rect 10560 8440 10566 8492
rect 11146 8440 11152 8492
rect 11204 8440 11210 8492
rect 11701 8483 11759 8489
rect 11701 8480 11713 8483
rect 11256 8452 11713 8480
rect 10594 8372 10600 8424
rect 10652 8412 10658 8424
rect 11256 8412 11284 8452
rect 11701 8449 11713 8452
rect 11747 8449 11759 8483
rect 11701 8443 11759 8449
rect 14936 8412 14964 8588
rect 15565 8551 15623 8557
rect 15565 8517 15577 8551
rect 15611 8548 15623 8551
rect 15654 8548 15660 8560
rect 15611 8520 15660 8548
rect 15611 8517 15623 8520
rect 15565 8511 15623 8517
rect 15654 8508 15660 8520
rect 15712 8508 15718 8560
rect 16850 8508 16856 8560
rect 16908 8548 16914 8560
rect 19904 8548 19932 8588
rect 20162 8576 20168 8628
rect 20220 8616 20226 8628
rect 20625 8619 20683 8625
rect 20625 8616 20637 8619
rect 20220 8588 20637 8616
rect 20220 8576 20226 8588
rect 20625 8585 20637 8588
rect 20671 8585 20683 8619
rect 20625 8579 20683 8585
rect 21085 8619 21143 8625
rect 21085 8585 21097 8619
rect 21131 8616 21143 8619
rect 21174 8616 21180 8628
rect 21131 8588 21180 8616
rect 21131 8585 21143 8588
rect 21085 8579 21143 8585
rect 21174 8576 21180 8588
rect 21232 8576 21238 8628
rect 25130 8616 25136 8628
rect 21284 8588 25136 8616
rect 21284 8548 21312 8588
rect 25130 8576 25136 8588
rect 25188 8576 25194 8628
rect 25222 8576 25228 8628
rect 25280 8616 25286 8628
rect 25409 8619 25467 8625
rect 25409 8616 25421 8619
rect 25280 8588 25421 8616
rect 25280 8576 25286 8588
rect 25409 8585 25421 8588
rect 25455 8585 25467 8619
rect 25409 8579 25467 8585
rect 31294 8576 31300 8628
rect 31352 8576 31358 8628
rect 34977 8619 35035 8625
rect 34977 8585 34989 8619
rect 35023 8585 35035 8619
rect 34977 8579 35035 8585
rect 26050 8548 26056 8560
rect 16908 8520 18184 8548
rect 19904 8520 21312 8548
rect 22066 8520 23612 8548
rect 16908 8508 16914 8520
rect 15473 8483 15531 8489
rect 15473 8449 15485 8483
rect 15519 8480 15531 8483
rect 16206 8480 16212 8492
rect 15519 8452 16212 8480
rect 15519 8449 15531 8452
rect 15473 8443 15531 8449
rect 16206 8440 16212 8452
rect 16264 8440 16270 8492
rect 17236 8489 17264 8520
rect 17221 8483 17279 8489
rect 17221 8449 17233 8483
rect 17267 8449 17279 8483
rect 17221 8443 17279 8449
rect 17488 8483 17546 8489
rect 17488 8449 17500 8483
rect 17534 8480 17546 8483
rect 18046 8480 18052 8492
rect 17534 8452 18052 8480
rect 17534 8449 17546 8452
rect 17488 8443 17546 8449
rect 18046 8440 18052 8452
rect 18104 8440 18110 8492
rect 18156 8480 18184 8520
rect 19702 8480 19708 8492
rect 18156 8452 19708 8480
rect 19702 8440 19708 8452
rect 19760 8440 19766 8492
rect 19797 8483 19855 8489
rect 19797 8449 19809 8483
rect 19843 8480 19855 8483
rect 20898 8480 20904 8492
rect 19843 8452 20904 8480
rect 19843 8449 19855 8452
rect 19797 8443 19855 8449
rect 20898 8440 20904 8452
rect 20956 8440 20962 8492
rect 20993 8483 21051 8489
rect 20993 8449 21005 8483
rect 21039 8480 21051 8483
rect 21266 8480 21272 8492
rect 21039 8452 21272 8480
rect 21039 8449 21051 8452
rect 20993 8443 21051 8449
rect 21266 8440 21272 8452
rect 21324 8440 21330 8492
rect 15378 8412 15384 8424
rect 10652 8384 11284 8412
rect 11808 8384 14964 8412
rect 15028 8384 15384 8412
rect 10652 8372 10658 8384
rect 11808 8344 11836 8384
rect 15028 8344 15056 8384
rect 15378 8372 15384 8384
rect 15436 8372 15442 8424
rect 15654 8372 15660 8424
rect 15712 8372 15718 8424
rect 19889 8415 19947 8421
rect 19889 8381 19901 8415
rect 19935 8412 19947 8415
rect 19978 8412 19984 8424
rect 19935 8384 19984 8412
rect 19935 8381 19947 8384
rect 19889 8375 19947 8381
rect 19978 8372 19984 8384
rect 20036 8372 20042 8424
rect 20070 8372 20076 8424
rect 20128 8412 20134 8424
rect 21177 8415 21235 8421
rect 21177 8412 21189 8415
rect 20128 8384 21189 8412
rect 20128 8372 20134 8384
rect 21177 8381 21189 8384
rect 21223 8412 21235 8415
rect 22066 8412 22094 8520
rect 22462 8489 22468 8492
rect 22456 8443 22468 8489
rect 22462 8440 22468 8443
rect 22520 8440 22526 8492
rect 21223 8384 22094 8412
rect 21223 8381 21235 8384
rect 21177 8375 21235 8381
rect 22186 8372 22192 8424
rect 22244 8372 22250 8424
rect 9416 8316 11836 8344
rect 13004 8316 15056 8344
rect 15105 8347 15163 8353
rect 5350 8236 5356 8288
rect 5408 8236 5414 8288
rect 7742 8236 7748 8288
rect 7800 8276 7806 8288
rect 8312 8276 8340 8316
rect 7800 8248 8340 8276
rect 7800 8236 7806 8248
rect 11514 8236 11520 8288
rect 11572 8276 11578 8288
rect 13004 8276 13032 8316
rect 15105 8313 15117 8347
rect 15151 8344 15163 8347
rect 16850 8344 16856 8356
rect 15151 8316 16856 8344
rect 15151 8313 15163 8316
rect 15105 8307 15163 8313
rect 16850 8304 16856 8316
rect 16908 8304 16914 8356
rect 19429 8347 19487 8353
rect 19429 8313 19441 8347
rect 19475 8344 19487 8347
rect 21910 8344 21916 8356
rect 19475 8316 21916 8344
rect 19475 8313 19487 8316
rect 19429 8307 19487 8313
rect 21910 8304 21916 8316
rect 21968 8304 21974 8356
rect 23584 8353 23612 8520
rect 25424 8520 26056 8548
rect 25424 8489 25452 8520
rect 26050 8508 26056 8520
rect 26108 8548 26114 8560
rect 26421 8551 26479 8557
rect 26421 8548 26433 8551
rect 26108 8520 26433 8548
rect 26108 8508 26114 8520
rect 26421 8517 26433 8520
rect 26467 8548 26479 8551
rect 27430 8548 27436 8560
rect 26467 8520 27436 8548
rect 26467 8517 26479 8520
rect 26421 8511 26479 8517
rect 27430 8508 27436 8520
rect 27488 8508 27494 8560
rect 28077 8551 28135 8557
rect 28077 8517 28089 8551
rect 28123 8548 28135 8551
rect 28166 8548 28172 8560
rect 28123 8520 28172 8548
rect 28123 8517 28135 8520
rect 28077 8511 28135 8517
rect 28166 8508 28172 8520
rect 28224 8508 28230 8560
rect 31113 8551 31171 8557
rect 31113 8517 31125 8551
rect 31159 8548 31171 8551
rect 31846 8548 31852 8560
rect 31159 8520 31852 8548
rect 31159 8517 31171 8520
rect 31113 8511 31171 8517
rect 31846 8508 31852 8520
rect 31904 8508 31910 8560
rect 34992 8548 35020 8579
rect 35618 8576 35624 8628
rect 35676 8576 35682 8628
rect 35805 8619 35863 8625
rect 35805 8585 35817 8619
rect 35851 8616 35863 8619
rect 37458 8616 37464 8628
rect 35851 8588 37464 8616
rect 35851 8585 35863 8588
rect 35805 8579 35863 8585
rect 37458 8576 37464 8588
rect 37516 8576 37522 8628
rect 39390 8576 39396 8628
rect 39448 8576 39454 8628
rect 40678 8616 40684 8628
rect 39868 8588 40684 8616
rect 35529 8551 35587 8557
rect 35529 8548 35541 8551
rect 34992 8520 35541 8548
rect 35529 8517 35541 8520
rect 35575 8548 35587 8551
rect 35710 8548 35716 8560
rect 35575 8520 35716 8548
rect 35575 8517 35587 8520
rect 35529 8511 35587 8517
rect 35710 8508 35716 8520
rect 35768 8508 35774 8560
rect 36078 8508 36084 8560
rect 36136 8548 36142 8560
rect 36265 8551 36323 8557
rect 36265 8548 36277 8551
rect 36136 8520 36277 8548
rect 36136 8508 36142 8520
rect 36265 8517 36277 8520
rect 36311 8517 36323 8551
rect 36265 8511 36323 8517
rect 36481 8551 36539 8557
rect 36481 8517 36493 8551
rect 36527 8548 36539 8551
rect 37366 8548 37372 8560
rect 36527 8520 37372 8548
rect 36527 8517 36539 8520
rect 36481 8511 36539 8517
rect 37366 8508 37372 8520
rect 37424 8508 37430 8560
rect 38746 8508 38752 8560
rect 38804 8548 38810 8560
rect 39868 8548 39896 8588
rect 40678 8576 40684 8588
rect 40736 8616 40742 8628
rect 41690 8616 41696 8628
rect 40736 8588 41696 8616
rect 40736 8576 40742 8588
rect 41690 8576 41696 8588
rect 41748 8576 41754 8628
rect 42702 8616 42708 8628
rect 41800 8588 42708 8616
rect 38804 8520 39896 8548
rect 38804 8508 38810 8520
rect 25409 8483 25467 8489
rect 25409 8449 25421 8483
rect 25455 8449 25467 8483
rect 25409 8443 25467 8449
rect 25958 8440 25964 8492
rect 26016 8480 26022 8492
rect 26145 8483 26203 8489
rect 26145 8480 26157 8483
rect 26016 8452 26157 8480
rect 26016 8440 26022 8452
rect 26145 8449 26157 8452
rect 26191 8480 26203 8483
rect 27249 8483 27307 8489
rect 27249 8480 27261 8483
rect 26191 8452 27261 8480
rect 26191 8449 26203 8452
rect 26145 8443 26203 8449
rect 27249 8449 27261 8452
rect 27295 8449 27307 8483
rect 27249 8443 27307 8449
rect 28629 8483 28687 8489
rect 28629 8449 28641 8483
rect 28675 8480 28687 8483
rect 29638 8480 29644 8492
rect 28675 8452 29644 8480
rect 28675 8449 28687 8452
rect 28629 8443 28687 8449
rect 29638 8440 29644 8452
rect 29696 8480 29702 8492
rect 30466 8480 30472 8492
rect 29696 8452 30472 8480
rect 29696 8440 29702 8452
rect 30466 8440 30472 8452
rect 30524 8440 30530 8492
rect 31021 8483 31079 8489
rect 31021 8449 31033 8483
rect 31067 8449 31079 8483
rect 31021 8443 31079 8449
rect 31389 8483 31447 8489
rect 31389 8449 31401 8483
rect 31435 8480 31447 8483
rect 31570 8480 31576 8492
rect 31435 8452 31576 8480
rect 31435 8449 31447 8452
rect 31389 8443 31447 8449
rect 23569 8347 23627 8353
rect 23569 8313 23581 8347
rect 23615 8344 23627 8347
rect 23842 8344 23848 8356
rect 23615 8316 23848 8344
rect 23615 8313 23627 8316
rect 23569 8307 23627 8313
rect 23842 8304 23848 8316
rect 23900 8304 23906 8356
rect 27154 8304 27160 8356
rect 27212 8344 27218 8356
rect 27522 8344 27528 8356
rect 27212 8316 27528 8344
rect 27212 8304 27218 8316
rect 27522 8304 27528 8316
rect 27580 8344 27586 8356
rect 29270 8344 29276 8356
rect 27580 8316 29276 8344
rect 27580 8304 27586 8316
rect 29270 8304 29276 8316
rect 29328 8344 29334 8356
rect 29917 8347 29975 8353
rect 29917 8344 29929 8347
rect 29328 8316 29929 8344
rect 29328 8304 29334 8316
rect 29917 8313 29929 8316
rect 29963 8313 29975 8347
rect 31036 8344 31064 8443
rect 31570 8440 31576 8452
rect 31628 8440 31634 8492
rect 34609 8483 34667 8489
rect 34609 8449 34621 8483
rect 34655 8449 34667 8483
rect 34609 8443 34667 8449
rect 31205 8415 31263 8421
rect 31205 8381 31217 8415
rect 31251 8412 31263 8415
rect 31478 8412 31484 8424
rect 31251 8384 31484 8412
rect 31251 8381 31263 8384
rect 31205 8375 31263 8381
rect 31478 8372 31484 8384
rect 31536 8412 31542 8424
rect 31662 8412 31668 8424
rect 31536 8384 31668 8412
rect 31536 8372 31542 8384
rect 31662 8372 31668 8384
rect 31720 8372 31726 8424
rect 34514 8372 34520 8424
rect 34572 8372 34578 8424
rect 34624 8412 34652 8443
rect 35434 8440 35440 8492
rect 35492 8440 35498 8492
rect 35802 8440 35808 8492
rect 35860 8440 35866 8492
rect 36354 8440 36360 8492
rect 36412 8480 36418 8492
rect 36412 8452 38332 8480
rect 36412 8440 36418 8452
rect 35986 8412 35992 8424
rect 34624 8384 35992 8412
rect 35986 8372 35992 8384
rect 36044 8412 36050 8424
rect 36538 8412 36544 8424
rect 36044 8384 36544 8412
rect 36044 8372 36050 8384
rect 36538 8372 36544 8384
rect 36596 8372 36602 8424
rect 31754 8344 31760 8356
rect 31036 8316 31760 8344
rect 29917 8307 29975 8313
rect 31754 8304 31760 8316
rect 31812 8304 31818 8356
rect 34146 8304 34152 8356
rect 34204 8344 34210 8356
rect 36262 8344 36268 8356
rect 34204 8316 36268 8344
rect 34204 8304 34210 8316
rect 36262 8304 36268 8316
rect 36320 8304 36326 8356
rect 36633 8347 36691 8353
rect 36633 8313 36645 8347
rect 36679 8344 36691 8347
rect 38010 8344 38016 8356
rect 36679 8316 38016 8344
rect 36679 8313 36691 8316
rect 36633 8307 36691 8313
rect 38010 8304 38016 8316
rect 38068 8304 38074 8356
rect 38304 8344 38332 8452
rect 38562 8440 38568 8492
rect 38620 8440 38626 8492
rect 39669 8483 39727 8489
rect 39669 8449 39681 8483
rect 39715 8449 39727 8483
rect 39669 8443 39727 8449
rect 39684 8412 39712 8443
rect 39758 8440 39764 8492
rect 39816 8440 39822 8492
rect 39868 8489 39896 8520
rect 40126 8508 40132 8560
rect 40184 8548 40190 8560
rect 41800 8557 41828 8588
rect 42702 8576 42708 8588
rect 42760 8576 42766 8628
rect 42886 8576 42892 8628
rect 42944 8576 42950 8628
rect 44174 8576 44180 8628
rect 44232 8576 44238 8628
rect 40497 8551 40555 8557
rect 40497 8548 40509 8551
rect 40184 8520 40509 8548
rect 40184 8508 40190 8520
rect 40497 8517 40509 8520
rect 40543 8548 40555 8551
rect 41785 8551 41843 8557
rect 41785 8548 41797 8551
rect 40543 8520 41797 8548
rect 40543 8517 40555 8520
rect 40497 8511 40555 8517
rect 41785 8517 41797 8520
rect 41831 8517 41843 8551
rect 41785 8511 41843 8517
rect 41969 8551 42027 8557
rect 41969 8517 41981 8551
rect 42015 8548 42027 8551
rect 42981 8551 43039 8557
rect 42981 8548 42993 8551
rect 42015 8520 42993 8548
rect 42015 8517 42027 8520
rect 41969 8511 42027 8517
rect 42981 8517 42993 8520
rect 43027 8517 43039 8551
rect 42981 8511 43039 8517
rect 39853 8483 39911 8489
rect 39853 8449 39865 8483
rect 39899 8449 39911 8483
rect 39853 8443 39911 8449
rect 39942 8440 39948 8492
rect 40000 8480 40006 8492
rect 40037 8483 40095 8489
rect 40037 8480 40049 8483
rect 40000 8452 40049 8480
rect 40000 8440 40006 8452
rect 40037 8449 40049 8452
rect 40083 8449 40095 8483
rect 40037 8443 40095 8449
rect 40954 8440 40960 8492
rect 41012 8440 41018 8492
rect 41322 8440 41328 8492
rect 41380 8480 41386 8492
rect 41601 8483 41659 8489
rect 41601 8480 41613 8483
rect 41380 8452 41613 8480
rect 41380 8440 41386 8452
rect 41601 8449 41613 8452
rect 41647 8449 41659 8483
rect 41601 8443 41659 8449
rect 41690 8440 41696 8492
rect 41748 8480 41754 8492
rect 42797 8483 42855 8489
rect 42797 8480 42809 8483
rect 41748 8452 42809 8480
rect 41748 8440 41754 8452
rect 42797 8449 42809 8452
rect 42843 8449 42855 8483
rect 42797 8443 42855 8449
rect 44358 8440 44364 8492
rect 44416 8440 44422 8492
rect 40865 8415 40923 8421
rect 40865 8412 40877 8415
rect 39684 8384 40877 8412
rect 40865 8381 40877 8384
rect 40911 8412 40923 8415
rect 41046 8412 41052 8424
rect 40911 8384 41052 8412
rect 40911 8381 40923 8384
rect 40865 8375 40923 8381
rect 41046 8372 41052 8384
rect 41104 8372 41110 8424
rect 41141 8347 41199 8353
rect 41141 8344 41153 8347
rect 38304 8316 41153 8344
rect 41141 8313 41153 8316
rect 41187 8313 41199 8347
rect 41141 8307 41199 8313
rect 42613 8347 42671 8353
rect 42613 8313 42625 8347
rect 42659 8313 42671 8347
rect 42613 8307 42671 8313
rect 11572 8248 13032 8276
rect 11572 8236 11578 8248
rect 18598 8236 18604 8288
rect 18656 8236 18662 8288
rect 29178 8236 29184 8288
rect 29236 8276 29242 8288
rect 36170 8276 36176 8288
rect 29236 8248 36176 8276
rect 29236 8236 29242 8248
rect 36170 8236 36176 8248
rect 36228 8236 36234 8288
rect 36446 8236 36452 8288
rect 36504 8236 36510 8288
rect 38654 8236 38660 8288
rect 38712 8236 38718 8288
rect 40402 8236 40408 8288
rect 40460 8276 40466 8288
rect 40589 8279 40647 8285
rect 40589 8276 40601 8279
rect 40460 8248 40601 8276
rect 40460 8236 40466 8248
rect 40589 8245 40601 8248
rect 40635 8245 40647 8279
rect 40589 8239 40647 8245
rect 41046 8236 41052 8288
rect 41104 8276 41110 8288
rect 42628 8276 42656 8307
rect 41104 8248 42656 8276
rect 41104 8236 41110 8248
rect 43162 8236 43168 8288
rect 43220 8236 43226 8288
rect 1104 8186 44896 8208
rect 1104 8134 6423 8186
rect 6475 8134 6487 8186
rect 6539 8134 6551 8186
rect 6603 8134 6615 8186
rect 6667 8134 6679 8186
rect 6731 8134 17370 8186
rect 17422 8134 17434 8186
rect 17486 8134 17498 8186
rect 17550 8134 17562 8186
rect 17614 8134 17626 8186
rect 17678 8134 28317 8186
rect 28369 8134 28381 8186
rect 28433 8134 28445 8186
rect 28497 8134 28509 8186
rect 28561 8134 28573 8186
rect 28625 8134 39264 8186
rect 39316 8134 39328 8186
rect 39380 8134 39392 8186
rect 39444 8134 39456 8186
rect 39508 8134 39520 8186
rect 39572 8134 44896 8186
rect 1104 8112 44896 8134
rect 6270 8032 6276 8084
rect 6328 8072 6334 8084
rect 6549 8075 6607 8081
rect 6549 8072 6561 8075
rect 6328 8044 6561 8072
rect 6328 8032 6334 8044
rect 6549 8041 6561 8044
rect 6595 8041 6607 8075
rect 9769 8075 9827 8081
rect 6549 8035 6607 8041
rect 6886 8044 9628 8072
rect 1581 8007 1639 8013
rect 1581 7973 1593 8007
rect 1627 8004 1639 8007
rect 6886 8004 6914 8044
rect 8202 8004 8208 8016
rect 1627 7976 6914 8004
rect 7852 7976 8208 8004
rect 1627 7973 1639 7976
rect 1581 7967 1639 7973
rect 3142 7896 3148 7948
rect 3200 7896 3206 7948
rect 3329 7939 3387 7945
rect 3329 7905 3341 7939
rect 3375 7936 3387 7939
rect 3375 7908 5212 7936
rect 3375 7905 3387 7908
rect 3329 7899 3387 7905
rect 934 7828 940 7880
rect 992 7868 998 7880
rect 1765 7871 1823 7877
rect 1765 7868 1777 7871
rect 992 7840 1777 7868
rect 992 7828 998 7840
rect 1765 7837 1777 7840
rect 1811 7837 1823 7871
rect 1765 7831 1823 7837
rect 5184 7800 5212 7908
rect 5261 7871 5319 7877
rect 5261 7837 5273 7871
rect 5307 7868 5319 7871
rect 5534 7868 5540 7880
rect 5307 7840 5540 7868
rect 5307 7837 5319 7840
rect 5261 7831 5319 7837
rect 5534 7828 5540 7840
rect 5592 7828 5598 7880
rect 5810 7828 5816 7880
rect 5868 7868 5874 7880
rect 7852 7868 7880 7976
rect 8202 7964 8208 7976
rect 8260 8004 8266 8016
rect 8260 7976 8432 8004
rect 8260 7964 8266 7976
rect 7926 7896 7932 7948
rect 7984 7936 7990 7948
rect 8404 7945 8432 7976
rect 8297 7939 8355 7945
rect 8297 7936 8309 7939
rect 7984 7908 8309 7936
rect 7984 7896 7990 7908
rect 8297 7905 8309 7908
rect 8343 7905 8355 7939
rect 8297 7899 8355 7905
rect 8389 7939 8447 7945
rect 8389 7905 8401 7939
rect 8435 7905 8447 7939
rect 8389 7899 8447 7905
rect 5868 7840 7880 7868
rect 5868 7828 5874 7840
rect 5442 7800 5448 7812
rect 5184 7772 5448 7800
rect 5442 7760 5448 7772
rect 5500 7800 5506 7812
rect 5828 7800 5856 7828
rect 5500 7772 5856 7800
rect 8205 7803 8263 7809
rect 5500 7760 5506 7772
rect 8205 7769 8217 7803
rect 8251 7800 8263 7803
rect 9122 7800 9128 7812
rect 8251 7772 9128 7800
rect 8251 7769 8263 7772
rect 8205 7763 8263 7769
rect 9122 7760 9128 7772
rect 9180 7760 9186 7812
rect 2685 7735 2743 7741
rect 2685 7701 2697 7735
rect 2731 7732 2743 7735
rect 2958 7732 2964 7744
rect 2731 7704 2964 7732
rect 2731 7701 2743 7704
rect 2685 7695 2743 7701
rect 2958 7692 2964 7704
rect 3016 7692 3022 7744
rect 3053 7735 3111 7741
rect 3053 7701 3065 7735
rect 3099 7732 3111 7735
rect 5258 7732 5264 7744
rect 3099 7704 5264 7732
rect 3099 7701 3111 7704
rect 3053 7695 3111 7701
rect 5258 7692 5264 7704
rect 5316 7692 5322 7744
rect 7282 7692 7288 7744
rect 7340 7732 7346 7744
rect 7837 7735 7895 7741
rect 7837 7732 7849 7735
rect 7340 7704 7849 7732
rect 7340 7692 7346 7704
rect 7837 7701 7849 7704
rect 7883 7701 7895 7735
rect 9600 7732 9628 8044
rect 9769 8041 9781 8075
rect 9815 8072 9827 8075
rect 10502 8072 10508 8084
rect 9815 8044 10508 8072
rect 9815 8041 9827 8044
rect 9769 8035 9827 8041
rect 10502 8032 10508 8044
rect 10560 8032 10566 8084
rect 10870 8032 10876 8084
rect 10928 8072 10934 8084
rect 10928 8044 11928 8072
rect 10928 8032 10934 8044
rect 11900 8013 11928 8044
rect 16206 8032 16212 8084
rect 16264 8032 16270 8084
rect 17773 8075 17831 8081
rect 17773 8041 17785 8075
rect 17819 8072 17831 8075
rect 18230 8072 18236 8084
rect 17819 8044 18236 8072
rect 17819 8041 17831 8044
rect 17773 8035 17831 8041
rect 18230 8032 18236 8044
rect 18288 8032 18294 8084
rect 20070 8072 20076 8084
rect 18340 8044 20076 8072
rect 11885 8007 11943 8013
rect 11885 7973 11897 8007
rect 11931 7973 11943 8007
rect 11885 7967 11943 7973
rect 11900 7936 11928 7967
rect 13081 7939 13139 7945
rect 13081 7936 13093 7939
rect 11900 7908 13093 7936
rect 13081 7905 13093 7908
rect 13127 7936 13139 7939
rect 13538 7936 13544 7948
rect 13127 7908 13544 7936
rect 13127 7905 13139 7908
rect 13081 7899 13139 7905
rect 13538 7896 13544 7908
rect 13596 7896 13602 7948
rect 18340 7945 18368 8044
rect 20070 8032 20076 8044
rect 20128 8032 20134 8084
rect 22462 8032 22468 8084
rect 22520 8072 22526 8084
rect 22557 8075 22615 8081
rect 22557 8072 22569 8075
rect 22520 8044 22569 8072
rect 22520 8032 22526 8044
rect 22557 8041 22569 8044
rect 22603 8041 22615 8075
rect 22557 8035 22615 8041
rect 27982 8032 27988 8084
rect 28040 8072 28046 8084
rect 28629 8075 28687 8081
rect 28629 8072 28641 8075
rect 28040 8044 28641 8072
rect 28040 8032 28046 8044
rect 28629 8041 28641 8044
rect 28675 8041 28687 8075
rect 32309 8075 32367 8081
rect 32309 8072 32321 8075
rect 28629 8035 28687 8041
rect 31680 8044 32321 8072
rect 31570 7964 31576 8016
rect 31628 8004 31634 8016
rect 31680 8013 31708 8044
rect 32309 8041 32321 8044
rect 32355 8041 32367 8075
rect 32309 8035 32367 8041
rect 32493 8075 32551 8081
rect 32493 8041 32505 8075
rect 32539 8072 32551 8075
rect 32950 8072 32956 8084
rect 32539 8044 32956 8072
rect 32539 8041 32551 8044
rect 32493 8035 32551 8041
rect 32950 8032 32956 8044
rect 33008 8032 33014 8084
rect 34241 8075 34299 8081
rect 34241 8041 34253 8075
rect 34287 8072 34299 8075
rect 36446 8072 36452 8084
rect 34287 8044 36452 8072
rect 34287 8041 34299 8044
rect 34241 8035 34299 8041
rect 36446 8032 36452 8044
rect 36504 8032 36510 8084
rect 36538 8032 36544 8084
rect 36596 8032 36602 8084
rect 36998 8032 37004 8084
rect 37056 8032 37062 8084
rect 37366 8032 37372 8084
rect 37424 8032 37430 8084
rect 39390 8032 39396 8084
rect 39448 8072 39454 8084
rect 41877 8075 41935 8081
rect 41877 8072 41889 8075
rect 39448 8044 41889 8072
rect 39448 8032 39454 8044
rect 41877 8041 41889 8044
rect 41923 8041 41935 8075
rect 41877 8035 41935 8041
rect 42337 8075 42395 8081
rect 42337 8041 42349 8075
rect 42383 8072 42395 8075
rect 42794 8072 42800 8084
rect 42383 8044 42800 8072
rect 42383 8041 42395 8044
rect 42337 8035 42395 8041
rect 42794 8032 42800 8044
rect 42852 8032 42858 8084
rect 31665 8007 31723 8013
rect 31665 8004 31677 8007
rect 31628 7976 31677 8004
rect 31628 7964 31634 7976
rect 31665 7973 31677 7976
rect 31711 7973 31723 8007
rect 31665 7967 31723 7973
rect 36170 7964 36176 8016
rect 36228 8004 36234 8016
rect 36228 7976 39436 8004
rect 36228 7964 36234 7976
rect 18325 7939 18383 7945
rect 18325 7936 18337 7939
rect 16776 7908 18337 7936
rect 9677 7871 9735 7877
rect 9677 7837 9689 7871
rect 9723 7868 9735 7871
rect 9858 7868 9864 7880
rect 9723 7840 9864 7868
rect 9723 7837 9735 7840
rect 9677 7831 9735 7837
rect 9858 7828 9864 7840
rect 9916 7828 9922 7880
rect 10505 7871 10563 7877
rect 10505 7837 10517 7871
rect 10551 7868 10563 7871
rect 10594 7868 10600 7880
rect 10551 7840 10600 7868
rect 10551 7837 10563 7840
rect 10505 7831 10563 7837
rect 10594 7828 10600 7840
rect 10652 7828 10658 7880
rect 12805 7871 12863 7877
rect 12805 7837 12817 7871
rect 12851 7868 12863 7871
rect 12894 7868 12900 7880
rect 12851 7840 12900 7868
rect 12851 7837 12863 7840
rect 12805 7831 12863 7837
rect 12894 7828 12900 7840
rect 12952 7828 12958 7880
rect 14829 7871 14887 7877
rect 14829 7837 14841 7871
rect 14875 7868 14887 7871
rect 14918 7868 14924 7880
rect 14875 7840 14924 7868
rect 14875 7837 14887 7840
rect 14829 7831 14887 7837
rect 14918 7828 14924 7840
rect 14976 7828 14982 7880
rect 15470 7868 15476 7880
rect 15028 7840 15476 7868
rect 9766 7760 9772 7812
rect 9824 7800 9830 7812
rect 10750 7803 10808 7809
rect 10750 7800 10762 7803
rect 9824 7772 10762 7800
rect 9824 7760 9830 7772
rect 10750 7769 10762 7772
rect 10796 7769 10808 7803
rect 15028 7800 15056 7840
rect 15470 7828 15476 7840
rect 15528 7828 15534 7880
rect 15654 7828 15660 7880
rect 15712 7868 15718 7880
rect 16776 7868 16804 7908
rect 18325 7905 18337 7908
rect 18371 7905 18383 7939
rect 18325 7899 18383 7905
rect 19886 7896 19892 7948
rect 19944 7896 19950 7948
rect 26142 7936 26148 7948
rect 25792 7908 26148 7936
rect 15712 7840 16804 7868
rect 15712 7828 15718 7840
rect 16850 7828 16856 7880
rect 16908 7828 16914 7880
rect 18141 7871 18199 7877
rect 18141 7837 18153 7871
rect 18187 7868 18199 7871
rect 18598 7868 18604 7880
rect 18187 7840 18604 7868
rect 18187 7837 18199 7840
rect 18141 7831 18199 7837
rect 18598 7828 18604 7840
rect 18656 7828 18662 7880
rect 19518 7828 19524 7880
rect 19576 7868 19582 7880
rect 20145 7871 20203 7877
rect 20145 7868 20157 7871
rect 19576 7840 20157 7868
rect 19576 7828 19582 7840
rect 20145 7837 20157 7840
rect 20191 7837 20203 7871
rect 20145 7831 20203 7837
rect 21910 7828 21916 7880
rect 21968 7828 21974 7880
rect 22741 7871 22799 7877
rect 22741 7837 22753 7871
rect 22787 7868 22799 7871
rect 23382 7868 23388 7880
rect 22787 7840 23388 7868
rect 22787 7837 22799 7840
rect 22741 7831 22799 7837
rect 23382 7828 23388 7840
rect 23440 7828 23446 7880
rect 23477 7871 23535 7877
rect 23477 7837 23489 7871
rect 23523 7868 23535 7871
rect 23566 7868 23572 7880
rect 23523 7840 23572 7868
rect 23523 7837 23535 7840
rect 23477 7831 23535 7837
rect 23566 7828 23572 7840
rect 23624 7828 23630 7880
rect 25792 7877 25820 7908
rect 26142 7896 26148 7908
rect 26200 7896 26206 7948
rect 26237 7939 26295 7945
rect 26237 7905 26249 7939
rect 26283 7936 26295 7939
rect 27154 7936 27160 7948
rect 26283 7908 27160 7936
rect 26283 7905 26295 7908
rect 26237 7899 26295 7905
rect 27154 7896 27160 7908
rect 27212 7896 27218 7948
rect 27890 7896 27896 7948
rect 27948 7936 27954 7948
rect 28077 7939 28135 7945
rect 28077 7936 28089 7939
rect 27948 7908 28089 7936
rect 27948 7896 27954 7908
rect 28077 7905 28089 7908
rect 28123 7936 28135 7939
rect 28902 7936 28908 7948
rect 28123 7908 28908 7936
rect 28123 7905 28135 7908
rect 28077 7899 28135 7905
rect 28902 7896 28908 7908
rect 28960 7896 28966 7948
rect 34072 7908 34284 7936
rect 25777 7871 25835 7877
rect 25777 7837 25789 7871
rect 25823 7837 25835 7871
rect 26605 7871 26663 7877
rect 26605 7868 26617 7871
rect 25777 7831 25835 7837
rect 26160 7840 26617 7868
rect 10750 7763 10808 7769
rect 10888 7772 15056 7800
rect 15096 7803 15154 7809
rect 10888 7732 10916 7772
rect 15096 7769 15108 7803
rect 15142 7800 15154 7803
rect 15142 7772 16712 7800
rect 15142 7769 15154 7772
rect 15096 7763 15154 7769
rect 9600 7704 10916 7732
rect 7837 7695 7895 7701
rect 12250 7692 12256 7744
rect 12308 7732 12314 7744
rect 12437 7735 12495 7741
rect 12437 7732 12449 7735
rect 12308 7704 12449 7732
rect 12308 7692 12314 7704
rect 12437 7701 12449 7704
rect 12483 7701 12495 7735
rect 12437 7695 12495 7701
rect 12894 7692 12900 7744
rect 12952 7692 12958 7744
rect 16684 7741 16712 7772
rect 17954 7760 17960 7812
rect 18012 7800 18018 7812
rect 18233 7803 18291 7809
rect 18233 7800 18245 7803
rect 18012 7772 18245 7800
rect 18012 7760 18018 7772
rect 18233 7769 18245 7772
rect 18279 7769 18291 7803
rect 26160 7800 26188 7840
rect 26605 7837 26617 7840
rect 26651 7837 26663 7871
rect 26605 7831 26663 7837
rect 27430 7828 27436 7880
rect 27488 7868 27494 7880
rect 28629 7871 28687 7877
rect 28629 7868 28641 7871
rect 27488 7840 28641 7868
rect 27488 7828 27494 7840
rect 28629 7837 28641 7840
rect 28675 7868 28687 7871
rect 29638 7868 29644 7880
rect 28675 7840 29644 7868
rect 28675 7837 28687 7840
rect 28629 7831 28687 7837
rect 29638 7828 29644 7840
rect 29696 7828 29702 7880
rect 29730 7828 29736 7880
rect 29788 7868 29794 7880
rect 30285 7871 30343 7877
rect 30285 7868 30297 7871
rect 29788 7840 30297 7868
rect 29788 7828 29794 7840
rect 30285 7837 30297 7840
rect 30331 7837 30343 7871
rect 30285 7831 30343 7837
rect 32582 7828 32588 7880
rect 32640 7868 32646 7880
rect 34072 7877 34100 7908
rect 34057 7871 34115 7877
rect 34057 7868 34069 7871
rect 32640 7840 34069 7868
rect 32640 7828 32646 7840
rect 34057 7837 34069 7840
rect 34103 7837 34115 7871
rect 34057 7831 34115 7837
rect 34149 7871 34207 7877
rect 34149 7837 34161 7871
rect 34195 7837 34207 7871
rect 34256 7868 34284 7908
rect 34330 7896 34336 7948
rect 34388 7896 34394 7948
rect 38654 7936 38660 7948
rect 37016 7908 38660 7936
rect 35066 7868 35072 7880
rect 34256 7840 35072 7868
rect 34149 7831 34207 7837
rect 27798 7800 27804 7812
rect 18233 7763 18291 7769
rect 25608 7772 26188 7800
rect 27646 7772 27804 7800
rect 16669 7735 16727 7741
rect 16669 7701 16681 7735
rect 16715 7701 16727 7735
rect 16669 7695 16727 7701
rect 21266 7692 21272 7744
rect 21324 7692 21330 7744
rect 21726 7692 21732 7744
rect 21784 7692 21790 7744
rect 23293 7735 23351 7741
rect 23293 7701 23305 7735
rect 23339 7732 23351 7735
rect 23382 7732 23388 7744
rect 23339 7704 23388 7732
rect 23339 7701 23351 7704
rect 23293 7695 23351 7701
rect 23382 7692 23388 7704
rect 23440 7692 23446 7744
rect 25608 7741 25636 7772
rect 27798 7760 27804 7772
rect 27856 7760 27862 7812
rect 30558 7809 30564 7812
rect 30552 7763 30564 7809
rect 30558 7760 30564 7763
rect 30616 7760 30622 7812
rect 31938 7760 31944 7812
rect 31996 7800 32002 7812
rect 32125 7803 32183 7809
rect 32125 7800 32137 7803
rect 31996 7772 32137 7800
rect 31996 7760 32002 7772
rect 32125 7769 32137 7772
rect 32171 7769 32183 7803
rect 34164 7800 34192 7831
rect 35066 7828 35072 7840
rect 35124 7828 35130 7880
rect 35158 7828 35164 7880
rect 35216 7828 35222 7880
rect 37016 7877 37044 7908
rect 38654 7896 38660 7908
rect 38712 7936 38718 7948
rect 38712 7908 39252 7936
rect 38712 7896 38718 7908
rect 37001 7871 37059 7877
rect 37001 7868 37013 7871
rect 35360 7840 37013 7868
rect 35360 7800 35388 7840
rect 37001 7837 37013 7840
rect 37047 7837 37059 7871
rect 37001 7831 37059 7837
rect 37090 7828 37096 7880
rect 37148 7828 37154 7880
rect 37182 7828 37188 7880
rect 37240 7868 37246 7880
rect 37240 7840 37964 7868
rect 37240 7828 37246 7840
rect 34164 7772 35388 7800
rect 35428 7803 35486 7809
rect 32125 7763 32183 7769
rect 35428 7769 35440 7803
rect 35474 7800 35486 7803
rect 37936 7800 37964 7840
rect 38010 7828 38016 7880
rect 38068 7828 38074 7880
rect 38746 7828 38752 7880
rect 38804 7868 38810 7880
rect 39224 7877 39252 7908
rect 39117 7871 39175 7877
rect 39117 7868 39129 7871
rect 38804 7840 39129 7868
rect 38804 7828 38810 7840
rect 39117 7837 39129 7840
rect 39163 7837 39175 7871
rect 39117 7831 39175 7837
rect 39209 7871 39267 7877
rect 39209 7837 39221 7871
rect 39255 7837 39267 7871
rect 39209 7831 39267 7837
rect 39298 7828 39304 7880
rect 39356 7828 39362 7880
rect 39408 7868 39436 7976
rect 40494 7896 40500 7948
rect 40552 7896 40558 7948
rect 39485 7871 39543 7877
rect 39485 7868 39497 7871
rect 39408 7840 39497 7868
rect 39485 7837 39497 7840
rect 39531 7868 39543 7871
rect 41046 7868 41052 7880
rect 39531 7840 41052 7868
rect 39531 7837 39543 7840
rect 39485 7831 39543 7837
rect 41046 7828 41052 7840
rect 41104 7828 41110 7880
rect 42521 7871 42579 7877
rect 42521 7837 42533 7871
rect 42567 7868 42579 7871
rect 43162 7868 43168 7880
rect 42567 7840 43168 7868
rect 42567 7837 42579 7840
rect 42521 7831 42579 7837
rect 43162 7828 43168 7840
rect 43220 7828 43226 7880
rect 44358 7828 44364 7880
rect 44416 7828 44422 7880
rect 39574 7800 39580 7812
rect 35474 7772 37872 7800
rect 37936 7772 39580 7800
rect 35474 7769 35486 7772
rect 35428 7763 35486 7769
rect 25593 7735 25651 7741
rect 25593 7701 25605 7735
rect 25639 7701 25651 7735
rect 25593 7695 25651 7701
rect 32335 7735 32393 7741
rect 32335 7701 32347 7735
rect 32381 7732 32393 7735
rect 34422 7732 34428 7744
rect 32381 7704 34428 7732
rect 32381 7701 32393 7704
rect 32335 7695 32393 7701
rect 34422 7692 34428 7704
rect 34480 7692 34486 7744
rect 36262 7692 36268 7744
rect 36320 7732 36326 7744
rect 37182 7732 37188 7744
rect 36320 7704 37188 7732
rect 36320 7692 36326 7704
rect 37182 7692 37188 7704
rect 37240 7692 37246 7744
rect 37844 7741 37872 7772
rect 39574 7760 39580 7772
rect 39632 7760 39638 7812
rect 40764 7803 40822 7809
rect 40764 7769 40776 7803
rect 40810 7800 40822 7803
rect 41414 7800 41420 7812
rect 40810 7772 41420 7800
rect 40810 7769 40822 7772
rect 40764 7763 40822 7769
rect 41414 7760 41420 7772
rect 41472 7760 41478 7812
rect 37829 7735 37887 7741
rect 37829 7701 37841 7735
rect 37875 7701 37887 7735
rect 37829 7695 37887 7701
rect 38841 7735 38899 7741
rect 38841 7701 38853 7735
rect 38887 7732 38899 7735
rect 41598 7732 41604 7744
rect 38887 7704 41604 7732
rect 38887 7701 38899 7704
rect 38841 7695 38899 7701
rect 41598 7692 41604 7704
rect 41656 7692 41662 7744
rect 43438 7692 43444 7744
rect 43496 7732 43502 7744
rect 44177 7735 44235 7741
rect 44177 7732 44189 7735
rect 43496 7704 44189 7732
rect 43496 7692 43502 7704
rect 44177 7701 44189 7704
rect 44223 7701 44235 7735
rect 44177 7695 44235 7701
rect 1104 7642 45051 7664
rect 1104 7590 11896 7642
rect 11948 7590 11960 7642
rect 12012 7590 12024 7642
rect 12076 7590 12088 7642
rect 12140 7590 12152 7642
rect 12204 7590 22843 7642
rect 22895 7590 22907 7642
rect 22959 7590 22971 7642
rect 23023 7590 23035 7642
rect 23087 7590 23099 7642
rect 23151 7590 33790 7642
rect 33842 7590 33854 7642
rect 33906 7590 33918 7642
rect 33970 7590 33982 7642
rect 34034 7590 34046 7642
rect 34098 7590 44737 7642
rect 44789 7590 44801 7642
rect 44853 7590 44865 7642
rect 44917 7590 44929 7642
rect 44981 7590 44993 7642
rect 45045 7590 45051 7642
rect 1104 7568 45051 7590
rect 3881 7531 3939 7537
rect 3881 7497 3893 7531
rect 3927 7528 3939 7531
rect 3970 7528 3976 7540
rect 3927 7500 3976 7528
rect 3927 7497 3939 7500
rect 3881 7491 3939 7497
rect 3970 7488 3976 7500
rect 4028 7488 4034 7540
rect 5261 7531 5319 7537
rect 5261 7497 5273 7531
rect 5307 7528 5319 7531
rect 5350 7528 5356 7540
rect 5307 7500 5356 7528
rect 5307 7497 5319 7500
rect 5261 7491 5319 7497
rect 5350 7488 5356 7500
rect 5408 7488 5414 7540
rect 9122 7488 9128 7540
rect 9180 7488 9186 7540
rect 11701 7531 11759 7537
rect 11701 7497 11713 7531
rect 11747 7528 11759 7531
rect 11790 7528 11796 7540
rect 11747 7500 11796 7528
rect 11747 7497 11759 7500
rect 11701 7491 11759 7497
rect 11790 7488 11796 7500
rect 11848 7488 11854 7540
rect 12437 7531 12495 7537
rect 12437 7497 12449 7531
rect 12483 7528 12495 7531
rect 14458 7528 14464 7540
rect 12483 7500 14464 7528
rect 12483 7497 12495 7500
rect 12437 7491 12495 7497
rect 14458 7488 14464 7500
rect 14516 7488 14522 7540
rect 31021 7531 31079 7537
rect 31021 7497 31033 7531
rect 31067 7528 31079 7531
rect 31110 7528 31116 7540
rect 31067 7500 31116 7528
rect 31067 7497 31079 7500
rect 31021 7491 31079 7497
rect 31110 7488 31116 7500
rect 31168 7488 31174 7540
rect 31386 7488 31392 7540
rect 31444 7488 31450 7540
rect 32950 7528 32956 7540
rect 31496 7500 32956 7528
rect 2593 7463 2651 7469
rect 2593 7429 2605 7463
rect 2639 7460 2651 7463
rect 5534 7460 5540 7472
rect 2639 7432 5540 7460
rect 2639 7429 2651 7432
rect 2593 7423 2651 7429
rect 5534 7420 5540 7432
rect 5592 7420 5598 7472
rect 6914 7420 6920 7472
rect 6972 7460 6978 7472
rect 14918 7460 14924 7472
rect 6972 7432 7788 7460
rect 6972 7420 6978 7432
rect 7760 7404 7788 7432
rect 13280 7432 14924 7460
rect 2133 7395 2191 7401
rect 2133 7361 2145 7395
rect 2179 7392 2191 7395
rect 2179 7364 4844 7392
rect 2179 7361 2191 7364
rect 2133 7355 2191 7361
rect 4816 7265 4844 7364
rect 5166 7352 5172 7404
rect 5224 7352 5230 7404
rect 7282 7352 7288 7404
rect 7340 7352 7346 7404
rect 7742 7352 7748 7404
rect 7800 7352 7806 7404
rect 8001 7395 8059 7401
rect 8001 7392 8013 7395
rect 7852 7364 8013 7392
rect 5074 7284 5080 7336
rect 5132 7324 5138 7336
rect 5442 7324 5448 7336
rect 5132 7296 5448 7324
rect 5132 7284 5138 7296
rect 5442 7284 5448 7296
rect 5500 7284 5506 7336
rect 7852 7324 7880 7364
rect 8001 7361 8013 7364
rect 8047 7361 8059 7395
rect 9858 7392 9864 7404
rect 9916 7396 9922 7404
rect 9819 7364 9864 7392
rect 8001 7355 8059 7361
rect 9858 7352 9864 7364
rect 9916 7392 9996 7396
rect 10965 7395 11023 7401
rect 10965 7392 10977 7395
rect 9916 7368 10977 7392
rect 9916 7352 9922 7368
rect 9968 7364 10977 7368
rect 10965 7361 10977 7364
rect 11011 7361 11023 7395
rect 10965 7355 11023 7361
rect 11885 7395 11943 7401
rect 11885 7361 11897 7395
rect 11931 7392 11943 7395
rect 12250 7392 12256 7404
rect 11931 7364 12256 7392
rect 11931 7361 11943 7364
rect 11885 7355 11943 7361
rect 7116 7296 7880 7324
rect 10980 7324 11008 7355
rect 12250 7352 12256 7364
rect 12308 7352 12314 7404
rect 12345 7395 12403 7401
rect 12345 7361 12357 7395
rect 12391 7392 12403 7395
rect 12618 7392 12624 7404
rect 12391 7364 12624 7392
rect 12391 7361 12403 7364
rect 12345 7355 12403 7361
rect 12360 7324 12388 7355
rect 12618 7352 12624 7364
rect 12676 7352 12682 7404
rect 13280 7401 13308 7432
rect 14918 7420 14924 7432
rect 14976 7420 14982 7472
rect 20156 7463 20214 7469
rect 20156 7429 20168 7463
rect 20202 7460 20214 7463
rect 21726 7460 21732 7472
rect 20202 7432 21732 7460
rect 20202 7429 20214 7432
rect 20156 7423 20214 7429
rect 21726 7420 21732 7432
rect 21784 7420 21790 7472
rect 23382 7469 23388 7472
rect 23376 7460 23388 7469
rect 23343 7432 23388 7460
rect 23376 7423 23388 7432
rect 23382 7420 23388 7423
rect 23440 7420 23446 7472
rect 27890 7420 27896 7472
rect 27948 7420 27954 7472
rect 28902 7420 28908 7472
rect 28960 7460 28966 7472
rect 28960 7432 30328 7460
rect 28960 7420 28966 7432
rect 13265 7395 13323 7401
rect 13265 7361 13277 7395
rect 13311 7361 13323 7395
rect 13265 7355 13323 7361
rect 13354 7352 13360 7404
rect 13412 7392 13418 7404
rect 13521 7395 13579 7401
rect 13521 7392 13533 7395
rect 13412 7364 13533 7392
rect 13412 7352 13418 7364
rect 13521 7361 13533 7364
rect 13567 7361 13579 7395
rect 13521 7355 13579 7361
rect 15470 7352 15476 7404
rect 15528 7352 15534 7404
rect 16206 7352 16212 7404
rect 16264 7392 16270 7404
rect 17221 7395 17279 7401
rect 17221 7392 17233 7395
rect 16264 7364 17233 7392
rect 16264 7352 16270 7364
rect 17221 7361 17233 7364
rect 17267 7361 17279 7395
rect 17221 7355 17279 7361
rect 19886 7352 19892 7404
rect 19944 7352 19950 7404
rect 25958 7352 25964 7404
rect 26016 7352 26022 7404
rect 29178 7352 29184 7404
rect 29236 7352 29242 7404
rect 29638 7352 29644 7404
rect 29696 7352 29702 7404
rect 30300 7401 30328 7432
rect 30650 7420 30656 7472
rect 30708 7460 30714 7472
rect 31496 7460 31524 7500
rect 32950 7488 32956 7500
rect 33008 7488 33014 7540
rect 34330 7488 34336 7540
rect 34388 7528 34394 7540
rect 37090 7528 37096 7540
rect 34388 7500 37096 7528
rect 34388 7488 34394 7500
rect 37090 7488 37096 7500
rect 37148 7528 37154 7540
rect 37553 7531 37611 7537
rect 37553 7528 37565 7531
rect 37148 7500 37565 7528
rect 37148 7488 37154 7500
rect 37553 7497 37565 7500
rect 37599 7497 37611 7531
rect 38397 7531 38455 7537
rect 38397 7528 38409 7531
rect 37553 7491 37611 7497
rect 37660 7500 38409 7528
rect 30708 7432 31524 7460
rect 31573 7463 31631 7469
rect 30708 7420 30714 7432
rect 31573 7429 31585 7463
rect 31619 7460 31631 7463
rect 31846 7460 31852 7472
rect 31619 7432 31852 7460
rect 31619 7429 31631 7432
rect 31573 7423 31631 7429
rect 31846 7420 31852 7432
rect 31904 7420 31910 7472
rect 31938 7420 31944 7472
rect 31996 7460 32002 7472
rect 33413 7463 33471 7469
rect 33413 7460 33425 7463
rect 31996 7432 33425 7460
rect 31996 7420 32002 7432
rect 33413 7429 33425 7432
rect 33459 7429 33471 7463
rect 33413 7423 33471 7429
rect 33643 7429 33701 7435
rect 33643 7426 33655 7429
rect 30285 7395 30343 7401
rect 30285 7361 30297 7395
rect 30331 7392 30343 7395
rect 31205 7395 31263 7401
rect 31205 7392 31217 7395
rect 30331 7364 31217 7392
rect 30331 7361 30343 7364
rect 30285 7355 30343 7361
rect 31205 7361 31217 7364
rect 31251 7392 31263 7395
rect 31386 7392 31392 7404
rect 31251 7364 31392 7392
rect 31251 7361 31263 7364
rect 31205 7355 31263 7361
rect 31386 7352 31392 7364
rect 31444 7352 31450 7404
rect 31665 7395 31723 7401
rect 31665 7361 31677 7395
rect 31711 7392 31723 7395
rect 31754 7392 31760 7404
rect 31711 7364 31760 7392
rect 31711 7361 31723 7364
rect 31665 7355 31723 7361
rect 31754 7352 31760 7364
rect 31812 7392 31818 7404
rect 32214 7392 32220 7404
rect 31812 7364 32220 7392
rect 31812 7352 31818 7364
rect 32214 7352 32220 7364
rect 32272 7352 32278 7404
rect 32582 7352 32588 7404
rect 32640 7352 32646 7404
rect 32674 7352 32680 7404
rect 32732 7352 32738 7404
rect 32766 7352 32772 7404
rect 32824 7352 32830 7404
rect 32950 7352 32956 7404
rect 33008 7352 33014 7404
rect 33042 7352 33048 7404
rect 33100 7392 33106 7404
rect 33628 7395 33655 7426
rect 33689 7404 33701 7429
rect 33778 7420 33784 7472
rect 33836 7460 33842 7472
rect 37660 7460 37688 7500
rect 38397 7497 38409 7500
rect 38443 7528 38455 7531
rect 38443 7500 38516 7528
rect 38443 7497 38455 7500
rect 38397 7491 38455 7497
rect 33836 7432 37688 7460
rect 38197 7463 38255 7469
rect 33836 7420 33842 7432
rect 38197 7429 38209 7463
rect 38243 7429 38255 7463
rect 38197 7423 38255 7429
rect 33689 7395 33692 7404
rect 33628 7392 33692 7395
rect 33100 7364 33692 7392
rect 33100 7352 33106 7364
rect 33686 7352 33692 7364
rect 33744 7352 33750 7404
rect 34330 7352 34336 7404
rect 34388 7392 34394 7404
rect 34517 7395 34575 7401
rect 34517 7392 34529 7395
rect 34388 7364 34529 7392
rect 34388 7352 34394 7364
rect 34517 7361 34529 7364
rect 34563 7361 34575 7395
rect 34517 7355 34575 7361
rect 35161 7395 35219 7401
rect 35161 7361 35173 7395
rect 35207 7392 35219 7395
rect 35342 7392 35348 7404
rect 35207 7364 35348 7392
rect 35207 7361 35219 7364
rect 35161 7355 35219 7361
rect 35342 7352 35348 7364
rect 35400 7352 35406 7404
rect 35986 7352 35992 7404
rect 36044 7392 36050 7404
rect 37461 7395 37519 7401
rect 37461 7392 37473 7395
rect 36044 7364 37473 7392
rect 36044 7352 36050 7364
rect 37461 7361 37473 7364
rect 37507 7361 37519 7395
rect 37461 7355 37519 7361
rect 15562 7324 15568 7336
rect 10980 7296 12388 7324
rect 14476 7296 15568 7324
rect 7116 7265 7144 7296
rect 4801 7259 4859 7265
rect 4801 7225 4813 7259
rect 4847 7225 4859 7259
rect 4801 7219 4859 7225
rect 7101 7259 7159 7265
rect 7101 7225 7113 7259
rect 7147 7225 7159 7259
rect 7101 7219 7159 7225
rect 1949 7191 2007 7197
rect 1949 7157 1961 7191
rect 1995 7188 2007 7191
rect 4246 7188 4252 7200
rect 1995 7160 4252 7188
rect 1995 7157 2007 7160
rect 1949 7151 2007 7157
rect 4246 7148 4252 7160
rect 4304 7148 4310 7200
rect 4982 7148 4988 7200
rect 5040 7188 5046 7200
rect 5442 7188 5448 7200
rect 5040 7160 5448 7188
rect 5040 7148 5046 7160
rect 5442 7148 5448 7160
rect 5500 7148 5506 7200
rect 9861 7191 9919 7197
rect 9861 7157 9873 7191
rect 9907 7188 9919 7191
rect 10962 7188 10968 7200
rect 9907 7160 10968 7188
rect 9907 7157 9919 7160
rect 9861 7151 9919 7157
rect 10962 7148 10968 7160
rect 11020 7148 11026 7200
rect 11054 7148 11060 7200
rect 11112 7148 11118 7200
rect 12894 7148 12900 7200
rect 12952 7188 12958 7200
rect 14476 7188 14504 7296
rect 15562 7284 15568 7296
rect 15620 7284 15626 7336
rect 15654 7284 15660 7336
rect 15712 7284 15718 7336
rect 22186 7284 22192 7336
rect 22244 7324 22250 7336
rect 23109 7327 23167 7333
rect 23109 7324 23121 7327
rect 22244 7296 23121 7324
rect 22244 7284 22250 7296
rect 23109 7293 23121 7296
rect 23155 7293 23167 7327
rect 23109 7287 23167 7293
rect 20898 7216 20904 7268
rect 20956 7256 20962 7268
rect 21269 7259 21327 7265
rect 21269 7256 21281 7259
rect 20956 7228 21281 7256
rect 20956 7216 20962 7228
rect 21269 7225 21281 7228
rect 21315 7256 21327 7259
rect 21818 7256 21824 7268
rect 21315 7228 21824 7256
rect 21315 7225 21327 7228
rect 21269 7219 21327 7225
rect 21818 7216 21824 7228
rect 21876 7216 21882 7268
rect 12952 7160 14504 7188
rect 14645 7191 14703 7197
rect 12952 7148 12958 7160
rect 14645 7157 14657 7191
rect 14691 7188 14703 7191
rect 15010 7188 15016 7200
rect 14691 7160 15016 7188
rect 14691 7157 14703 7160
rect 14645 7151 14703 7157
rect 15010 7148 15016 7160
rect 15068 7148 15074 7200
rect 15102 7148 15108 7200
rect 15160 7148 15166 7200
rect 17313 7191 17371 7197
rect 17313 7157 17325 7191
rect 17359 7188 17371 7191
rect 17954 7188 17960 7200
rect 17359 7160 17960 7188
rect 17359 7157 17371 7160
rect 17313 7151 17371 7157
rect 17954 7148 17960 7160
rect 18012 7148 18018 7200
rect 23124 7188 23152 7287
rect 26234 7284 26240 7336
rect 26292 7284 26298 7336
rect 27154 7284 27160 7336
rect 27212 7284 27218 7336
rect 27433 7327 27491 7333
rect 27433 7293 27445 7327
rect 27479 7324 27491 7327
rect 28718 7324 28724 7336
rect 27479 7296 28724 7324
rect 27479 7293 27491 7296
rect 27433 7287 27491 7293
rect 28718 7284 28724 7296
rect 28776 7284 28782 7336
rect 31297 7327 31355 7333
rect 31297 7293 31309 7327
rect 31343 7324 31355 7327
rect 31570 7324 31576 7336
rect 31343 7296 31576 7324
rect 31343 7293 31355 7296
rect 31297 7287 31355 7293
rect 31570 7284 31576 7296
rect 31628 7324 31634 7336
rect 32398 7324 32404 7336
rect 31628 7296 32404 7324
rect 31628 7284 31634 7296
rect 32398 7284 32404 7296
rect 32456 7284 32462 7336
rect 35250 7284 35256 7336
rect 35308 7324 35314 7336
rect 35437 7327 35495 7333
rect 35437 7324 35449 7327
rect 35308 7296 35449 7324
rect 35308 7284 35314 7296
rect 35437 7293 35449 7296
rect 35483 7324 35495 7327
rect 35618 7324 35624 7336
rect 35483 7296 35624 7324
rect 35483 7293 35495 7296
rect 35437 7287 35495 7293
rect 35618 7284 35624 7296
rect 35676 7284 35682 7336
rect 36262 7284 36268 7336
rect 36320 7284 36326 7336
rect 36357 7327 36415 7333
rect 36357 7293 36369 7327
rect 36403 7293 36415 7327
rect 36357 7287 36415 7293
rect 36474 7327 36532 7333
rect 36474 7293 36486 7327
rect 36520 7324 36532 7327
rect 36722 7324 36728 7336
rect 36520 7296 36728 7324
rect 36520 7293 36532 7296
rect 36474 7287 36532 7293
rect 31846 7216 31852 7268
rect 31904 7256 31910 7268
rect 32582 7256 32588 7268
rect 31904 7228 32588 7256
rect 31904 7216 31910 7228
rect 32582 7216 32588 7228
rect 32640 7216 32646 7268
rect 34238 7216 34244 7268
rect 34296 7256 34302 7268
rect 34977 7259 35035 7265
rect 34977 7256 34989 7259
rect 34296 7228 34989 7256
rect 34296 7216 34302 7228
rect 34977 7225 34989 7228
rect 35023 7225 35035 7259
rect 34977 7219 35035 7225
rect 35066 7216 35072 7268
rect 35124 7256 35130 7268
rect 35345 7259 35403 7265
rect 35345 7256 35357 7259
rect 35124 7228 35357 7256
rect 35124 7216 35130 7228
rect 35345 7225 35357 7228
rect 35391 7225 35403 7259
rect 36372 7256 36400 7287
rect 36722 7284 36728 7296
rect 36780 7284 36786 7336
rect 37182 7284 37188 7336
rect 37240 7324 37246 7336
rect 38212 7324 38240 7423
rect 38488 7392 38516 7500
rect 38562 7488 38568 7540
rect 38620 7488 38626 7540
rect 39209 7531 39267 7537
rect 39209 7497 39221 7531
rect 39255 7528 39267 7531
rect 39298 7528 39304 7540
rect 39255 7500 39304 7528
rect 39255 7497 39267 7500
rect 39209 7491 39267 7497
rect 39298 7488 39304 7500
rect 39356 7488 39362 7540
rect 39574 7488 39580 7540
rect 39632 7528 39638 7540
rect 40681 7531 40739 7537
rect 40681 7528 40693 7531
rect 39632 7500 40693 7528
rect 39632 7488 39638 7500
rect 40681 7497 40693 7500
rect 40727 7497 40739 7531
rect 40681 7491 40739 7497
rect 41414 7488 41420 7540
rect 41472 7488 41478 7540
rect 40313 7463 40371 7469
rect 40313 7429 40325 7463
rect 40359 7460 40371 7463
rect 40359 7432 42656 7460
rect 40359 7429 40371 7432
rect 40313 7423 40371 7429
rect 39853 7395 39911 7401
rect 39853 7392 39865 7395
rect 38488 7364 39865 7392
rect 39853 7361 39865 7364
rect 39899 7392 39911 7395
rect 40957 7395 41015 7401
rect 40957 7392 40969 7395
rect 39899 7390 40448 7392
rect 40604 7390 40969 7392
rect 39899 7364 40969 7390
rect 39899 7361 39911 7364
rect 40420 7362 40632 7364
rect 39853 7355 39911 7361
rect 40957 7361 40969 7364
rect 41003 7361 41015 7395
rect 40957 7355 41015 7361
rect 41598 7352 41604 7404
rect 41656 7352 41662 7404
rect 42628 7401 42656 7432
rect 42613 7395 42671 7401
rect 42613 7361 42625 7395
rect 42659 7361 42671 7395
rect 42613 7355 42671 7361
rect 42797 7395 42855 7401
rect 42797 7361 42809 7395
rect 42843 7361 42855 7395
rect 42797 7355 42855 7361
rect 39390 7324 39396 7336
rect 37240 7296 39396 7324
rect 37240 7284 37246 7296
rect 39390 7284 39396 7296
rect 39448 7284 39454 7336
rect 39485 7327 39543 7333
rect 39485 7293 39497 7327
rect 39531 7293 39543 7327
rect 39485 7287 39543 7293
rect 39500 7256 39528 7287
rect 39758 7284 39764 7336
rect 39816 7284 39822 7336
rect 40497 7327 40555 7333
rect 40497 7293 40509 7327
rect 40543 7293 40555 7327
rect 40497 7287 40555 7293
rect 40589 7327 40647 7333
rect 40589 7293 40601 7327
rect 40635 7324 40647 7327
rect 40770 7324 40776 7336
rect 40635 7296 40776 7324
rect 40635 7293 40647 7296
rect 40589 7287 40647 7293
rect 40218 7256 40224 7268
rect 36372 7228 40224 7256
rect 35345 7219 35403 7225
rect 23382 7188 23388 7200
rect 23124 7160 23388 7188
rect 23382 7148 23388 7160
rect 23440 7148 23446 7200
rect 24394 7148 24400 7200
rect 24452 7188 24458 7200
rect 24489 7191 24547 7197
rect 24489 7188 24501 7191
rect 24452 7160 24501 7188
rect 24452 7148 24458 7160
rect 24489 7157 24501 7160
rect 24535 7157 24547 7191
rect 24489 7151 24547 7157
rect 27614 7148 27620 7200
rect 27672 7188 27678 7200
rect 29733 7191 29791 7197
rect 29733 7188 29745 7191
rect 27672 7160 29745 7188
rect 27672 7148 27678 7160
rect 29733 7157 29745 7160
rect 29779 7157 29791 7191
rect 29733 7151 29791 7157
rect 30377 7191 30435 7197
rect 30377 7157 30389 7191
rect 30423 7188 30435 7191
rect 30650 7188 30656 7200
rect 30423 7160 30656 7188
rect 30423 7157 30435 7160
rect 30377 7151 30435 7157
rect 30650 7148 30656 7160
rect 30708 7148 30714 7200
rect 31478 7148 31484 7200
rect 31536 7188 31542 7200
rect 32030 7188 32036 7200
rect 31536 7160 32036 7188
rect 31536 7148 31542 7160
rect 32030 7148 32036 7160
rect 32088 7148 32094 7200
rect 32306 7148 32312 7200
rect 32364 7148 32370 7200
rect 32398 7148 32404 7200
rect 32456 7188 32462 7200
rect 33597 7191 33655 7197
rect 33597 7188 33609 7191
rect 32456 7160 33609 7188
rect 32456 7148 32462 7160
rect 33597 7157 33609 7160
rect 33643 7157 33655 7191
rect 33597 7151 33655 7157
rect 33778 7148 33784 7200
rect 33836 7148 33842 7200
rect 34333 7191 34391 7197
rect 34333 7157 34345 7191
rect 34379 7188 34391 7191
rect 34790 7188 34796 7200
rect 34379 7160 34796 7188
rect 34379 7157 34391 7160
rect 34333 7151 34391 7157
rect 34790 7148 34796 7160
rect 34848 7148 34854 7200
rect 36630 7148 36636 7200
rect 36688 7148 36694 7200
rect 38396 7197 38424 7228
rect 40218 7216 40224 7228
rect 40276 7216 40282 7268
rect 40310 7216 40316 7268
rect 40368 7256 40374 7268
rect 40512 7256 40540 7287
rect 40770 7284 40776 7296
rect 40828 7284 40834 7336
rect 40862 7284 40868 7336
rect 40920 7284 40926 7336
rect 41414 7284 41420 7336
rect 41472 7324 41478 7336
rect 42812 7324 42840 7355
rect 41472 7296 42840 7324
rect 41472 7284 41478 7296
rect 40368 7228 40540 7256
rect 40368 7216 40374 7228
rect 38381 7191 38439 7197
rect 38381 7157 38393 7191
rect 38427 7157 38439 7191
rect 38381 7151 38439 7157
rect 40126 7148 40132 7200
rect 40184 7188 40190 7200
rect 42613 7191 42671 7197
rect 42613 7188 42625 7191
rect 40184 7160 42625 7188
rect 40184 7148 40190 7160
rect 42613 7157 42625 7160
rect 42659 7157 42671 7191
rect 42613 7151 42671 7157
rect 1104 7098 44896 7120
rect 1104 7046 6423 7098
rect 6475 7046 6487 7098
rect 6539 7046 6551 7098
rect 6603 7046 6615 7098
rect 6667 7046 6679 7098
rect 6731 7046 17370 7098
rect 17422 7046 17434 7098
rect 17486 7046 17498 7098
rect 17550 7046 17562 7098
rect 17614 7046 17626 7098
rect 17678 7046 28317 7098
rect 28369 7046 28381 7098
rect 28433 7046 28445 7098
rect 28497 7046 28509 7098
rect 28561 7046 28573 7098
rect 28625 7046 39264 7098
rect 39316 7046 39328 7098
rect 39380 7046 39392 7098
rect 39444 7046 39456 7098
rect 39508 7046 39520 7098
rect 39572 7046 44896 7098
rect 1104 7024 44896 7046
rect 3142 6944 3148 6996
rect 3200 6984 3206 6996
rect 3421 6987 3479 6993
rect 3421 6984 3433 6987
rect 3200 6956 3433 6984
rect 3200 6944 3206 6956
rect 3421 6953 3433 6956
rect 3467 6953 3479 6987
rect 3421 6947 3479 6953
rect 9388 6987 9446 6993
rect 9388 6953 9400 6987
rect 9434 6984 9446 6987
rect 10134 6984 10140 6996
rect 9434 6956 10140 6984
rect 9434 6953 9446 6956
rect 9388 6947 9446 6953
rect 10134 6944 10140 6956
rect 10192 6944 10198 6996
rect 10594 6944 10600 6996
rect 10652 6984 10658 6996
rect 11790 6984 11796 6996
rect 10652 6956 11796 6984
rect 10652 6944 10658 6956
rect 11790 6944 11796 6956
rect 11848 6944 11854 6996
rect 12345 6987 12403 6993
rect 12345 6953 12357 6987
rect 12391 6984 12403 6987
rect 13354 6984 13360 6996
rect 12391 6956 13360 6984
rect 12391 6953 12403 6956
rect 12345 6947 12403 6953
rect 13354 6944 13360 6956
rect 13412 6944 13418 6996
rect 15654 6984 15660 6996
rect 15304 6956 15660 6984
rect 12989 6919 13047 6925
rect 12989 6885 13001 6919
rect 13035 6885 13047 6919
rect 15304 6916 15332 6956
rect 15654 6944 15660 6956
rect 15712 6984 15718 6996
rect 20990 6984 20996 6996
rect 15712 6956 17632 6984
rect 15712 6944 15718 6956
rect 12989 6879 13047 6885
rect 14844 6888 15332 6916
rect 6914 6808 6920 6860
rect 6972 6848 6978 6860
rect 9125 6851 9183 6857
rect 9125 6848 9137 6851
rect 6972 6820 9137 6848
rect 6972 6808 6978 6820
rect 9125 6817 9137 6820
rect 9171 6848 9183 6851
rect 9398 6848 9404 6860
rect 9171 6820 9404 6848
rect 9171 6817 9183 6820
rect 9125 6811 9183 6817
rect 9398 6808 9404 6820
rect 9456 6848 9462 6860
rect 10594 6848 10600 6860
rect 9456 6820 10600 6848
rect 9456 6808 9462 6820
rect 10594 6808 10600 6820
rect 10652 6808 10658 6860
rect 2041 6783 2099 6789
rect 2041 6749 2053 6783
rect 2087 6780 2099 6783
rect 3878 6780 3884 6792
rect 2087 6752 3884 6780
rect 2087 6749 2099 6752
rect 2041 6743 2099 6749
rect 3878 6740 3884 6752
rect 3936 6780 3942 6792
rect 3973 6783 4031 6789
rect 3973 6780 3985 6783
rect 3936 6752 3985 6780
rect 3936 6740 3942 6752
rect 3973 6749 3985 6752
rect 4019 6749 4031 6783
rect 3973 6743 4031 6749
rect 4240 6783 4298 6789
rect 4240 6749 4252 6783
rect 4286 6780 4298 6783
rect 5350 6780 5356 6792
rect 4286 6752 5356 6780
rect 4286 6749 4298 6752
rect 4240 6743 4298 6749
rect 5350 6740 5356 6752
rect 5408 6740 5414 6792
rect 6178 6740 6184 6792
rect 6236 6780 6242 6792
rect 6549 6783 6607 6789
rect 6549 6780 6561 6783
rect 6236 6752 6561 6780
rect 6236 6740 6242 6752
rect 6549 6749 6561 6752
rect 6595 6749 6607 6783
rect 6549 6743 6607 6749
rect 7558 6740 7564 6792
rect 7616 6780 7622 6792
rect 8297 6783 8355 6789
rect 8297 6780 8309 6783
rect 7616 6752 8309 6780
rect 7616 6740 7622 6752
rect 8297 6749 8309 6752
rect 8343 6749 8355 6783
rect 8297 6743 8355 6749
rect 11054 6740 11060 6792
rect 11112 6780 11118 6792
rect 11885 6783 11943 6789
rect 11885 6780 11897 6783
rect 11112 6752 11897 6780
rect 11112 6740 11118 6752
rect 11885 6749 11897 6752
rect 11931 6749 11943 6783
rect 11885 6743 11943 6749
rect 12529 6783 12587 6789
rect 12529 6749 12541 6783
rect 12575 6780 12587 6783
rect 13004 6780 13032 6879
rect 13446 6808 13452 6860
rect 13504 6808 13510 6860
rect 13633 6851 13691 6857
rect 13633 6817 13645 6851
rect 13679 6848 13691 6851
rect 14844 6848 14872 6888
rect 13679 6820 14872 6848
rect 13679 6817 13691 6820
rect 13633 6811 13691 6817
rect 14918 6808 14924 6860
rect 14976 6848 14982 6860
rect 15289 6851 15347 6857
rect 15289 6848 15301 6851
rect 14976 6820 15301 6848
rect 14976 6808 14982 6820
rect 15289 6817 15301 6820
rect 15335 6817 15347 6851
rect 17604 6848 17632 6956
rect 20456 6956 20996 6984
rect 20456 6928 20484 6956
rect 20990 6944 20996 6956
rect 21048 6984 21054 6996
rect 21450 6984 21456 6996
rect 21048 6956 21456 6984
rect 21048 6944 21054 6956
rect 21450 6944 21456 6956
rect 21508 6944 21514 6996
rect 31573 6987 31631 6993
rect 31573 6953 31585 6987
rect 31619 6984 31631 6987
rect 32766 6984 32772 6996
rect 31619 6956 32772 6984
rect 31619 6953 31631 6956
rect 31573 6947 31631 6953
rect 32766 6944 32772 6956
rect 32824 6944 32830 6996
rect 35713 6987 35771 6993
rect 35713 6953 35725 6987
rect 35759 6984 35771 6987
rect 36998 6984 37004 6996
rect 35759 6956 37004 6984
rect 35759 6953 35771 6956
rect 35713 6947 35771 6953
rect 36998 6944 37004 6956
rect 37056 6944 37062 6996
rect 40218 6944 40224 6996
rect 40276 6984 40282 6996
rect 40770 6984 40776 6996
rect 40276 6956 40776 6984
rect 40276 6944 40282 6956
rect 40770 6944 40776 6956
rect 40828 6984 40834 6996
rect 40828 6956 41000 6984
rect 40828 6944 40834 6956
rect 20438 6916 20444 6928
rect 19306 6888 20444 6916
rect 17681 6851 17739 6857
rect 17681 6848 17693 6851
rect 17604 6820 17693 6848
rect 15289 6811 15347 6817
rect 17681 6817 17693 6820
rect 17727 6817 17739 6851
rect 17681 6811 17739 6817
rect 18598 6808 18604 6860
rect 18656 6808 18662 6860
rect 19306 6848 19334 6888
rect 20438 6876 20444 6888
rect 20496 6876 20502 6928
rect 20898 6916 20904 6928
rect 20548 6888 20904 6916
rect 20548 6857 20576 6888
rect 20898 6876 20904 6888
rect 20956 6876 20962 6928
rect 21266 6876 21272 6928
rect 21324 6916 21330 6928
rect 21634 6916 21640 6928
rect 21324 6888 21640 6916
rect 21324 6876 21330 6888
rect 21634 6876 21640 6888
rect 21692 6876 21698 6928
rect 32398 6916 32404 6928
rect 31864 6888 32404 6916
rect 18800 6820 19334 6848
rect 20533 6851 20591 6857
rect 12575 6752 13032 6780
rect 13357 6783 13415 6789
rect 12575 6749 12587 6752
rect 12529 6743 12587 6749
rect 13357 6749 13369 6783
rect 13403 6780 13415 6783
rect 14461 6783 14519 6789
rect 13403 6752 14412 6780
rect 13403 6749 13415 6752
rect 13357 6743 13415 6749
rect 2308 6715 2366 6721
rect 2308 6681 2320 6715
rect 2354 6712 2366 6715
rect 4430 6712 4436 6724
rect 2354 6684 4436 6712
rect 2354 6681 2366 6684
rect 2308 6675 2366 6681
rect 4430 6672 4436 6684
rect 4488 6712 4494 6724
rect 10686 6712 10692 6724
rect 4488 6684 5396 6712
rect 10626 6684 10692 6712
rect 4488 6672 4494 6684
rect 5368 6653 5396 6684
rect 10686 6672 10692 6684
rect 10744 6672 10750 6724
rect 14182 6712 14188 6724
rect 10796 6684 14188 6712
rect 5353 6647 5411 6653
rect 5353 6613 5365 6647
rect 5399 6613 5411 6647
rect 5353 6607 5411 6613
rect 6365 6647 6423 6653
rect 6365 6613 6377 6647
rect 6411 6644 6423 6647
rect 6822 6644 6828 6656
rect 6411 6616 6828 6644
rect 6411 6613 6423 6616
rect 6365 6607 6423 6613
rect 6822 6604 6828 6616
rect 6880 6604 6886 6656
rect 8481 6647 8539 6653
rect 8481 6613 8493 6647
rect 8527 6644 8539 6647
rect 10796 6644 10824 6684
rect 14182 6672 14188 6684
rect 14240 6672 14246 6724
rect 14384 6712 14412 6752
rect 14461 6749 14473 6783
rect 14507 6780 14519 6783
rect 15102 6780 15108 6792
rect 14507 6752 15108 6780
rect 14507 6749 14519 6752
rect 14461 6743 14519 6749
rect 15102 6740 15108 6752
rect 15160 6740 15166 6792
rect 18506 6740 18512 6792
rect 18564 6740 18570 6792
rect 15010 6712 15016 6724
rect 14384 6684 15016 6712
rect 15010 6672 15016 6684
rect 15068 6672 15074 6724
rect 15562 6721 15568 6724
rect 15556 6675 15568 6721
rect 15562 6672 15568 6675
rect 15620 6672 15626 6724
rect 17497 6715 17555 6721
rect 17497 6712 17509 6715
rect 16684 6684 17509 6712
rect 8527 6616 10824 6644
rect 8527 6613 8539 6616
rect 8481 6607 8539 6613
rect 10870 6604 10876 6656
rect 10928 6604 10934 6656
rect 11606 6604 11612 6656
rect 11664 6644 11670 6656
rect 11701 6647 11759 6653
rect 11701 6644 11713 6647
rect 11664 6616 11713 6644
rect 11664 6604 11670 6616
rect 11701 6613 11713 6616
rect 11747 6613 11759 6647
rect 11701 6607 11759 6613
rect 14277 6647 14335 6653
rect 14277 6613 14289 6647
rect 14323 6644 14335 6647
rect 14550 6644 14556 6656
rect 14323 6616 14556 6644
rect 14323 6613 14335 6616
rect 14277 6607 14335 6613
rect 14550 6604 14556 6616
rect 14608 6604 14614 6656
rect 16684 6653 16712 6684
rect 17497 6681 17509 6684
rect 17543 6712 17555 6715
rect 17770 6712 17776 6724
rect 17543 6684 17776 6712
rect 17543 6681 17555 6684
rect 17497 6675 17555 6681
rect 17770 6672 17776 6684
rect 17828 6672 17834 6724
rect 18138 6672 18144 6724
rect 18196 6712 18202 6724
rect 18800 6712 18828 6820
rect 20533 6817 20545 6851
rect 20579 6817 20591 6851
rect 21284 6848 21312 6876
rect 20533 6811 20591 6817
rect 20640 6820 21312 6848
rect 21376 6820 22094 6848
rect 20165 6783 20223 6789
rect 20165 6780 20177 6783
rect 18196 6684 18828 6712
rect 18892 6752 20177 6780
rect 18196 6672 18202 6684
rect 16669 6647 16727 6653
rect 16669 6613 16681 6647
rect 16715 6613 16727 6647
rect 16669 6607 16727 6613
rect 17126 6604 17132 6656
rect 17184 6604 17190 6656
rect 17218 6604 17224 6656
rect 17276 6644 17282 6656
rect 17589 6647 17647 6653
rect 17589 6644 17601 6647
rect 17276 6616 17601 6644
rect 17276 6604 17282 6616
rect 17589 6613 17601 6616
rect 17635 6644 17647 6647
rect 17862 6644 17868 6656
rect 17635 6616 17868 6644
rect 17635 6613 17647 6616
rect 17589 6607 17647 6613
rect 17862 6604 17868 6616
rect 17920 6604 17926 6656
rect 18892 6653 18920 6752
rect 20165 6749 20177 6752
rect 20211 6749 20223 6783
rect 20165 6743 20223 6749
rect 20349 6783 20407 6789
rect 20349 6749 20361 6783
rect 20395 6749 20407 6783
rect 20349 6743 20407 6749
rect 20364 6712 20392 6743
rect 20438 6740 20444 6792
rect 20496 6780 20502 6792
rect 20496 6752 20541 6780
rect 20496 6740 20502 6752
rect 20640 6712 20668 6820
rect 21376 6789 21404 6820
rect 20717 6783 20775 6789
rect 20717 6749 20729 6783
rect 20763 6749 20775 6783
rect 20717 6743 20775 6749
rect 21361 6783 21419 6789
rect 21361 6749 21373 6783
rect 21407 6749 21419 6783
rect 21361 6743 21419 6749
rect 20364 6684 20668 6712
rect 20732 6712 20760 6743
rect 21450 6740 21456 6792
rect 21508 6780 21514 6792
rect 21508 6752 21553 6780
rect 21508 6740 21514 6752
rect 21634 6740 21640 6792
rect 21692 6740 21698 6792
rect 21818 6740 21824 6792
rect 21876 6789 21882 6792
rect 21876 6780 21884 6789
rect 21876 6752 21921 6780
rect 21876 6743 21884 6752
rect 21876 6740 21882 6743
rect 21726 6712 21732 6724
rect 20732 6684 21732 6712
rect 21726 6672 21732 6684
rect 21784 6672 21790 6724
rect 22066 6712 22094 6820
rect 23750 6808 23756 6860
rect 23808 6808 23814 6860
rect 23842 6808 23848 6860
rect 23900 6808 23906 6860
rect 24673 6851 24731 6857
rect 24673 6817 24685 6851
rect 24719 6817 24731 6851
rect 24673 6811 24731 6817
rect 25133 6851 25191 6857
rect 25133 6817 25145 6851
rect 25179 6817 25191 6851
rect 27614 6848 27620 6860
rect 25133 6811 25191 6817
rect 26804 6820 27620 6848
rect 23661 6783 23719 6789
rect 23661 6749 23673 6783
rect 23707 6780 23719 6783
rect 24394 6780 24400 6792
rect 23707 6752 24400 6780
rect 23707 6749 23719 6752
rect 23661 6743 23719 6749
rect 24394 6740 24400 6752
rect 24452 6780 24458 6792
rect 24688 6780 24716 6811
rect 24452 6752 24716 6780
rect 24765 6783 24823 6789
rect 24452 6740 24458 6752
rect 24765 6749 24777 6783
rect 24811 6780 24823 6783
rect 25038 6780 25044 6792
rect 24811 6752 25044 6780
rect 24811 6749 24823 6752
rect 24765 6743 24823 6749
rect 25038 6740 25044 6752
rect 25096 6740 25102 6792
rect 25148 6712 25176 6811
rect 25961 6783 26019 6789
rect 25961 6749 25973 6783
rect 26007 6780 26019 6783
rect 26050 6780 26056 6792
rect 26007 6752 26056 6780
rect 26007 6749 26019 6752
rect 25961 6743 26019 6749
rect 26050 6740 26056 6752
rect 26108 6740 26114 6792
rect 26804 6789 26832 6820
rect 27614 6808 27620 6820
rect 27672 6808 27678 6860
rect 31864 6857 31892 6888
rect 32398 6876 32404 6888
rect 32456 6876 32462 6928
rect 32582 6876 32588 6928
rect 32640 6916 32646 6928
rect 39758 6916 39764 6928
rect 32640 6888 39764 6916
rect 32640 6876 32646 6888
rect 31849 6851 31907 6857
rect 31849 6817 31861 6851
rect 31895 6817 31907 6851
rect 31849 6811 31907 6817
rect 32214 6808 32220 6860
rect 32272 6848 32278 6860
rect 33042 6848 33048 6860
rect 32272 6820 33048 6848
rect 32272 6808 32278 6820
rect 33042 6808 33048 6820
rect 33100 6808 33106 6860
rect 26789 6783 26847 6789
rect 26789 6749 26801 6783
rect 26835 6749 26847 6783
rect 26789 6743 26847 6749
rect 27246 6740 27252 6792
rect 27304 6740 27310 6792
rect 29730 6740 29736 6792
rect 29788 6740 29794 6792
rect 31757 6783 31815 6789
rect 31757 6749 31769 6783
rect 31803 6749 31815 6783
rect 31757 6743 31815 6749
rect 32125 6783 32183 6789
rect 32125 6749 32137 6783
rect 32171 6780 32183 6783
rect 32582 6780 32588 6792
rect 32171 6752 32588 6780
rect 32171 6749 32183 6752
rect 32125 6743 32183 6749
rect 22066 6684 25176 6712
rect 28445 6715 28503 6721
rect 28445 6681 28457 6715
rect 28491 6712 28503 6715
rect 28718 6712 28724 6724
rect 28491 6684 28724 6712
rect 28491 6681 28503 6684
rect 28445 6675 28503 6681
rect 28718 6672 28724 6684
rect 28776 6672 28782 6724
rect 30000 6715 30058 6721
rect 30000 6681 30012 6715
rect 30046 6712 30058 6715
rect 31018 6712 31024 6724
rect 30046 6684 31024 6712
rect 30046 6681 30058 6684
rect 30000 6675 30058 6681
rect 31018 6672 31024 6684
rect 31076 6672 31082 6724
rect 31772 6712 31800 6743
rect 32582 6740 32588 6752
rect 32640 6740 32646 6792
rect 32677 6783 32735 6789
rect 32677 6749 32689 6783
rect 32723 6780 32735 6783
rect 33778 6780 33784 6792
rect 32723 6752 33784 6780
rect 32723 6749 32735 6752
rect 32677 6743 32735 6749
rect 33778 6740 33784 6752
rect 33836 6740 33842 6792
rect 34164 6789 34192 6888
rect 39758 6876 39764 6888
rect 39816 6916 39822 6928
rect 40862 6916 40868 6928
rect 39816 6888 40868 6916
rect 39816 6876 39822 6888
rect 40862 6876 40868 6888
rect 40920 6876 40926 6928
rect 35158 6808 35164 6860
rect 35216 6848 35222 6860
rect 40402 6848 40408 6860
rect 35216 6820 40408 6848
rect 35216 6808 35222 6820
rect 40402 6808 40408 6820
rect 40460 6848 40466 6860
rect 40972 6848 41000 6956
rect 40460 6820 40816 6848
rect 40972 6820 41460 6848
rect 40460 6808 40466 6820
rect 40788 6792 40816 6820
rect 33965 6783 34023 6789
rect 33965 6749 33977 6783
rect 34011 6749 34023 6783
rect 33965 6743 34023 6749
rect 34149 6783 34207 6789
rect 34149 6749 34161 6783
rect 34195 6749 34207 6783
rect 34149 6743 34207 6749
rect 31938 6712 31944 6724
rect 31128 6684 31944 6712
rect 18877 6647 18935 6653
rect 18877 6613 18889 6647
rect 18923 6613 18935 6647
rect 18877 6607 18935 6613
rect 20714 6604 20720 6656
rect 20772 6644 20778 6656
rect 20901 6647 20959 6653
rect 20901 6644 20913 6647
rect 20772 6616 20913 6644
rect 20772 6604 20778 6616
rect 20901 6613 20913 6616
rect 20947 6613 20959 6647
rect 20901 6607 20959 6613
rect 22002 6604 22008 6656
rect 22060 6604 22066 6656
rect 23293 6647 23351 6653
rect 23293 6613 23305 6647
rect 23339 6644 23351 6647
rect 23566 6644 23572 6656
rect 23339 6616 23572 6644
rect 23339 6613 23351 6616
rect 23293 6607 23351 6613
rect 23566 6604 23572 6616
rect 23624 6604 23630 6656
rect 25777 6647 25835 6653
rect 25777 6613 25789 6647
rect 25823 6644 25835 6647
rect 25866 6644 25872 6656
rect 25823 6616 25872 6644
rect 25823 6613 25835 6616
rect 25777 6607 25835 6613
rect 25866 6604 25872 6616
rect 25924 6604 25930 6656
rect 26605 6647 26663 6653
rect 26605 6613 26617 6647
rect 26651 6644 26663 6647
rect 27890 6644 27896 6656
rect 26651 6616 27896 6644
rect 26651 6613 26663 6616
rect 26605 6607 26663 6613
rect 27890 6604 27896 6616
rect 27948 6604 27954 6656
rect 30374 6604 30380 6656
rect 30432 6644 30438 6656
rect 31128 6653 31156 6684
rect 31938 6672 31944 6684
rect 31996 6672 32002 6724
rect 33980 6712 34008 6743
rect 34882 6740 34888 6792
rect 34940 6780 34946 6792
rect 35345 6783 35403 6789
rect 35345 6780 35357 6783
rect 34940 6752 35357 6780
rect 34940 6740 34946 6752
rect 35345 6749 35357 6752
rect 35391 6749 35403 6783
rect 35345 6743 35403 6749
rect 35713 6783 35771 6789
rect 35713 6749 35725 6783
rect 35759 6749 35771 6783
rect 35713 6743 35771 6749
rect 35526 6712 35532 6724
rect 32140 6684 34008 6712
rect 34072 6684 35532 6712
rect 31113 6647 31171 6653
rect 31113 6644 31125 6647
rect 30432 6616 31125 6644
rect 30432 6604 30438 6616
rect 31113 6613 31125 6616
rect 31159 6613 31171 6647
rect 31113 6607 31171 6613
rect 32030 6604 32036 6656
rect 32088 6644 32094 6656
rect 32140 6644 32168 6684
rect 32088 6616 32168 6644
rect 32088 6604 32094 6616
rect 32674 6604 32680 6656
rect 32732 6644 32738 6656
rect 32769 6647 32827 6653
rect 32769 6644 32781 6647
rect 32732 6616 32781 6644
rect 32732 6604 32738 6616
rect 32769 6613 32781 6616
rect 32815 6644 32827 6647
rect 34072 6644 34100 6684
rect 35526 6672 35532 6684
rect 35584 6672 35590 6724
rect 35728 6712 35756 6743
rect 35802 6740 35808 6792
rect 35860 6780 35866 6792
rect 35860 6752 36492 6780
rect 35860 6740 35866 6752
rect 35986 6712 35992 6724
rect 35728 6684 35992 6712
rect 35986 6672 35992 6684
rect 36044 6712 36050 6724
rect 36354 6712 36360 6724
rect 36044 6684 36360 6712
rect 36044 6672 36050 6684
rect 36354 6672 36360 6684
rect 36412 6672 36418 6724
rect 32815 6616 34100 6644
rect 32815 6613 32827 6616
rect 32769 6607 32827 6613
rect 34146 6604 34152 6656
rect 34204 6644 34210 6656
rect 34333 6647 34391 6653
rect 34333 6644 34345 6647
rect 34204 6616 34345 6644
rect 34204 6604 34210 6616
rect 34333 6613 34345 6616
rect 34379 6613 34391 6647
rect 34333 6607 34391 6613
rect 35342 6604 35348 6656
rect 35400 6644 35406 6656
rect 35897 6647 35955 6653
rect 35897 6644 35909 6647
rect 35400 6616 35909 6644
rect 35400 6604 35406 6616
rect 35897 6613 35909 6616
rect 35943 6644 35955 6647
rect 36262 6644 36268 6656
rect 35943 6616 36268 6644
rect 35943 6613 35955 6616
rect 35897 6607 35955 6613
rect 36262 6604 36268 6616
rect 36320 6604 36326 6656
rect 36464 6644 36492 6752
rect 36538 6740 36544 6792
rect 36596 6740 36602 6792
rect 36630 6740 36636 6792
rect 36688 6780 36694 6792
rect 36725 6783 36783 6789
rect 36725 6780 36737 6783
rect 36688 6752 36737 6780
rect 36688 6740 36694 6752
rect 36725 6749 36737 6752
rect 36771 6749 36783 6783
rect 36725 6743 36783 6749
rect 36906 6740 36912 6792
rect 36964 6740 36970 6792
rect 37369 6783 37427 6789
rect 37369 6749 37381 6783
rect 37415 6749 37427 6783
rect 37369 6743 37427 6749
rect 39485 6783 39543 6789
rect 39485 6749 39497 6783
rect 39531 6780 39543 6783
rect 40126 6780 40132 6792
rect 39531 6752 40132 6780
rect 39531 6749 39543 6752
rect 39485 6743 39543 6749
rect 36556 6712 36584 6740
rect 37384 6712 37412 6743
rect 40126 6740 40132 6752
rect 40184 6740 40190 6792
rect 40218 6740 40224 6792
rect 40276 6740 40282 6792
rect 40494 6740 40500 6792
rect 40552 6740 40558 6792
rect 40678 6740 40684 6792
rect 40736 6740 40742 6792
rect 40770 6740 40776 6792
rect 40828 6780 40834 6792
rect 41325 6783 41383 6789
rect 41325 6780 41337 6783
rect 40828 6752 41337 6780
rect 40828 6740 40834 6752
rect 41325 6749 41337 6752
rect 41371 6749 41383 6783
rect 41432 6780 41460 6820
rect 43438 6808 43444 6860
rect 43496 6808 43502 6860
rect 43349 6783 43407 6789
rect 41432 6752 42748 6780
rect 41325 6743 41383 6749
rect 41570 6715 41628 6721
rect 41570 6712 41582 6715
rect 36556 6684 37412 6712
rect 39316 6684 41582 6712
rect 36633 6647 36691 6653
rect 36633 6644 36645 6647
rect 36464 6616 36645 6644
rect 36633 6613 36645 6616
rect 36679 6644 36691 6647
rect 37366 6644 37372 6656
rect 36679 6616 37372 6644
rect 36679 6613 36691 6616
rect 36633 6607 36691 6613
rect 37366 6604 37372 6616
rect 37424 6604 37430 6656
rect 37461 6647 37519 6653
rect 37461 6613 37473 6647
rect 37507 6644 37519 6647
rect 37642 6644 37648 6656
rect 37507 6616 37648 6644
rect 37507 6613 37519 6616
rect 37461 6607 37519 6613
rect 37642 6604 37648 6616
rect 37700 6604 37706 6656
rect 39316 6653 39344 6684
rect 41570 6681 41582 6684
rect 41616 6681 41628 6715
rect 41570 6675 41628 6681
rect 39301 6647 39359 6653
rect 39301 6613 39313 6647
rect 39347 6613 39359 6647
rect 39301 6607 39359 6613
rect 40037 6647 40095 6653
rect 40037 6613 40049 6647
rect 40083 6644 40095 6647
rect 41414 6644 41420 6656
rect 40083 6616 41420 6644
rect 40083 6613 40095 6616
rect 40037 6607 40095 6613
rect 41414 6604 41420 6616
rect 41472 6604 41478 6656
rect 42720 6653 42748 6752
rect 43349 6749 43361 6783
rect 43395 6749 43407 6783
rect 43349 6743 43407 6749
rect 42705 6647 42763 6653
rect 42705 6613 42717 6647
rect 42751 6644 42763 6647
rect 43364 6644 43392 6743
rect 42751 6616 43392 6644
rect 42751 6613 42763 6616
rect 42705 6607 42763 6613
rect 43714 6604 43720 6656
rect 43772 6604 43778 6656
rect 1104 6554 45051 6576
rect 1104 6502 11896 6554
rect 11948 6502 11960 6554
rect 12012 6502 12024 6554
rect 12076 6502 12088 6554
rect 12140 6502 12152 6554
rect 12204 6502 22843 6554
rect 22895 6502 22907 6554
rect 22959 6502 22971 6554
rect 23023 6502 23035 6554
rect 23087 6502 23099 6554
rect 23151 6502 33790 6554
rect 33842 6502 33854 6554
rect 33906 6502 33918 6554
rect 33970 6502 33982 6554
rect 34034 6502 34046 6554
rect 34098 6502 44737 6554
rect 44789 6502 44801 6554
rect 44853 6502 44865 6554
rect 44917 6502 44929 6554
rect 44981 6502 44993 6554
rect 45045 6502 45051 6554
rect 1104 6480 45051 6502
rect 3421 6443 3479 6449
rect 3421 6409 3433 6443
rect 3467 6440 3479 6443
rect 4338 6440 4344 6452
rect 3467 6412 4344 6440
rect 3467 6409 3479 6412
rect 3421 6403 3479 6409
rect 4338 6400 4344 6412
rect 4396 6400 4402 6452
rect 5166 6400 5172 6452
rect 5224 6440 5230 6452
rect 5353 6443 5411 6449
rect 5353 6440 5365 6443
rect 5224 6412 5365 6440
rect 5224 6400 5230 6412
rect 5353 6409 5365 6412
rect 5399 6440 5411 6443
rect 5994 6440 6000 6452
rect 5399 6412 6000 6440
rect 5399 6409 5411 6412
rect 5353 6403 5411 6409
rect 5994 6400 6000 6412
rect 6052 6400 6058 6452
rect 9950 6400 9956 6452
rect 10008 6440 10014 6452
rect 10321 6443 10379 6449
rect 10321 6440 10333 6443
rect 10008 6412 10333 6440
rect 10008 6400 10014 6412
rect 10321 6409 10333 6412
rect 10367 6409 10379 6443
rect 10321 6403 10379 6409
rect 10686 6400 10692 6452
rect 10744 6440 10750 6452
rect 10781 6443 10839 6449
rect 10781 6440 10793 6443
rect 10744 6412 10793 6440
rect 10744 6400 10750 6412
rect 10781 6409 10793 6412
rect 10827 6409 10839 6443
rect 10781 6403 10839 6409
rect 15562 6400 15568 6452
rect 15620 6400 15626 6452
rect 17954 6400 17960 6452
rect 18012 6400 18018 6452
rect 19242 6440 19248 6452
rect 18064 6412 19248 6440
rect 4246 6381 4252 6384
rect 4240 6372 4252 6381
rect 2056 6344 4016 6372
rect 4207 6344 4252 6372
rect 2056 6313 2084 6344
rect 2041 6307 2099 6313
rect 2041 6273 2053 6307
rect 2087 6273 2099 6307
rect 2041 6267 2099 6273
rect 2308 6307 2366 6313
rect 2308 6273 2320 6307
rect 2354 6304 2366 6307
rect 2354 6276 3924 6304
rect 2354 6273 2366 6276
rect 2308 6267 2366 6273
rect 3896 6100 3924 6276
rect 3988 6248 4016 6344
rect 4240 6335 4252 6344
rect 4246 6332 4252 6335
rect 4304 6332 4310 6384
rect 9861 6375 9919 6381
rect 9861 6341 9873 6375
rect 9907 6372 9919 6375
rect 10870 6372 10876 6384
rect 9907 6344 10876 6372
rect 9907 6341 9919 6344
rect 9861 6335 9919 6341
rect 10870 6332 10876 6344
rect 10928 6332 10934 6384
rect 12526 6332 12532 6384
rect 12584 6372 12590 6384
rect 12989 6375 13047 6381
rect 12989 6372 13001 6375
rect 12584 6344 13001 6372
rect 12584 6332 12590 6344
rect 12989 6341 13001 6344
rect 13035 6372 13047 6375
rect 13262 6372 13268 6384
rect 13035 6344 13268 6372
rect 13035 6341 13047 6344
rect 12989 6335 13047 6341
rect 13262 6332 13268 6344
rect 13320 6332 13326 6384
rect 14737 6375 14795 6381
rect 14737 6341 14749 6375
rect 14783 6372 14795 6375
rect 14918 6372 14924 6384
rect 14783 6344 14924 6372
rect 14783 6341 14795 6344
rect 14737 6335 14795 6341
rect 14918 6332 14924 6344
rect 14976 6332 14982 6384
rect 15010 6332 15016 6384
rect 15068 6372 15074 6384
rect 18064 6372 18092 6412
rect 19242 6400 19248 6412
rect 19300 6400 19306 6452
rect 21726 6400 21732 6452
rect 21784 6440 21790 6452
rect 23201 6443 23259 6449
rect 23201 6440 23213 6443
rect 21784 6412 23213 6440
rect 21784 6400 21790 6412
rect 23201 6409 23213 6412
rect 23247 6409 23259 6443
rect 23201 6403 23259 6409
rect 27246 6400 27252 6452
rect 27304 6400 27310 6452
rect 30469 6443 30527 6449
rect 30469 6409 30481 6443
rect 30515 6440 30527 6443
rect 30558 6440 30564 6452
rect 30515 6412 30564 6440
rect 30515 6409 30527 6412
rect 30469 6403 30527 6409
rect 30558 6400 30564 6412
rect 30616 6400 30622 6452
rect 30650 6400 30656 6452
rect 30708 6400 30714 6452
rect 31018 6400 31024 6452
rect 31076 6440 31082 6452
rect 31113 6443 31171 6449
rect 31113 6440 31125 6443
rect 31076 6412 31125 6440
rect 31076 6400 31082 6412
rect 31113 6409 31125 6412
rect 31159 6409 31171 6443
rect 31113 6403 31171 6409
rect 31386 6400 31392 6452
rect 31444 6440 31450 6452
rect 33870 6440 33876 6452
rect 31444 6412 33876 6440
rect 31444 6400 31450 6412
rect 33870 6400 33876 6412
rect 33928 6440 33934 6452
rect 34422 6440 34428 6452
rect 33928 6412 34428 6440
rect 33928 6400 33934 6412
rect 34422 6400 34428 6412
rect 34480 6440 34486 6452
rect 34480 6412 36124 6440
rect 34480 6400 34486 6412
rect 15068 6344 18092 6372
rect 15068 6332 15074 6344
rect 18598 6332 18604 6384
rect 18656 6372 18662 6384
rect 18656 6344 20484 6372
rect 18656 6332 18662 6344
rect 4522 6264 4528 6316
rect 4580 6304 4586 6316
rect 5997 6307 6055 6313
rect 5997 6304 6009 6307
rect 4580 6276 6009 6304
rect 4580 6264 4586 6276
rect 5997 6273 6009 6276
rect 6043 6273 6055 6307
rect 5997 6267 6055 6273
rect 8478 6264 8484 6316
rect 8536 6264 8542 6316
rect 9030 6264 9036 6316
rect 9088 6304 9094 6316
rect 9125 6307 9183 6313
rect 9125 6304 9137 6307
rect 9088 6276 9137 6304
rect 9088 6264 9094 6276
rect 9125 6273 9137 6276
rect 9171 6273 9183 6307
rect 9125 6267 9183 6273
rect 10962 6264 10968 6316
rect 11020 6264 11026 6316
rect 15749 6307 15807 6313
rect 15749 6273 15761 6307
rect 15795 6304 15807 6307
rect 17126 6304 17132 6316
rect 15795 6276 17132 6304
rect 15795 6273 15807 6276
rect 15749 6267 15807 6273
rect 17126 6264 17132 6276
rect 17184 6264 17190 6316
rect 17954 6307 18012 6313
rect 17954 6273 17966 6307
rect 18000 6304 18012 6307
rect 18230 6304 18236 6316
rect 18000 6276 18236 6304
rect 18000 6273 18012 6276
rect 17954 6267 18012 6273
rect 18230 6264 18236 6276
rect 18288 6264 18294 6316
rect 19150 6264 19156 6316
rect 19208 6264 19214 6316
rect 19242 6264 19248 6316
rect 19300 6264 19306 6316
rect 19334 6264 19340 6316
rect 19392 6264 19398 6316
rect 19521 6307 19579 6313
rect 19521 6273 19533 6307
rect 19567 6273 19579 6307
rect 19521 6267 19579 6273
rect 19981 6307 20039 6313
rect 19981 6273 19993 6307
rect 20027 6304 20039 6307
rect 20346 6304 20352 6316
rect 20027 6276 20352 6304
rect 20027 6273 20039 6276
rect 19981 6267 20039 6273
rect 3970 6196 3976 6248
rect 4028 6196 4034 6248
rect 8938 6196 8944 6248
rect 8996 6196 9002 6248
rect 15470 6196 15476 6248
rect 15528 6236 15534 6248
rect 18417 6239 18475 6245
rect 18417 6236 18429 6239
rect 15528 6208 18429 6236
rect 15528 6196 15534 6208
rect 18417 6205 18429 6208
rect 18463 6236 18475 6239
rect 19426 6236 19432 6248
rect 18463 6208 19432 6236
rect 18463 6205 18475 6208
rect 18417 6199 18475 6205
rect 19426 6196 19432 6208
rect 19484 6196 19490 6248
rect 5813 6171 5871 6177
rect 5813 6168 5825 6171
rect 4908 6140 5825 6168
rect 4908 6100 4936 6140
rect 5813 6137 5825 6140
rect 5859 6137 5871 6171
rect 5813 6131 5871 6137
rect 10134 6128 10140 6180
rect 10192 6168 10198 6180
rect 10229 6171 10287 6177
rect 10229 6168 10241 6171
rect 10192 6140 10241 6168
rect 10192 6128 10198 6140
rect 10229 6137 10241 6140
rect 10275 6168 10287 6171
rect 10870 6168 10876 6180
rect 10275 6140 10876 6168
rect 10275 6137 10287 6140
rect 10229 6131 10287 6137
rect 10870 6128 10876 6140
rect 10928 6128 10934 6180
rect 17773 6171 17831 6177
rect 17773 6137 17785 6171
rect 17819 6168 17831 6171
rect 19536 6168 19564 6267
rect 20346 6264 20352 6276
rect 20404 6264 20410 6316
rect 20456 6313 20484 6344
rect 23750 6332 23756 6384
rect 23808 6332 23814 6384
rect 23969 6375 24027 6381
rect 23969 6341 23981 6375
rect 24015 6372 24027 6375
rect 24578 6372 24584 6384
rect 24015 6344 24584 6372
rect 24015 6341 24027 6344
rect 23969 6335 24027 6341
rect 24578 6332 24584 6344
rect 24636 6332 24642 6384
rect 25866 6332 25872 6384
rect 25924 6332 25930 6384
rect 30668 6372 30696 6400
rect 27356 6344 30696 6372
rect 33321 6375 33379 6381
rect 20441 6307 20499 6313
rect 20441 6273 20453 6307
rect 20487 6304 20499 6307
rect 22738 6304 22744 6316
rect 20487 6276 22744 6304
rect 20487 6273 20499 6276
rect 20441 6267 20499 6273
rect 22738 6264 22744 6276
rect 22796 6264 22802 6316
rect 23106 6264 23112 6316
rect 23164 6264 23170 6316
rect 27062 6264 27068 6316
rect 27120 6304 27126 6316
rect 27356 6313 27384 6344
rect 33321 6341 33333 6375
rect 33367 6372 33379 6375
rect 34241 6375 34299 6381
rect 34241 6372 34253 6375
rect 33367 6344 34253 6372
rect 33367 6341 33379 6344
rect 33321 6335 33379 6341
rect 34241 6341 34253 6344
rect 34287 6341 34299 6375
rect 34241 6335 34299 6341
rect 35066 6332 35072 6384
rect 35124 6372 35130 6384
rect 35124 6344 35664 6372
rect 35124 6332 35130 6344
rect 27157 6307 27215 6313
rect 27157 6304 27169 6307
rect 27120 6276 27169 6304
rect 27120 6264 27126 6276
rect 27157 6273 27169 6276
rect 27203 6273 27215 6307
rect 27157 6267 27215 6273
rect 27341 6307 27399 6313
rect 27341 6273 27353 6307
rect 27387 6273 27399 6307
rect 27341 6267 27399 6273
rect 27614 6264 27620 6316
rect 27672 6304 27678 6316
rect 28629 6307 28687 6313
rect 28629 6304 28641 6307
rect 27672 6276 28641 6304
rect 27672 6264 27678 6276
rect 28629 6273 28641 6276
rect 28675 6273 28687 6307
rect 28629 6267 28687 6273
rect 29270 6264 29276 6316
rect 29328 6264 29334 6316
rect 29733 6307 29791 6313
rect 29733 6273 29745 6307
rect 29779 6273 29791 6307
rect 29733 6267 29791 6273
rect 30653 6307 30711 6313
rect 30653 6273 30665 6307
rect 30699 6304 30711 6307
rect 30742 6304 30748 6316
rect 30699 6276 30748 6304
rect 30699 6273 30711 6276
rect 30653 6267 30711 6273
rect 20162 6196 20168 6248
rect 20220 6196 20226 6248
rect 20806 6196 20812 6248
rect 20864 6196 20870 6248
rect 23474 6196 23480 6248
rect 23532 6236 23538 6248
rect 24486 6236 24492 6248
rect 23532 6208 24492 6236
rect 23532 6196 23538 6208
rect 24486 6196 24492 6208
rect 24544 6236 24550 6248
rect 24581 6239 24639 6245
rect 24581 6236 24593 6239
rect 24544 6208 24593 6236
rect 24544 6196 24550 6208
rect 24581 6205 24593 6208
rect 24627 6205 24639 6239
rect 24857 6239 24915 6245
rect 24857 6236 24869 6239
rect 24581 6199 24639 6205
rect 24688 6208 24869 6236
rect 17819 6140 19564 6168
rect 20073 6171 20131 6177
rect 17819 6137 17831 6140
rect 17773 6131 17831 6137
rect 20073 6137 20085 6171
rect 20119 6168 20131 6171
rect 22554 6168 22560 6180
rect 20119 6140 22560 6168
rect 20119 6137 20131 6140
rect 20073 6131 20131 6137
rect 22554 6128 22560 6140
rect 22612 6128 22618 6180
rect 23014 6128 23020 6180
rect 23072 6168 23078 6180
rect 24688 6168 24716 6208
rect 24857 6205 24869 6208
rect 24903 6205 24915 6239
rect 24857 6199 24915 6205
rect 29178 6196 29184 6248
rect 29236 6236 29242 6248
rect 29748 6236 29776 6267
rect 30742 6264 30748 6276
rect 30800 6264 30806 6316
rect 31297 6307 31355 6313
rect 31297 6273 31309 6307
rect 31343 6304 31355 6307
rect 32306 6304 32312 6316
rect 31343 6276 32312 6304
rect 31343 6273 31355 6276
rect 31297 6267 31355 6273
rect 32306 6264 32312 6276
rect 32364 6264 32370 6316
rect 33229 6307 33287 6313
rect 33229 6273 33241 6307
rect 33275 6273 33287 6307
rect 33229 6267 33287 6273
rect 29236 6208 29776 6236
rect 29236 6196 29242 6208
rect 30006 6196 30012 6248
rect 30064 6196 30070 6248
rect 23072 6140 24716 6168
rect 33244 6168 33272 6267
rect 33870 6264 33876 6316
rect 33928 6264 33934 6316
rect 33965 6307 34023 6313
rect 33965 6273 33977 6307
rect 34011 6304 34023 6307
rect 34054 6304 34060 6316
rect 34011 6276 34060 6304
rect 34011 6273 34023 6276
rect 33965 6267 34023 6273
rect 34054 6264 34060 6276
rect 34112 6264 34118 6316
rect 34149 6307 34207 6313
rect 34149 6273 34161 6307
rect 34195 6273 34207 6307
rect 34149 6267 34207 6273
rect 34333 6307 34391 6313
rect 34333 6273 34345 6307
rect 34379 6304 34391 6307
rect 35342 6304 35348 6316
rect 34379 6276 35348 6304
rect 34379 6273 34391 6276
rect 34333 6267 34391 6273
rect 33686 6196 33692 6248
rect 33744 6236 33750 6248
rect 34164 6236 34192 6267
rect 35342 6264 35348 6276
rect 35400 6264 35406 6316
rect 35434 6264 35440 6316
rect 35492 6264 35498 6316
rect 35636 6313 35664 6344
rect 35621 6307 35679 6313
rect 35621 6273 35633 6307
rect 35667 6273 35679 6307
rect 35621 6267 35679 6273
rect 35713 6307 35771 6313
rect 35713 6273 35725 6307
rect 35759 6304 35771 6307
rect 35986 6304 35992 6316
rect 35759 6276 35992 6304
rect 35759 6273 35771 6276
rect 35713 6267 35771 6273
rect 35986 6264 35992 6276
rect 36044 6264 36050 6316
rect 36096 6304 36124 6412
rect 36446 6400 36452 6452
rect 36504 6440 36510 6452
rect 37550 6440 37556 6452
rect 36504 6412 37556 6440
rect 36504 6400 36510 6412
rect 37550 6400 37556 6412
rect 37608 6400 37614 6452
rect 43714 6440 43720 6452
rect 38580 6412 43720 6440
rect 36262 6332 36268 6384
rect 36320 6372 36326 6384
rect 36320 6344 36676 6372
rect 36320 6332 36326 6344
rect 36648 6313 36676 6344
rect 36633 6307 36691 6313
rect 36096 6276 36584 6304
rect 34514 6236 34520 6248
rect 33744 6208 34520 6236
rect 33744 6196 33750 6208
rect 34514 6196 34520 6208
rect 34572 6196 34578 6248
rect 36556 6245 36584 6276
rect 36633 6273 36645 6307
rect 36679 6273 36691 6307
rect 36633 6267 36691 6273
rect 37366 6264 37372 6316
rect 37424 6304 37430 6316
rect 37461 6307 37519 6313
rect 37461 6304 37473 6307
rect 37424 6276 37473 6304
rect 37424 6264 37430 6276
rect 37461 6273 37473 6276
rect 37507 6273 37519 6307
rect 37461 6267 37519 6273
rect 37642 6264 37648 6316
rect 37700 6264 37706 6316
rect 38473 6307 38531 6313
rect 38473 6273 38485 6307
rect 38519 6304 38531 6307
rect 38580 6304 38608 6412
rect 43714 6400 43720 6412
rect 43772 6400 43778 6452
rect 40865 6375 40923 6381
rect 40865 6341 40877 6375
rect 40911 6372 40923 6375
rect 41325 6375 41383 6381
rect 41325 6372 41337 6375
rect 40911 6344 41337 6372
rect 40911 6341 40923 6344
rect 40865 6335 40923 6341
rect 41325 6341 41337 6344
rect 41371 6341 41383 6375
rect 41325 6335 41383 6341
rect 41432 6344 41644 6372
rect 38519 6276 38608 6304
rect 38519 6273 38531 6276
rect 38473 6267 38531 6273
rect 38654 6264 38660 6316
rect 38712 6264 38718 6316
rect 39022 6264 39028 6316
rect 39080 6304 39086 6316
rect 40589 6307 40647 6313
rect 40589 6304 40601 6307
rect 39080 6276 40601 6304
rect 39080 6264 39086 6276
rect 40589 6273 40601 6276
rect 40635 6273 40647 6307
rect 41432 6304 41460 6344
rect 40589 6267 40647 6273
rect 40779 6276 41460 6304
rect 35253 6239 35311 6245
rect 35253 6205 35265 6239
rect 35299 6236 35311 6239
rect 36449 6239 36507 6245
rect 36449 6236 36461 6239
rect 35299 6228 35388 6236
rect 35452 6228 36461 6236
rect 35299 6208 36461 6228
rect 35299 6205 35311 6208
rect 35253 6199 35311 6205
rect 35360 6200 35480 6208
rect 36449 6205 36461 6208
rect 36495 6205 36507 6239
rect 36449 6199 36507 6205
rect 36541 6239 36599 6245
rect 36541 6205 36553 6239
rect 36587 6236 36599 6239
rect 37274 6236 37280 6248
rect 36587 6208 37280 6236
rect 36587 6205 36599 6208
rect 36541 6199 36599 6205
rect 37274 6196 37280 6208
rect 37332 6196 37338 6248
rect 37660 6236 37688 6264
rect 38749 6239 38807 6245
rect 38749 6236 38761 6239
rect 37660 6208 38761 6236
rect 35529 6171 35587 6177
rect 33244 6140 34008 6168
rect 23072 6128 23078 6140
rect 3896 6072 4936 6100
rect 8294 6060 8300 6112
rect 8352 6060 8358 6112
rect 9306 6060 9312 6112
rect 9364 6060 9370 6112
rect 18322 6060 18328 6112
rect 18380 6060 18386 6112
rect 18877 6103 18935 6109
rect 18877 6069 18889 6103
rect 18923 6100 18935 6103
rect 20622 6100 20628 6112
rect 18923 6072 20628 6100
rect 18923 6069 18935 6072
rect 18877 6063 18935 6069
rect 20622 6060 20628 6072
rect 20680 6060 20686 6112
rect 22462 6060 22468 6112
rect 22520 6100 22526 6112
rect 23937 6103 23995 6109
rect 23937 6100 23949 6103
rect 22520 6072 23949 6100
rect 22520 6060 22526 6072
rect 23937 6069 23949 6072
rect 23983 6069 23995 6103
rect 23937 6063 23995 6069
rect 24118 6060 24124 6112
rect 24176 6060 24182 6112
rect 24854 6060 24860 6112
rect 24912 6100 24918 6112
rect 26329 6103 26387 6109
rect 26329 6100 26341 6103
rect 24912 6072 26341 6100
rect 24912 6060 24918 6072
rect 26329 6069 26341 6072
rect 26375 6069 26387 6103
rect 26329 6063 26387 6069
rect 28445 6103 28503 6109
rect 28445 6069 28457 6103
rect 28491 6100 28503 6103
rect 28994 6100 29000 6112
rect 28491 6072 29000 6100
rect 28491 6069 28503 6072
rect 28445 6063 28503 6069
rect 28994 6060 29000 6072
rect 29052 6060 29058 6112
rect 29086 6060 29092 6112
rect 29144 6060 29150 6112
rect 29822 6060 29828 6112
rect 29880 6060 29886 6112
rect 29914 6060 29920 6112
rect 29972 6060 29978 6112
rect 33410 6060 33416 6112
rect 33468 6100 33474 6112
rect 33873 6103 33931 6109
rect 33873 6100 33885 6103
rect 33468 6072 33885 6100
rect 33468 6060 33474 6072
rect 33873 6069 33885 6072
rect 33919 6069 33931 6103
rect 33980 6100 34008 6140
rect 35529 6137 35541 6171
rect 35575 6168 35587 6171
rect 35618 6168 35624 6180
rect 35575 6140 35624 6168
rect 35575 6137 35587 6140
rect 35529 6131 35587 6137
rect 35618 6128 35624 6140
rect 35676 6128 35682 6180
rect 37660 6168 37688 6208
rect 38749 6205 38761 6208
rect 38795 6205 38807 6239
rect 38749 6199 38807 6205
rect 38841 6239 38899 6245
rect 38841 6205 38853 6239
rect 38887 6205 38899 6239
rect 38841 6199 38899 6205
rect 36188 6140 37688 6168
rect 34974 6100 34980 6112
rect 33980 6072 34980 6100
rect 33873 6063 33931 6069
rect 34974 6060 34980 6072
rect 35032 6100 35038 6112
rect 35342 6100 35348 6112
rect 35032 6072 35348 6100
rect 35032 6060 35038 6072
rect 35342 6060 35348 6072
rect 35400 6060 35406 6112
rect 35434 6060 35440 6112
rect 35492 6100 35498 6112
rect 36188 6100 36216 6140
rect 38562 6128 38568 6180
rect 38620 6168 38626 6180
rect 38856 6168 38884 6199
rect 38620 6140 38884 6168
rect 40604 6168 40632 6267
rect 40678 6196 40684 6248
rect 40736 6236 40742 6248
rect 40779 6236 40807 6276
rect 41506 6264 41512 6316
rect 41564 6264 41570 6316
rect 41616 6313 41644 6344
rect 41601 6307 41659 6313
rect 41601 6273 41613 6307
rect 41647 6273 41659 6307
rect 41601 6267 41659 6273
rect 42797 6307 42855 6313
rect 42797 6273 42809 6307
rect 42843 6273 42855 6307
rect 42797 6267 42855 6273
rect 40736 6208 40807 6236
rect 40865 6239 40923 6245
rect 40736 6196 40742 6208
rect 40865 6205 40877 6239
rect 40911 6236 40923 6239
rect 40954 6236 40960 6248
rect 40911 6208 40960 6236
rect 40911 6205 40923 6208
rect 40865 6199 40923 6205
rect 40954 6196 40960 6208
rect 41012 6196 41018 6248
rect 41397 6239 41455 6245
rect 41397 6205 41409 6239
rect 41443 6236 41455 6239
rect 42812 6236 42840 6267
rect 41443 6208 42840 6236
rect 41443 6205 41455 6208
rect 41397 6199 41455 6205
rect 41506 6168 41512 6180
rect 40604 6140 41512 6168
rect 38620 6128 38626 6140
rect 41506 6128 41512 6140
rect 41564 6128 41570 6180
rect 35492 6072 36216 6100
rect 35492 6060 35498 6072
rect 36262 6060 36268 6112
rect 36320 6060 36326 6112
rect 36906 6060 36912 6112
rect 36964 6100 36970 6112
rect 37461 6103 37519 6109
rect 37461 6100 37473 6103
rect 36964 6072 37473 6100
rect 36964 6060 36970 6072
rect 37461 6069 37473 6072
rect 37507 6069 37519 6103
rect 37461 6063 37519 6069
rect 38746 6060 38752 6112
rect 38804 6100 38810 6112
rect 39209 6103 39267 6109
rect 39209 6100 39221 6103
rect 38804 6072 39221 6100
rect 38804 6060 38810 6072
rect 39209 6069 39221 6072
rect 39255 6069 39267 6103
rect 39209 6063 39267 6069
rect 42610 6060 42616 6112
rect 42668 6060 42674 6112
rect 1104 6010 44896 6032
rect 1104 5958 6423 6010
rect 6475 5958 6487 6010
rect 6539 5958 6551 6010
rect 6603 5958 6615 6010
rect 6667 5958 6679 6010
rect 6731 5958 17370 6010
rect 17422 5958 17434 6010
rect 17486 5958 17498 6010
rect 17550 5958 17562 6010
rect 17614 5958 17626 6010
rect 17678 5958 28317 6010
rect 28369 5958 28381 6010
rect 28433 5958 28445 6010
rect 28497 5958 28509 6010
rect 28561 5958 28573 6010
rect 28625 5958 39264 6010
rect 39316 5958 39328 6010
rect 39380 5958 39392 6010
rect 39444 5958 39456 6010
rect 39508 5958 39520 6010
rect 39572 5958 44896 6010
rect 1104 5936 44896 5958
rect 934 5856 940 5908
rect 992 5896 998 5908
rect 1765 5899 1823 5905
rect 1765 5896 1777 5899
rect 992 5868 1777 5896
rect 992 5856 998 5868
rect 1765 5865 1777 5868
rect 1811 5865 1823 5899
rect 1765 5859 1823 5865
rect 5258 5856 5264 5908
rect 5316 5896 5322 5908
rect 5353 5899 5411 5905
rect 5353 5896 5365 5899
rect 5316 5868 5365 5896
rect 5316 5856 5322 5868
rect 5353 5865 5365 5868
rect 5399 5865 5411 5899
rect 5353 5859 5411 5865
rect 11701 5899 11759 5905
rect 11701 5865 11713 5899
rect 11747 5896 11759 5899
rect 11790 5896 11796 5908
rect 11747 5868 11796 5896
rect 11747 5865 11759 5868
rect 11701 5859 11759 5865
rect 11790 5856 11796 5868
rect 11848 5856 11854 5908
rect 14292 5868 15240 5896
rect 8938 5828 8944 5840
rect 5828 5800 8944 5828
rect 2958 5652 2964 5704
rect 3016 5652 3022 5704
rect 3970 5652 3976 5704
rect 4028 5692 4034 5704
rect 4028 5664 4384 5692
rect 4028 5652 4034 5664
rect 4218 5627 4276 5633
rect 4218 5624 4230 5627
rect 2792 5596 4230 5624
rect 2792 5565 2820 5596
rect 4218 5593 4230 5596
rect 4264 5593 4276 5627
rect 4356 5624 4384 5664
rect 4706 5652 4712 5704
rect 4764 5692 4770 5704
rect 5442 5692 5448 5704
rect 4764 5664 5448 5692
rect 4764 5652 4770 5664
rect 5442 5652 5448 5664
rect 5500 5692 5506 5704
rect 5828 5701 5856 5800
rect 8588 5769 8616 5800
rect 8938 5788 8944 5800
rect 8996 5788 9002 5840
rect 8573 5763 8631 5769
rect 8573 5729 8585 5763
rect 8619 5729 8631 5763
rect 8573 5723 8631 5729
rect 13725 5763 13783 5769
rect 13725 5729 13737 5763
rect 13771 5760 13783 5763
rect 14292 5760 14320 5868
rect 15212 5828 15240 5868
rect 15470 5856 15476 5908
rect 15528 5896 15534 5908
rect 15657 5899 15715 5905
rect 15657 5896 15669 5899
rect 15528 5868 15669 5896
rect 15528 5856 15534 5868
rect 15657 5865 15669 5868
rect 15703 5865 15715 5899
rect 15657 5859 15715 5865
rect 17773 5899 17831 5905
rect 17773 5865 17785 5899
rect 17819 5896 17831 5899
rect 18138 5896 18144 5908
rect 17819 5868 18144 5896
rect 17819 5865 17831 5868
rect 17773 5859 17831 5865
rect 18138 5856 18144 5868
rect 18196 5856 18202 5908
rect 18325 5899 18383 5905
rect 18325 5865 18337 5899
rect 18371 5896 18383 5899
rect 19334 5896 19340 5908
rect 18371 5868 19340 5896
rect 18371 5865 18383 5868
rect 18325 5859 18383 5865
rect 19334 5856 19340 5868
rect 19392 5856 19398 5908
rect 19981 5899 20039 5905
rect 19981 5865 19993 5899
rect 20027 5896 20039 5899
rect 20162 5896 20168 5908
rect 20027 5868 20168 5896
rect 20027 5865 20039 5868
rect 19981 5859 20039 5865
rect 20162 5856 20168 5868
rect 20220 5856 20226 5908
rect 20346 5856 20352 5908
rect 20404 5896 20410 5908
rect 20901 5899 20959 5905
rect 20901 5896 20913 5899
rect 20404 5868 20913 5896
rect 20404 5856 20410 5868
rect 20901 5865 20913 5868
rect 20947 5865 20959 5899
rect 20901 5859 20959 5865
rect 23014 5856 23020 5908
rect 23072 5856 23078 5908
rect 23106 5856 23112 5908
rect 23164 5896 23170 5908
rect 23845 5899 23903 5905
rect 23845 5896 23857 5899
rect 23164 5868 23857 5896
rect 23164 5856 23170 5868
rect 23845 5865 23857 5868
rect 23891 5896 23903 5899
rect 23891 5868 24532 5896
rect 23891 5865 23903 5868
rect 23845 5859 23903 5865
rect 16114 5828 16120 5840
rect 15212 5800 16120 5828
rect 16114 5788 16120 5800
rect 16172 5788 16178 5840
rect 17954 5788 17960 5840
rect 18012 5828 18018 5840
rect 18785 5831 18843 5837
rect 18785 5828 18797 5831
rect 18012 5800 18797 5828
rect 18012 5788 18018 5800
rect 18785 5797 18797 5800
rect 18831 5797 18843 5831
rect 18785 5791 18843 5797
rect 19150 5788 19156 5840
rect 19208 5828 19214 5840
rect 23382 5828 23388 5840
rect 19208 5800 23388 5828
rect 19208 5788 19214 5800
rect 13771 5732 14320 5760
rect 13771 5729 13783 5732
rect 13725 5723 13783 5729
rect 15746 5720 15752 5772
rect 15804 5760 15810 5772
rect 15804 5732 17724 5760
rect 15804 5720 15810 5732
rect 17696 5704 17724 5732
rect 18230 5720 18236 5772
rect 18288 5760 18294 5772
rect 18288 5732 18920 5760
rect 18288 5720 18294 5732
rect 5813 5695 5871 5701
rect 5813 5692 5825 5695
rect 5500 5664 5825 5692
rect 5500 5652 5506 5664
rect 5813 5661 5825 5664
rect 5859 5661 5871 5695
rect 5813 5655 5871 5661
rect 5994 5652 6000 5704
rect 6052 5652 6058 5704
rect 7561 5695 7619 5701
rect 7561 5661 7573 5695
rect 7607 5692 7619 5695
rect 8205 5695 8263 5701
rect 8205 5692 8217 5695
rect 7607 5664 8217 5692
rect 7607 5661 7619 5664
rect 7561 5655 7619 5661
rect 8205 5661 8217 5664
rect 8251 5661 8263 5695
rect 8205 5655 8263 5661
rect 8386 5652 8392 5704
rect 8444 5652 8450 5704
rect 10413 5695 10471 5701
rect 10413 5661 10425 5695
rect 10459 5692 10471 5695
rect 12526 5692 12532 5704
rect 10459 5664 12532 5692
rect 10459 5661 10471 5664
rect 10413 5655 10471 5661
rect 12526 5652 12532 5664
rect 12584 5652 12590 5704
rect 12618 5652 12624 5704
rect 12676 5652 12682 5704
rect 13354 5652 13360 5704
rect 13412 5692 13418 5704
rect 13449 5695 13507 5701
rect 13449 5692 13461 5695
rect 13412 5664 13461 5692
rect 13412 5652 13418 5664
rect 13449 5661 13461 5664
rect 13495 5661 13507 5695
rect 13449 5655 13507 5661
rect 13538 5652 13544 5704
rect 13596 5652 13602 5704
rect 13814 5652 13820 5704
rect 13872 5692 13878 5704
rect 14277 5695 14335 5701
rect 14277 5692 14289 5695
rect 13872 5664 14289 5692
rect 13872 5652 13878 5664
rect 14277 5661 14289 5664
rect 14323 5692 14335 5695
rect 14918 5692 14924 5704
rect 14323 5664 14924 5692
rect 14323 5661 14335 5664
rect 14277 5655 14335 5661
rect 14918 5652 14924 5664
rect 14976 5652 14982 5704
rect 16298 5652 16304 5704
rect 16356 5652 16362 5704
rect 17678 5652 17684 5704
rect 17736 5652 17742 5704
rect 17770 5652 17776 5704
rect 17828 5692 17834 5704
rect 18509 5695 18567 5701
rect 18509 5692 18521 5695
rect 17828 5664 18521 5692
rect 17828 5652 17834 5664
rect 6914 5624 6920 5636
rect 4356 5596 6920 5624
rect 4218 5587 4276 5593
rect 6914 5584 6920 5596
rect 6972 5584 6978 5636
rect 7929 5627 7987 5633
rect 7929 5593 7941 5627
rect 7975 5624 7987 5627
rect 8404 5624 8432 5652
rect 7975 5596 8432 5624
rect 12636 5624 12664 5652
rect 14550 5633 14556 5636
rect 14544 5624 14556 5633
rect 12636 5596 13860 5624
rect 14511 5596 14556 5624
rect 7975 5593 7987 5596
rect 7929 5587 7987 5593
rect 2777 5559 2835 5565
rect 2777 5525 2789 5559
rect 2823 5525 2835 5559
rect 2777 5519 2835 5525
rect 6178 5516 6184 5568
rect 6236 5516 6242 5568
rect 7190 5516 7196 5568
rect 7248 5556 7254 5568
rect 7377 5559 7435 5565
rect 7377 5556 7389 5559
rect 7248 5528 7389 5556
rect 7248 5516 7254 5528
rect 7377 5525 7389 5528
rect 7423 5525 7435 5559
rect 7377 5519 7435 5525
rect 12710 5516 12716 5568
rect 12768 5516 12774 5568
rect 12802 5516 12808 5568
rect 12860 5556 12866 5568
rect 13725 5559 13783 5565
rect 13725 5556 13737 5559
rect 12860 5528 13737 5556
rect 12860 5516 12866 5528
rect 13725 5525 13737 5528
rect 13771 5525 13783 5559
rect 13832 5556 13860 5596
rect 14544 5587 14556 5596
rect 14550 5584 14556 5587
rect 14608 5584 14614 5636
rect 14936 5624 14964 5652
rect 16574 5624 16580 5636
rect 14936 5596 16580 5624
rect 16574 5584 16580 5596
rect 16632 5584 16638 5636
rect 14458 5556 14464 5568
rect 13832 5528 14464 5556
rect 13725 5519 13783 5525
rect 14458 5516 14464 5528
rect 14516 5516 14522 5568
rect 15838 5516 15844 5568
rect 15896 5556 15902 5568
rect 16117 5559 16175 5565
rect 16117 5556 16129 5559
rect 15896 5528 16129 5556
rect 15896 5516 15902 5528
rect 16117 5525 16129 5528
rect 16163 5525 16175 5559
rect 18248 5556 18276 5664
rect 18509 5661 18521 5664
rect 18555 5661 18567 5695
rect 18509 5655 18567 5661
rect 18598 5652 18604 5704
rect 18656 5652 18662 5704
rect 18892 5701 18920 5732
rect 19444 5701 19472 5800
rect 23382 5788 23388 5800
rect 23440 5788 23446 5840
rect 24029 5831 24087 5837
rect 24029 5797 24041 5831
rect 24075 5797 24087 5831
rect 24504 5828 24532 5868
rect 24578 5856 24584 5908
rect 24636 5856 24642 5908
rect 26050 5856 26056 5908
rect 26108 5856 26114 5908
rect 27614 5856 27620 5908
rect 27672 5856 27678 5908
rect 28629 5899 28687 5905
rect 28629 5865 28641 5899
rect 28675 5896 28687 5899
rect 29270 5896 29276 5908
rect 28675 5868 29276 5896
rect 28675 5865 28687 5868
rect 28629 5859 28687 5865
rect 29270 5856 29276 5868
rect 29328 5856 29334 5908
rect 34149 5899 34207 5905
rect 34149 5865 34161 5899
rect 34195 5896 34207 5899
rect 34238 5896 34244 5908
rect 34195 5868 34244 5896
rect 34195 5865 34207 5868
rect 34149 5859 34207 5865
rect 34238 5856 34244 5868
rect 34296 5856 34302 5908
rect 34330 5856 34336 5908
rect 34388 5856 34394 5908
rect 35158 5896 35164 5908
rect 34900 5868 35164 5896
rect 24504 5800 24808 5828
rect 24029 5791 24087 5797
rect 19518 5720 19524 5772
rect 19576 5760 19582 5772
rect 22002 5760 22008 5772
rect 19576 5732 19840 5760
rect 19576 5720 19582 5732
rect 19812 5701 19840 5732
rect 20548 5732 22008 5760
rect 20548 5701 20576 5732
rect 22002 5720 22008 5732
rect 22060 5720 22066 5772
rect 24044 5760 24072 5791
rect 22388 5732 24072 5760
rect 18877 5695 18935 5701
rect 18877 5661 18889 5695
rect 18923 5661 18935 5695
rect 18877 5655 18935 5661
rect 19429 5695 19487 5701
rect 19429 5661 19441 5695
rect 19475 5661 19487 5695
rect 19705 5695 19763 5701
rect 19705 5692 19717 5695
rect 19429 5655 19487 5661
rect 19536 5664 19717 5692
rect 18322 5584 18328 5636
rect 18380 5624 18386 5636
rect 19536 5624 19564 5664
rect 19705 5661 19717 5664
rect 19751 5661 19763 5695
rect 19705 5655 19763 5661
rect 19797 5695 19855 5701
rect 19797 5661 19809 5695
rect 19843 5661 19855 5695
rect 19797 5655 19855 5661
rect 20533 5695 20591 5701
rect 20533 5661 20545 5695
rect 20579 5661 20591 5695
rect 20533 5655 20591 5661
rect 18380 5596 19564 5624
rect 18380 5584 18386 5596
rect 19610 5584 19616 5636
rect 19668 5584 19674 5636
rect 19720 5624 19748 5655
rect 20622 5652 20628 5704
rect 20680 5652 20686 5704
rect 20714 5652 20720 5704
rect 20772 5652 20778 5704
rect 21174 5652 21180 5704
rect 21232 5692 21238 5704
rect 22388 5701 22416 5732
rect 21361 5695 21419 5701
rect 21361 5692 21373 5695
rect 21232 5664 21373 5692
rect 21232 5652 21238 5664
rect 21361 5661 21373 5664
rect 21407 5661 21419 5695
rect 22373 5695 22431 5701
rect 22373 5692 22385 5695
rect 21361 5655 21419 5661
rect 22066 5664 22385 5692
rect 21453 5627 21511 5633
rect 21453 5624 21465 5627
rect 19720 5596 21465 5624
rect 21453 5593 21465 5596
rect 21499 5593 21511 5627
rect 21453 5587 21511 5593
rect 20806 5556 20812 5568
rect 18248 5528 20812 5556
rect 16117 5519 16175 5525
rect 20806 5516 20812 5528
rect 20864 5516 20870 5568
rect 20898 5516 20904 5568
rect 20956 5556 20962 5568
rect 22066 5556 22094 5664
rect 22373 5661 22385 5664
rect 22419 5661 22431 5695
rect 22373 5655 22431 5661
rect 23201 5695 23259 5701
rect 23201 5661 23213 5695
rect 23247 5692 23259 5695
rect 24118 5692 24124 5704
rect 23247 5664 24124 5692
rect 23247 5661 23259 5664
rect 23201 5655 23259 5661
rect 24118 5652 24124 5664
rect 24176 5652 24182 5704
rect 24780 5701 24808 5800
rect 29730 5788 29736 5840
rect 29788 5828 29794 5840
rect 29788 5800 31754 5828
rect 29788 5788 29794 5800
rect 29914 5760 29920 5772
rect 28644 5732 29920 5760
rect 24765 5695 24823 5701
rect 24765 5661 24777 5695
rect 24811 5692 24823 5695
rect 24854 5692 24860 5704
rect 24811 5664 24860 5692
rect 24811 5661 24823 5664
rect 24765 5655 24823 5661
rect 24854 5652 24860 5664
rect 24912 5652 24918 5704
rect 25038 5652 25044 5704
rect 25096 5652 25102 5704
rect 25866 5652 25872 5704
rect 25924 5692 25930 5704
rect 26234 5692 26240 5704
rect 25924 5664 26240 5692
rect 25924 5652 25930 5664
rect 26234 5652 26240 5664
rect 26292 5692 26298 5704
rect 28644 5701 28672 5732
rect 29914 5720 29920 5732
rect 29972 5720 29978 5772
rect 30285 5763 30343 5769
rect 30285 5729 30297 5763
rect 30331 5760 30343 5763
rect 30650 5760 30656 5772
rect 30331 5732 30656 5760
rect 30331 5729 30343 5732
rect 30285 5723 30343 5729
rect 30650 5720 30656 5732
rect 30708 5720 30714 5772
rect 31726 5760 31754 5800
rect 34900 5769 34928 5868
rect 35158 5856 35164 5868
rect 35216 5856 35222 5908
rect 35526 5856 35532 5908
rect 35584 5896 35590 5908
rect 36265 5899 36323 5905
rect 35584 5868 35848 5896
rect 35584 5856 35590 5868
rect 35820 5828 35848 5868
rect 36265 5865 36277 5899
rect 36311 5896 36323 5899
rect 36538 5896 36544 5908
rect 36311 5868 36544 5896
rect 36311 5865 36323 5868
rect 36265 5859 36323 5865
rect 36538 5856 36544 5868
rect 36596 5856 36602 5908
rect 36909 5899 36967 5905
rect 36909 5865 36921 5899
rect 36955 5896 36967 5899
rect 37182 5896 37188 5908
rect 36955 5868 37188 5896
rect 36955 5865 36967 5868
rect 36909 5859 36967 5865
rect 37182 5856 37188 5868
rect 37240 5856 37246 5908
rect 37274 5856 37280 5908
rect 37332 5896 37338 5908
rect 40310 5896 40316 5908
rect 37332 5868 40316 5896
rect 37332 5856 37338 5868
rect 40310 5856 40316 5868
rect 40368 5856 40374 5908
rect 40494 5828 40500 5840
rect 35820 5800 40500 5828
rect 40494 5788 40500 5800
rect 40552 5788 40558 5840
rect 32953 5763 33011 5769
rect 32953 5760 32965 5763
rect 31726 5732 32965 5760
rect 32953 5729 32965 5732
rect 32999 5760 33011 5763
rect 34885 5763 34943 5769
rect 34885 5760 34897 5763
rect 32999 5732 34897 5760
rect 32999 5729 33011 5732
rect 32953 5723 33011 5729
rect 34885 5729 34897 5732
rect 34931 5729 34943 5763
rect 34885 5723 34943 5729
rect 37642 5720 37648 5772
rect 37700 5760 37706 5772
rect 39022 5760 39028 5772
rect 37700 5732 38148 5760
rect 37700 5720 37706 5732
rect 27525 5695 27583 5701
rect 27525 5692 27537 5695
rect 26292 5664 27537 5692
rect 26292 5652 26298 5664
rect 27525 5661 27537 5664
rect 27571 5661 27583 5695
rect 27525 5655 27583 5661
rect 28629 5695 28687 5701
rect 28629 5661 28641 5695
rect 28675 5661 28687 5695
rect 28629 5655 28687 5661
rect 28905 5695 28963 5701
rect 28905 5661 28917 5695
rect 28951 5692 28963 5695
rect 29822 5692 29828 5704
rect 28951 5664 29828 5692
rect 28951 5661 28963 5664
rect 28905 5655 28963 5661
rect 23661 5627 23719 5633
rect 23661 5593 23673 5627
rect 23707 5593 23719 5627
rect 23661 5587 23719 5593
rect 23877 5627 23935 5633
rect 23877 5593 23889 5627
rect 23923 5624 23935 5627
rect 25056 5624 25084 5652
rect 28920 5624 28948 5655
rect 29822 5652 29828 5664
rect 29880 5652 29886 5704
rect 30374 5652 30380 5704
rect 30432 5652 30438 5704
rect 30466 5652 30472 5704
rect 30524 5692 30530 5704
rect 31205 5695 31263 5701
rect 31205 5692 31217 5695
rect 30524 5664 31217 5692
rect 30524 5652 30530 5664
rect 31205 5661 31217 5664
rect 31251 5661 31263 5695
rect 31205 5655 31263 5661
rect 34054 5652 34060 5704
rect 34112 5652 34118 5704
rect 34241 5695 34299 5701
rect 34241 5661 34253 5695
rect 34287 5692 34299 5695
rect 34422 5692 34428 5704
rect 34287 5664 34428 5692
rect 34287 5661 34299 5664
rect 34241 5655 34299 5661
rect 34422 5652 34428 5664
rect 34480 5652 34486 5704
rect 34790 5652 34796 5704
rect 34848 5692 34854 5704
rect 35141 5695 35199 5701
rect 35141 5692 35153 5695
rect 34848 5664 35153 5692
rect 34848 5652 34854 5664
rect 35141 5661 35153 5664
rect 35187 5661 35199 5695
rect 35141 5655 35199 5661
rect 38010 5652 38016 5704
rect 38068 5652 38074 5704
rect 38120 5701 38148 5732
rect 38396 5732 39028 5760
rect 38396 5701 38424 5732
rect 39022 5720 39028 5732
rect 39080 5720 39086 5772
rect 40770 5720 40776 5772
rect 40828 5720 40834 5772
rect 38562 5701 38568 5704
rect 38106 5695 38164 5701
rect 38106 5661 38118 5695
rect 38152 5661 38164 5695
rect 38381 5695 38439 5701
rect 38381 5692 38393 5695
rect 38106 5655 38164 5661
rect 38212 5664 38393 5692
rect 23923 5596 28948 5624
rect 33873 5627 33931 5633
rect 23923 5593 23935 5596
rect 23877 5587 23935 5593
rect 33873 5593 33885 5627
rect 33919 5624 33931 5627
rect 34882 5624 34888 5636
rect 33919 5596 34888 5624
rect 33919 5593 33931 5596
rect 33873 5587 33931 5593
rect 20956 5528 22094 5556
rect 20956 5516 20962 5528
rect 22462 5516 22468 5568
rect 22520 5516 22526 5568
rect 23676 5556 23704 5587
rect 34882 5584 34888 5596
rect 34940 5584 34946 5636
rect 35342 5584 35348 5636
rect 35400 5624 35406 5636
rect 36722 5624 36728 5636
rect 35400 5596 36728 5624
rect 35400 5584 35406 5596
rect 36722 5584 36728 5596
rect 36780 5584 36786 5636
rect 36906 5584 36912 5636
rect 36964 5633 36970 5636
rect 36964 5627 36983 5633
rect 36971 5593 36983 5627
rect 36964 5587 36983 5593
rect 36964 5584 36970 5587
rect 37366 5584 37372 5636
rect 37424 5624 37430 5636
rect 38212 5624 38240 5664
rect 38381 5661 38393 5664
rect 38427 5661 38439 5695
rect 38381 5655 38439 5661
rect 38519 5695 38568 5701
rect 38519 5661 38531 5695
rect 38565 5661 38568 5695
rect 38519 5655 38568 5661
rect 38562 5652 38568 5655
rect 38620 5652 38626 5704
rect 38654 5652 38660 5704
rect 38712 5652 38718 5704
rect 41040 5695 41098 5701
rect 41040 5661 41052 5695
rect 41086 5692 41098 5695
rect 42610 5692 42616 5704
rect 41086 5664 42616 5692
rect 41086 5661 41098 5664
rect 41040 5655 41098 5661
rect 42610 5652 42616 5664
rect 42668 5652 42674 5704
rect 37424 5596 38240 5624
rect 38289 5627 38347 5633
rect 37424 5584 37430 5596
rect 38289 5593 38301 5627
rect 38335 5593 38347 5627
rect 38672 5624 38700 5652
rect 43898 5624 43904 5636
rect 38289 5587 38347 5593
rect 38488 5596 43904 5624
rect 24302 5556 24308 5568
rect 23676 5528 24308 5556
rect 24302 5516 24308 5528
rect 24360 5556 24366 5568
rect 24949 5559 25007 5565
rect 24949 5556 24961 5559
rect 24360 5528 24961 5556
rect 24360 5516 24366 5528
rect 24949 5525 24961 5528
rect 24995 5556 25007 5559
rect 25222 5556 25228 5568
rect 24995 5528 25228 5556
rect 24995 5525 25007 5528
rect 24949 5519 25007 5525
rect 25222 5516 25228 5528
rect 25280 5556 25286 5568
rect 28813 5559 28871 5565
rect 28813 5556 28825 5559
rect 25280 5528 28825 5556
rect 25280 5516 25286 5528
rect 28813 5525 28825 5528
rect 28859 5556 28871 5559
rect 29178 5556 29184 5568
rect 28859 5528 29184 5556
rect 28859 5525 28871 5528
rect 28813 5519 28871 5525
rect 29178 5516 29184 5528
rect 29236 5516 29242 5568
rect 30742 5516 30748 5568
rect 30800 5516 30806 5568
rect 37090 5516 37096 5568
rect 37148 5516 37154 5568
rect 38304 5556 38332 5587
rect 38488 5556 38516 5596
rect 43898 5584 43904 5596
rect 43956 5584 43962 5636
rect 38304 5528 38516 5556
rect 38654 5516 38660 5568
rect 38712 5516 38718 5568
rect 41690 5516 41696 5568
rect 41748 5556 41754 5568
rect 42153 5559 42211 5565
rect 42153 5556 42165 5559
rect 41748 5528 42165 5556
rect 41748 5516 41754 5528
rect 42153 5525 42165 5528
rect 42199 5525 42211 5559
rect 42153 5519 42211 5525
rect 1104 5466 45051 5488
rect 1104 5414 11896 5466
rect 11948 5414 11960 5466
rect 12012 5414 12024 5466
rect 12076 5414 12088 5466
rect 12140 5414 12152 5466
rect 12204 5414 22843 5466
rect 22895 5414 22907 5466
rect 22959 5414 22971 5466
rect 23023 5414 23035 5466
rect 23087 5414 23099 5466
rect 23151 5414 33790 5466
rect 33842 5414 33854 5466
rect 33906 5414 33918 5466
rect 33970 5414 33982 5466
rect 34034 5414 34046 5466
rect 34098 5414 44737 5466
rect 44789 5414 44801 5466
rect 44853 5414 44865 5466
rect 44917 5414 44929 5466
rect 44981 5414 44993 5466
rect 45045 5414 45051 5466
rect 1104 5392 45051 5414
rect 4338 5312 4344 5364
rect 4396 5312 4402 5364
rect 4430 5312 4436 5364
rect 4488 5312 4494 5364
rect 10870 5312 10876 5364
rect 10928 5312 10934 5364
rect 12989 5355 13047 5361
rect 12989 5321 13001 5355
rect 13035 5352 13047 5355
rect 13262 5352 13268 5364
rect 13035 5324 13268 5352
rect 13035 5321 13047 5324
rect 12989 5315 13047 5321
rect 13262 5312 13268 5324
rect 13320 5312 13326 5364
rect 16025 5355 16083 5361
rect 16025 5352 16037 5355
rect 15948 5324 16037 5352
rect 7190 5244 7196 5296
rect 7248 5244 7254 5296
rect 9398 5284 9404 5296
rect 9140 5256 9404 5284
rect 4706 5176 4712 5228
rect 4764 5216 4770 5228
rect 5169 5219 5227 5225
rect 5169 5216 5181 5219
rect 4764 5188 5181 5216
rect 4764 5176 4770 5188
rect 5169 5185 5181 5188
rect 5215 5185 5227 5219
rect 5169 5179 5227 5185
rect 5258 5176 5264 5228
rect 5316 5216 5322 5228
rect 5353 5219 5411 5225
rect 5353 5216 5365 5219
rect 5316 5188 5365 5216
rect 5316 5176 5322 5188
rect 5353 5185 5365 5188
rect 5399 5185 5411 5219
rect 5353 5179 5411 5185
rect 6917 5219 6975 5225
rect 6917 5185 6929 5219
rect 6963 5185 6975 5219
rect 6917 5179 6975 5185
rect 934 5108 940 5160
rect 992 5148 998 5160
rect 1581 5151 1639 5157
rect 1581 5148 1593 5151
rect 992 5120 1593 5148
rect 992 5108 998 5120
rect 1581 5117 1593 5120
rect 1627 5117 1639 5151
rect 1581 5111 1639 5117
rect 1854 5108 1860 5160
rect 1912 5108 1918 5160
rect 4617 5151 4675 5157
rect 4617 5117 4629 5151
rect 4663 5148 4675 5151
rect 5074 5148 5080 5160
rect 4663 5120 5080 5148
rect 4663 5117 4675 5120
rect 4617 5111 4675 5117
rect 5074 5108 5080 5120
rect 5132 5108 5138 5160
rect 6932 5148 6960 5179
rect 8294 5176 8300 5228
rect 8352 5176 8358 5228
rect 9140 5225 9168 5256
rect 9398 5244 9404 5256
rect 9456 5244 9462 5296
rect 10410 5244 10416 5296
rect 10468 5244 10474 5296
rect 12802 5244 12808 5296
rect 12860 5244 12866 5296
rect 13722 5284 13728 5296
rect 13556 5256 13728 5284
rect 9125 5219 9183 5225
rect 9125 5216 9137 5219
rect 8404 5188 9137 5216
rect 8404 5148 8432 5188
rect 9125 5185 9137 5188
rect 9171 5185 9183 5219
rect 9125 5179 9183 5185
rect 12345 5219 12403 5225
rect 12345 5185 12357 5219
rect 12391 5216 12403 5219
rect 12710 5216 12716 5228
rect 12391 5188 12716 5216
rect 12391 5185 12403 5188
rect 12345 5179 12403 5185
rect 12710 5176 12716 5188
rect 12768 5176 12774 5228
rect 13081 5219 13139 5225
rect 13081 5185 13093 5219
rect 13127 5216 13139 5219
rect 13446 5216 13452 5228
rect 13127 5188 13452 5216
rect 13127 5185 13139 5188
rect 13081 5179 13139 5185
rect 13446 5176 13452 5188
rect 13504 5176 13510 5228
rect 13556 5225 13584 5256
rect 13722 5244 13728 5256
rect 13780 5244 13786 5296
rect 15838 5284 15844 5296
rect 15042 5256 15844 5284
rect 15838 5244 15844 5256
rect 15896 5244 15902 5296
rect 13541 5219 13599 5225
rect 13541 5185 13553 5219
rect 13587 5185 13599 5219
rect 13541 5179 13599 5185
rect 15746 5176 15752 5228
rect 15804 5176 15810 5228
rect 6932 5120 8432 5148
rect 8665 5151 8723 5157
rect 8665 5117 8677 5151
rect 8711 5148 8723 5151
rect 9401 5151 9459 5157
rect 9401 5148 9413 5151
rect 8711 5120 9413 5148
rect 8711 5117 8723 5120
rect 8665 5111 8723 5117
rect 9401 5117 9413 5120
rect 9447 5117 9459 5151
rect 9401 5111 9459 5117
rect 13814 5108 13820 5160
rect 13872 5108 13878 5160
rect 15289 5151 15347 5157
rect 15289 5117 15301 5151
rect 15335 5148 15347 5151
rect 15764 5148 15792 5176
rect 15948 5160 15976 5324
rect 16025 5321 16037 5324
rect 16071 5321 16083 5355
rect 16025 5315 16083 5321
rect 17155 5355 17213 5361
rect 17155 5321 17167 5355
rect 17201 5352 17213 5355
rect 17773 5355 17831 5361
rect 17773 5352 17785 5355
rect 17201 5324 17785 5352
rect 17201 5321 17213 5324
rect 17155 5315 17213 5321
rect 17773 5321 17785 5324
rect 17819 5321 17831 5355
rect 17773 5315 17831 5321
rect 17954 5312 17960 5364
rect 18012 5352 18018 5364
rect 20530 5352 20536 5364
rect 18012 5324 20536 5352
rect 18012 5312 18018 5324
rect 20530 5312 20536 5324
rect 20588 5312 20594 5364
rect 22462 5352 22468 5364
rect 20732 5324 22468 5352
rect 16942 5244 16948 5296
rect 17000 5244 17006 5296
rect 18506 5284 18512 5296
rect 18156 5256 18512 5284
rect 17678 5176 17684 5228
rect 17736 5216 17742 5228
rect 18156 5225 18184 5256
rect 18506 5244 18512 5256
rect 18564 5244 18570 5296
rect 18785 5287 18843 5293
rect 18785 5253 18797 5287
rect 18831 5253 18843 5287
rect 19001 5287 19059 5293
rect 19001 5284 19013 5287
rect 18785 5247 18843 5253
rect 18984 5253 19013 5284
rect 19047 5284 19059 5287
rect 19702 5284 19708 5296
rect 19047 5256 19708 5284
rect 19047 5253 19059 5256
rect 18984 5247 19059 5253
rect 18049 5219 18107 5225
rect 18049 5216 18061 5219
rect 17736 5188 18061 5216
rect 17736 5176 17742 5188
rect 18049 5185 18061 5188
rect 18095 5185 18107 5219
rect 18049 5179 18107 5185
rect 18141 5219 18199 5225
rect 18141 5185 18153 5219
rect 18187 5185 18199 5219
rect 18141 5179 18199 5185
rect 18230 5176 18236 5228
rect 18288 5216 18294 5228
rect 18800 5216 18828 5247
rect 18874 5216 18880 5228
rect 18288 5188 18880 5216
rect 18288 5176 18294 5188
rect 18874 5176 18880 5188
rect 18932 5176 18938 5228
rect 15335 5120 15792 5148
rect 15335 5117 15347 5120
rect 15289 5111 15347 5117
rect 15838 5108 15844 5160
rect 15896 5108 15902 5160
rect 15930 5108 15936 5160
rect 15988 5108 15994 5160
rect 16025 5143 16083 5149
rect 16025 5109 16037 5143
rect 16071 5140 16083 5143
rect 16114 5140 16120 5160
rect 16071 5112 16120 5140
rect 16071 5109 16083 5112
rect 16025 5103 16083 5109
rect 16114 5108 16120 5112
rect 16172 5148 16178 5160
rect 16942 5148 16948 5160
rect 16172 5120 16948 5148
rect 16172 5108 16178 5120
rect 16942 5108 16948 5120
rect 17000 5108 17006 5160
rect 17954 5108 17960 5160
rect 18012 5108 18018 5160
rect 18414 5108 18420 5160
rect 18472 5148 18478 5160
rect 18984 5148 19012 5247
rect 19702 5244 19708 5256
rect 19760 5244 19766 5296
rect 19797 5287 19855 5293
rect 19797 5253 19809 5287
rect 19843 5284 19855 5287
rect 20438 5284 20444 5296
rect 19843 5256 20444 5284
rect 19843 5253 19855 5256
rect 19797 5247 19855 5253
rect 19812 5216 19840 5247
rect 20438 5244 20444 5256
rect 20496 5244 20502 5296
rect 18472 5120 19012 5148
rect 19306 5188 19840 5216
rect 19981 5219 20039 5225
rect 18472 5108 18478 5120
rect 3973 5083 4031 5089
rect 3973 5049 3985 5083
rect 4019 5080 4031 5083
rect 4522 5080 4528 5092
rect 4019 5052 4528 5080
rect 4019 5049 4031 5052
rect 3973 5043 4031 5049
rect 4522 5040 4528 5052
rect 4580 5040 4586 5092
rect 18598 5080 18604 5092
rect 17144 5052 18604 5080
rect 5537 5015 5595 5021
rect 5537 4981 5549 5015
rect 5583 5012 5595 5015
rect 7190 5012 7196 5024
rect 5583 4984 7196 5012
rect 5583 4981 5595 4984
rect 5537 4975 5595 4981
rect 7190 4972 7196 4984
rect 7248 4972 7254 5024
rect 12158 4972 12164 5024
rect 12216 4972 12222 5024
rect 12805 5015 12863 5021
rect 12805 4981 12817 5015
rect 12851 5012 12863 5015
rect 12894 5012 12900 5024
rect 12851 4984 12900 5012
rect 12851 4981 12863 4984
rect 12805 4975 12863 4981
rect 12894 4972 12900 4984
rect 12952 4972 12958 5024
rect 17144 5021 17172 5052
rect 18598 5040 18604 5052
rect 18656 5040 18662 5092
rect 17129 5015 17187 5021
rect 17129 4981 17141 5015
rect 17175 4981 17187 5015
rect 17129 4975 17187 4981
rect 17313 5015 17371 5021
rect 17313 4981 17325 5015
rect 17359 5012 17371 5015
rect 17770 5012 17776 5024
rect 17359 4984 17776 5012
rect 17359 4981 17371 4984
rect 17313 4975 17371 4981
rect 17770 4972 17776 4984
rect 17828 4972 17834 5024
rect 18506 4972 18512 5024
rect 18564 5012 18570 5024
rect 18969 5015 19027 5021
rect 18969 5012 18981 5015
rect 18564 4984 18981 5012
rect 18564 4972 18570 4984
rect 18969 4981 18981 4984
rect 19015 4981 19027 5015
rect 18969 4975 19027 4981
rect 19058 4972 19064 5024
rect 19116 5012 19122 5024
rect 19153 5015 19211 5021
rect 19153 5012 19165 5015
rect 19116 4984 19165 5012
rect 19116 4972 19122 4984
rect 19153 4981 19165 4984
rect 19199 5012 19211 5015
rect 19306 5012 19334 5188
rect 19981 5185 19993 5219
rect 20027 5185 20039 5219
rect 19981 5179 20039 5185
rect 20625 5219 20683 5225
rect 20625 5185 20637 5219
rect 20671 5216 20683 5219
rect 20732 5216 20760 5324
rect 22462 5312 22468 5324
rect 22520 5312 22526 5364
rect 22738 5312 22744 5364
rect 22796 5312 22802 5364
rect 24026 5352 24032 5364
rect 23308 5324 24032 5352
rect 20898 5244 20904 5296
rect 20956 5284 20962 5296
rect 23308 5284 23336 5324
rect 24026 5312 24032 5324
rect 24084 5312 24090 5364
rect 28718 5312 28724 5364
rect 28776 5352 28782 5364
rect 28776 5324 41414 5352
rect 28776 5312 28782 5324
rect 20956 5256 21312 5284
rect 20956 5244 20962 5256
rect 20671 5188 20760 5216
rect 20809 5219 20867 5225
rect 20671 5185 20683 5188
rect 20625 5179 20683 5185
rect 20809 5185 20821 5219
rect 20855 5216 20867 5219
rect 20990 5216 20996 5228
rect 20855 5188 20996 5216
rect 20855 5185 20867 5188
rect 20809 5179 20867 5185
rect 19996 5148 20024 5179
rect 20990 5176 20996 5188
rect 21048 5176 21054 5228
rect 21284 5225 21312 5256
rect 22664 5256 23336 5284
rect 22664 5225 22692 5256
rect 23382 5244 23388 5296
rect 23440 5284 23446 5296
rect 26513 5287 26571 5293
rect 26513 5284 26525 5287
rect 23440 5256 26525 5284
rect 23440 5244 23446 5256
rect 23492 5225 23520 5256
rect 21269 5219 21327 5225
rect 21269 5185 21281 5219
rect 21315 5185 21327 5219
rect 21269 5179 21327 5185
rect 21453 5219 21511 5225
rect 21453 5185 21465 5219
rect 21499 5185 21511 5219
rect 21453 5179 21511 5185
rect 22649 5219 22707 5225
rect 22649 5185 22661 5219
rect 22695 5185 22707 5219
rect 22649 5179 22707 5185
rect 23293 5219 23351 5225
rect 23293 5185 23305 5219
rect 23339 5185 23351 5219
rect 23293 5179 23351 5185
rect 23477 5219 23535 5225
rect 23477 5185 23489 5219
rect 23523 5185 23535 5219
rect 23477 5179 23535 5185
rect 21174 5148 21180 5160
rect 19996 5120 21180 5148
rect 21174 5108 21180 5120
rect 21232 5148 21238 5160
rect 21468 5148 21496 5179
rect 23308 5148 23336 5179
rect 23934 5176 23940 5228
rect 23992 5176 23998 5228
rect 24044 5225 24072 5256
rect 26513 5253 26525 5256
rect 26559 5253 26571 5287
rect 26513 5247 26571 5253
rect 28994 5244 29000 5296
rect 29052 5244 29058 5296
rect 33612 5256 35204 5284
rect 24029 5219 24087 5225
rect 24029 5185 24041 5219
rect 24075 5185 24087 5219
rect 24029 5179 24087 5185
rect 24213 5219 24271 5225
rect 24213 5185 24225 5219
rect 24259 5185 24271 5219
rect 24213 5179 24271 5185
rect 24228 5148 24256 5179
rect 24302 5176 24308 5228
rect 24360 5176 24366 5228
rect 24397 5219 24455 5225
rect 24397 5185 24409 5219
rect 24443 5216 24455 5219
rect 24949 5219 25007 5225
rect 24949 5216 24961 5219
rect 24443 5188 24961 5216
rect 24443 5185 24455 5188
rect 24397 5179 24455 5185
rect 24949 5185 24961 5188
rect 24995 5185 25007 5219
rect 24949 5179 25007 5185
rect 24412 5148 24440 5179
rect 25222 5176 25228 5228
rect 25280 5176 25286 5228
rect 25314 5176 25320 5228
rect 25372 5176 25378 5228
rect 25961 5219 26019 5225
rect 25961 5185 25973 5219
rect 26007 5185 26019 5219
rect 25961 5179 26019 5185
rect 26421 5219 26479 5225
rect 26421 5185 26433 5219
rect 26467 5216 26479 5219
rect 27338 5216 27344 5228
rect 26467 5188 27344 5216
rect 26467 5185 26479 5188
rect 26421 5179 26479 5185
rect 21232 5120 21496 5148
rect 22066 5120 24256 5148
rect 24320 5120 24440 5148
rect 24489 5151 24547 5157
rect 21232 5108 21238 5120
rect 19794 5040 19800 5092
rect 19852 5080 19858 5092
rect 20625 5083 20683 5089
rect 20625 5080 20637 5083
rect 19852 5052 20637 5080
rect 19852 5040 19858 5052
rect 20625 5049 20637 5052
rect 20671 5049 20683 5083
rect 20625 5043 20683 5049
rect 19199 4984 19334 5012
rect 19199 4981 19211 4984
rect 19153 4975 19211 4981
rect 20162 4972 20168 5024
rect 20220 4972 20226 5024
rect 21358 4972 21364 5024
rect 21416 5012 21422 5024
rect 22066 5012 22094 5120
rect 22554 5040 22560 5092
rect 22612 5080 22618 5092
rect 24320 5080 24348 5120
rect 24489 5117 24501 5151
rect 24535 5148 24547 5151
rect 25976 5148 26004 5179
rect 27338 5176 27344 5188
rect 27396 5176 27402 5228
rect 33137 5219 33195 5225
rect 33137 5185 33149 5219
rect 33183 5216 33195 5219
rect 33410 5216 33416 5228
rect 33183 5188 33416 5216
rect 33183 5185 33195 5188
rect 33137 5179 33195 5185
rect 33410 5176 33416 5188
rect 33468 5176 33474 5228
rect 33612 5225 33640 5256
rect 35176 5228 35204 5256
rect 37550 5244 37556 5296
rect 37608 5244 37614 5296
rect 38654 5284 38660 5296
rect 38304 5256 38660 5284
rect 33597 5219 33655 5225
rect 33597 5185 33609 5219
rect 33643 5185 33655 5219
rect 33853 5219 33911 5225
rect 33853 5216 33865 5219
rect 33597 5179 33655 5185
rect 33704 5188 33865 5216
rect 24535 5120 26004 5148
rect 24535 5117 24547 5120
rect 24489 5111 24547 5117
rect 27154 5108 27160 5160
rect 27212 5148 27218 5160
rect 28077 5151 28135 5157
rect 28077 5148 28089 5151
rect 27212 5120 28089 5148
rect 27212 5108 27218 5120
rect 28077 5117 28089 5120
rect 28123 5148 28135 5151
rect 28353 5151 28411 5157
rect 28123 5120 28212 5148
rect 28123 5117 28135 5120
rect 28077 5111 28135 5117
rect 22612 5052 24348 5080
rect 22612 5040 22618 5052
rect 21416 4984 22094 5012
rect 23293 5015 23351 5021
rect 21416 4972 21422 4984
rect 23293 4981 23305 5015
rect 23339 5012 23351 5015
rect 23934 5012 23940 5024
rect 23339 4984 23940 5012
rect 23339 4981 23351 4984
rect 23293 4975 23351 4981
rect 23934 4972 23940 4984
rect 23992 4972 23998 5024
rect 25777 5015 25835 5021
rect 25777 4981 25789 5015
rect 25823 5012 25835 5015
rect 25866 5012 25872 5024
rect 25823 4984 25872 5012
rect 25823 4981 25835 4984
rect 25777 4975 25835 4981
rect 25866 4972 25872 4984
rect 25924 4972 25930 5024
rect 28184 5012 28212 5120
rect 28353 5117 28365 5151
rect 28399 5148 28411 5151
rect 29086 5148 29092 5160
rect 28399 5120 29092 5148
rect 28399 5117 28411 5120
rect 28353 5111 28411 5117
rect 29086 5108 29092 5120
rect 29144 5108 29150 5160
rect 29822 5108 29828 5160
rect 29880 5108 29886 5160
rect 33704 5148 33732 5188
rect 33853 5185 33865 5188
rect 33899 5185 33911 5219
rect 33853 5179 33911 5185
rect 35158 5176 35164 5228
rect 35216 5216 35222 5228
rect 35437 5219 35495 5225
rect 35437 5216 35449 5219
rect 35216 5188 35449 5216
rect 35216 5176 35222 5188
rect 35437 5185 35449 5188
rect 35483 5185 35495 5219
rect 35437 5179 35495 5185
rect 35526 5176 35532 5228
rect 35584 5216 35590 5228
rect 35693 5219 35751 5225
rect 35693 5216 35705 5219
rect 35584 5188 35705 5216
rect 35584 5176 35590 5188
rect 35693 5185 35705 5188
rect 35739 5185 35751 5219
rect 35693 5179 35751 5185
rect 37182 5176 37188 5228
rect 37240 5216 37246 5228
rect 38304 5225 38332 5256
rect 38654 5244 38660 5256
rect 38712 5244 38718 5296
rect 38746 5244 38752 5296
rect 38804 5293 38810 5296
rect 38804 5287 38832 5293
rect 38820 5253 38832 5287
rect 38804 5247 38832 5253
rect 38804 5244 38810 5247
rect 41386 5228 41414 5324
rect 41506 5312 41512 5364
rect 41564 5352 41570 5364
rect 41693 5355 41751 5361
rect 41693 5352 41705 5355
rect 41564 5324 41705 5352
rect 41564 5312 41570 5324
rect 41693 5321 41705 5324
rect 41739 5321 41751 5355
rect 41693 5315 41751 5321
rect 37461 5219 37519 5225
rect 37461 5216 37473 5219
rect 37240 5188 37473 5216
rect 37240 5176 37246 5188
rect 37461 5185 37473 5188
rect 37507 5185 37519 5219
rect 37461 5179 37519 5185
rect 38289 5219 38347 5225
rect 38289 5185 38301 5219
rect 38335 5185 38347 5219
rect 41386 5188 41420 5228
rect 38289 5179 38347 5185
rect 41414 5176 41420 5188
rect 41472 5176 41478 5228
rect 41690 5176 41696 5228
rect 41748 5176 41754 5228
rect 42794 5176 42800 5228
rect 42852 5176 42858 5228
rect 32968 5120 33732 5148
rect 32968 5089 32996 5120
rect 38562 5108 38568 5160
rect 38620 5108 38626 5160
rect 38657 5151 38715 5157
rect 38657 5117 38669 5151
rect 38703 5117 38715 5151
rect 38657 5111 38715 5117
rect 43993 5151 44051 5157
rect 43993 5117 44005 5151
rect 44039 5148 44051 5151
rect 44634 5148 44640 5160
rect 44039 5120 44640 5148
rect 44039 5117 44051 5120
rect 43993 5111 44051 5117
rect 32953 5083 33011 5089
rect 32953 5049 32965 5083
rect 32999 5049 33011 5083
rect 38672 5080 38700 5111
rect 44634 5108 44640 5120
rect 44692 5108 44698 5160
rect 32953 5043 33011 5049
rect 34900 5052 35112 5080
rect 29362 5012 29368 5024
rect 28184 4984 29368 5012
rect 29362 4972 29368 4984
rect 29420 4972 29426 5024
rect 30742 4972 30748 5024
rect 30800 5012 30806 5024
rect 34900 5012 34928 5052
rect 30800 4984 34928 5012
rect 30800 4972 30806 4984
rect 34974 4972 34980 5024
rect 35032 4972 35038 5024
rect 35084 5012 35112 5052
rect 36372 5052 38700 5080
rect 36372 5012 36400 5052
rect 38930 5040 38936 5092
rect 38988 5040 38994 5092
rect 35084 4984 36400 5012
rect 36817 5015 36875 5021
rect 36817 4981 36829 5015
rect 36863 5012 36875 5015
rect 37182 5012 37188 5024
rect 36863 4984 37188 5012
rect 36863 4981 36875 4984
rect 36817 4975 36875 4981
rect 37182 4972 37188 4984
rect 37240 4972 37246 5024
rect 1104 4922 44896 4944
rect 1104 4870 6423 4922
rect 6475 4870 6487 4922
rect 6539 4870 6551 4922
rect 6603 4870 6615 4922
rect 6667 4870 6679 4922
rect 6731 4870 17370 4922
rect 17422 4870 17434 4922
rect 17486 4870 17498 4922
rect 17550 4870 17562 4922
rect 17614 4870 17626 4922
rect 17678 4870 28317 4922
rect 28369 4870 28381 4922
rect 28433 4870 28445 4922
rect 28497 4870 28509 4922
rect 28561 4870 28573 4922
rect 28625 4870 39264 4922
rect 39316 4870 39328 4922
rect 39380 4870 39392 4922
rect 39444 4870 39456 4922
rect 39508 4870 39520 4922
rect 39572 4870 44896 4922
rect 1104 4848 44896 4870
rect 10410 4768 10416 4820
rect 10468 4768 10474 4820
rect 13354 4808 13360 4820
rect 11900 4780 13360 4808
rect 1854 4700 1860 4752
rect 1912 4740 1918 4752
rect 11900 4740 11928 4780
rect 13354 4768 13360 4780
rect 13412 4768 13418 4820
rect 14461 4811 14519 4817
rect 14461 4777 14473 4811
rect 14507 4808 14519 4811
rect 16298 4808 16304 4820
rect 14507 4780 16304 4808
rect 14507 4777 14519 4780
rect 14461 4771 14519 4777
rect 16298 4768 16304 4780
rect 16356 4768 16362 4820
rect 18414 4808 18420 4820
rect 16408 4780 18420 4808
rect 1912 4712 11928 4740
rect 1912 4700 1918 4712
rect 13262 4700 13268 4752
rect 13320 4740 13326 4752
rect 13541 4743 13599 4749
rect 13541 4740 13553 4743
rect 13320 4712 13553 4740
rect 13320 4700 13326 4712
rect 13541 4709 13553 4712
rect 13587 4709 13599 4743
rect 13541 4703 13599 4709
rect 4338 4632 4344 4684
rect 4396 4672 4402 4684
rect 4396 4644 4844 4672
rect 4396 4632 4402 4644
rect 4706 4564 4712 4616
rect 4764 4564 4770 4616
rect 4816 4613 4844 4644
rect 11790 4632 11796 4684
rect 11848 4632 11854 4684
rect 12069 4675 12127 4681
rect 12069 4641 12081 4675
rect 12115 4672 12127 4675
rect 12710 4672 12716 4684
rect 12115 4644 12716 4672
rect 12115 4641 12127 4644
rect 12069 4635 12127 4641
rect 12710 4632 12716 4644
rect 12768 4632 12774 4684
rect 15930 4672 15936 4684
rect 15028 4644 15936 4672
rect 4801 4607 4859 4613
rect 4801 4573 4813 4607
rect 4847 4573 4859 4607
rect 4801 4567 4859 4573
rect 9858 4564 9864 4616
rect 9916 4564 9922 4616
rect 9953 4607 10011 4613
rect 9953 4573 9965 4607
rect 9999 4604 10011 4607
rect 10597 4607 10655 4613
rect 10597 4604 10609 4607
rect 9999 4576 10609 4604
rect 9999 4573 10011 4576
rect 9953 4567 10011 4573
rect 10597 4573 10609 4576
rect 10643 4573 10655 4607
rect 10597 4567 10655 4573
rect 14458 4564 14464 4616
rect 14516 4564 14522 4616
rect 15028 4613 15056 4644
rect 15930 4632 15936 4644
rect 15988 4632 15994 4684
rect 15013 4607 15071 4613
rect 15013 4573 15025 4607
rect 15059 4573 15071 4607
rect 15013 4567 15071 4573
rect 15197 4607 15255 4613
rect 15197 4573 15209 4607
rect 15243 4604 15255 4607
rect 16408 4604 16436 4780
rect 18414 4768 18420 4780
rect 18472 4768 18478 4820
rect 18874 4768 18880 4820
rect 18932 4768 18938 4820
rect 21174 4768 21180 4820
rect 21232 4768 21238 4820
rect 23750 4768 23756 4820
rect 23808 4808 23814 4820
rect 24578 4808 24584 4820
rect 23808 4780 24584 4808
rect 23808 4768 23814 4780
rect 24578 4768 24584 4780
rect 24636 4808 24642 4820
rect 25314 4808 25320 4820
rect 24636 4780 25320 4808
rect 24636 4768 24642 4780
rect 25314 4768 25320 4780
rect 25372 4808 25378 4820
rect 25372 4780 26924 4808
rect 25372 4768 25378 4780
rect 21637 4743 21695 4749
rect 21637 4709 21649 4743
rect 21683 4709 21695 4743
rect 21637 4703 21695 4709
rect 16574 4632 16580 4684
rect 16632 4672 16638 4684
rect 17129 4675 17187 4681
rect 17129 4672 17141 4675
rect 16632 4644 17141 4672
rect 16632 4632 16638 4644
rect 17129 4641 17141 4644
rect 17175 4672 17187 4675
rect 18138 4672 18144 4684
rect 17175 4644 18144 4672
rect 17175 4641 17187 4644
rect 17129 4635 17187 4641
rect 18138 4632 18144 4644
rect 18196 4672 18202 4684
rect 19429 4675 19487 4681
rect 19429 4672 19441 4675
rect 18196 4644 19441 4672
rect 18196 4632 18202 4644
rect 19429 4641 19441 4644
rect 19475 4641 19487 4675
rect 19429 4635 19487 4641
rect 19705 4675 19763 4681
rect 19705 4641 19717 4675
rect 19751 4672 19763 4675
rect 21652 4672 21680 4703
rect 23934 4700 23940 4752
rect 23992 4740 23998 4752
rect 26896 4740 26924 4780
rect 27338 4768 27344 4820
rect 27396 4768 27402 4820
rect 34885 4811 34943 4817
rect 34885 4777 34897 4811
rect 34931 4808 34943 4811
rect 35526 4808 35532 4820
rect 34931 4780 35532 4808
rect 34931 4777 34943 4780
rect 34885 4771 34943 4777
rect 35526 4768 35532 4780
rect 35584 4768 35590 4820
rect 37093 4811 37151 4817
rect 37093 4777 37105 4811
rect 37139 4808 37151 4811
rect 38010 4808 38016 4820
rect 37139 4780 38016 4808
rect 37139 4777 37151 4780
rect 37093 4771 37151 4777
rect 38010 4768 38016 4780
rect 38068 4768 38074 4820
rect 38289 4811 38347 4817
rect 38289 4777 38301 4811
rect 38335 4808 38347 4811
rect 38562 4808 38568 4820
rect 38335 4780 38568 4808
rect 38335 4777 38347 4780
rect 38289 4771 38347 4777
rect 38562 4768 38568 4780
rect 38620 4768 38626 4820
rect 30006 4740 30012 4752
rect 23992 4712 25084 4740
rect 26896 4712 30012 4740
rect 23992 4700 23998 4712
rect 19751 4644 21680 4672
rect 19751 4641 19763 4644
rect 19705 4635 19763 4641
rect 23658 4632 23664 4684
rect 23716 4672 23722 4684
rect 24486 4672 24492 4684
rect 23716 4644 24492 4672
rect 23716 4632 23722 4644
rect 24486 4632 24492 4644
rect 24544 4672 24550 4684
rect 24544 4644 24900 4672
rect 24544 4632 24550 4644
rect 15243 4576 16436 4604
rect 15243 4573 15255 4576
rect 15197 4567 15255 4573
rect 12158 4496 12164 4548
rect 12216 4536 12222 4548
rect 12216 4508 12558 4536
rect 12216 4496 12222 4508
rect 13538 4496 13544 4548
rect 13596 4536 13602 4548
rect 15212 4536 15240 4567
rect 21818 4564 21824 4616
rect 21876 4564 21882 4616
rect 23753 4607 23811 4613
rect 23753 4573 23765 4607
rect 23799 4573 23811 4607
rect 23753 4567 23811 4573
rect 13596 4508 15240 4536
rect 13596 4496 13602 4508
rect 17402 4496 17408 4548
rect 17460 4496 17466 4548
rect 19426 4536 19432 4548
rect 18630 4508 19432 4536
rect 19426 4496 19432 4508
rect 19484 4496 19490 4548
rect 20714 4496 20720 4548
rect 20772 4496 20778 4548
rect 23768 4536 23796 4567
rect 24026 4564 24032 4616
rect 24084 4564 24090 4616
rect 24578 4564 24584 4616
rect 24636 4564 24642 4616
rect 24765 4607 24823 4613
rect 24765 4573 24777 4607
rect 24811 4573 24823 4607
rect 24765 4567 24823 4573
rect 24780 4536 24808 4567
rect 23768 4508 24808 4536
rect 24872 4536 24900 4644
rect 25056 4613 25084 4712
rect 30006 4700 30012 4712
rect 30064 4700 30070 4752
rect 25593 4675 25651 4681
rect 25593 4641 25605 4675
rect 25639 4672 25651 4675
rect 29362 4672 29368 4684
rect 25639 4644 29368 4672
rect 25639 4641 25651 4644
rect 25593 4635 25651 4641
rect 25041 4607 25099 4613
rect 25041 4573 25053 4607
rect 25087 4573 25099 4607
rect 25041 4567 25099 4573
rect 25608 4536 25636 4635
rect 29362 4632 29368 4644
rect 29420 4632 29426 4684
rect 36817 4675 36875 4681
rect 36817 4641 36829 4675
rect 36863 4641 36875 4675
rect 36817 4635 36875 4641
rect 28994 4564 29000 4616
rect 29052 4604 29058 4616
rect 29917 4607 29975 4613
rect 29917 4604 29929 4607
rect 29052 4576 29929 4604
rect 29052 4564 29058 4576
rect 29917 4573 29929 4576
rect 29963 4573 29975 4607
rect 29917 4567 29975 4573
rect 30558 4564 30564 4616
rect 30616 4564 30622 4616
rect 35069 4607 35127 4613
rect 35069 4573 35081 4607
rect 35115 4604 35127 4607
rect 36262 4604 36268 4616
rect 35115 4576 36268 4604
rect 35115 4573 35127 4576
rect 35069 4567 35127 4573
rect 36262 4564 36268 4576
rect 36320 4564 36326 4616
rect 36722 4564 36728 4616
rect 36780 4564 36786 4616
rect 36832 4604 36860 4635
rect 37182 4632 37188 4684
rect 37240 4672 37246 4684
rect 38105 4675 38163 4681
rect 37240 4644 38056 4672
rect 37240 4632 37246 4644
rect 37458 4604 37464 4616
rect 36832 4576 37464 4604
rect 37458 4564 37464 4576
rect 37516 4564 37522 4616
rect 38028 4613 38056 4644
rect 38105 4641 38117 4675
rect 38151 4672 38163 4675
rect 44174 4672 44180 4684
rect 38151 4644 44180 4672
rect 38151 4641 38163 4644
rect 38105 4635 38163 4641
rect 44174 4632 44180 4644
rect 44232 4632 44238 4684
rect 38013 4607 38071 4613
rect 38013 4573 38025 4607
rect 38059 4573 38071 4607
rect 38013 4567 38071 4573
rect 24872 4508 25636 4536
rect 25866 4496 25872 4548
rect 25924 4496 25930 4548
rect 26878 4496 26884 4548
rect 26936 4496 26942 4548
rect 4985 4471 5043 4477
rect 4985 4437 4997 4471
rect 5031 4468 5043 4471
rect 5626 4468 5632 4480
rect 5031 4440 5632 4468
rect 5031 4437 5043 4440
rect 4985 4431 5043 4437
rect 5626 4428 5632 4440
rect 5684 4428 5690 4480
rect 15102 4428 15108 4480
rect 15160 4428 15166 4480
rect 23569 4471 23627 4477
rect 23569 4437 23581 4471
rect 23615 4468 23627 4471
rect 24026 4468 24032 4480
rect 23615 4440 24032 4468
rect 23615 4437 23627 4440
rect 23569 4431 23627 4437
rect 24026 4428 24032 4440
rect 24084 4428 24090 4480
rect 24118 4428 24124 4480
rect 24176 4468 24182 4480
rect 24949 4471 25007 4477
rect 24949 4468 24961 4471
rect 24176 4440 24961 4468
rect 24176 4428 24182 4440
rect 24949 4437 24961 4440
rect 24995 4468 25007 4471
rect 25406 4468 25412 4480
rect 24995 4440 25412 4468
rect 24995 4437 25007 4440
rect 24949 4431 25007 4437
rect 25406 4428 25412 4440
rect 25464 4428 25470 4480
rect 29730 4428 29736 4480
rect 29788 4428 29794 4480
rect 30374 4428 30380 4480
rect 30432 4428 30438 4480
rect 1104 4378 45051 4400
rect 1104 4326 11896 4378
rect 11948 4326 11960 4378
rect 12012 4326 12024 4378
rect 12076 4326 12088 4378
rect 12140 4326 12152 4378
rect 12204 4326 22843 4378
rect 22895 4326 22907 4378
rect 22959 4326 22971 4378
rect 23023 4326 23035 4378
rect 23087 4326 23099 4378
rect 23151 4326 33790 4378
rect 33842 4326 33854 4378
rect 33906 4326 33918 4378
rect 33970 4326 33982 4378
rect 34034 4326 34046 4378
rect 34098 4326 44737 4378
rect 44789 4326 44801 4378
rect 44853 4326 44865 4378
rect 44917 4326 44929 4378
rect 44981 4326 44993 4378
rect 45045 4326 45051 4378
rect 1104 4304 45051 4326
rect 12710 4224 12716 4276
rect 12768 4224 12774 4276
rect 13814 4224 13820 4276
rect 13872 4264 13878 4276
rect 14093 4267 14151 4273
rect 14093 4264 14105 4267
rect 13872 4236 14105 4264
rect 13872 4224 13878 4236
rect 14093 4233 14105 4236
rect 14139 4233 14151 4267
rect 14093 4227 14151 4233
rect 16942 4224 16948 4276
rect 17000 4264 17006 4276
rect 17000 4236 17080 4264
rect 17000 4224 17006 4236
rect 17052 4196 17080 4236
rect 17402 4224 17408 4276
rect 17460 4264 17466 4276
rect 17681 4267 17739 4273
rect 17681 4264 17693 4267
rect 17460 4236 17693 4264
rect 17460 4224 17466 4236
rect 17681 4233 17693 4236
rect 17727 4233 17739 4267
rect 17681 4227 17739 4233
rect 18598 4224 18604 4276
rect 18656 4224 18662 4276
rect 20162 4224 20168 4276
rect 20220 4273 20226 4276
rect 20220 4267 20244 4273
rect 20232 4233 20244 4267
rect 20220 4227 20244 4233
rect 20220 4224 20226 4227
rect 23750 4224 23756 4276
rect 23808 4224 23814 4276
rect 25406 4224 25412 4276
rect 25464 4224 25470 4276
rect 25869 4267 25927 4273
rect 25869 4233 25881 4267
rect 25915 4233 25927 4267
rect 25869 4227 25927 4233
rect 19981 4199 20039 4205
rect 19981 4196 19993 4199
rect 17052 4168 19993 4196
rect 19981 4165 19993 4168
rect 20027 4196 20039 4199
rect 23768 4196 23796 4224
rect 25884 4196 25912 4227
rect 20027 4168 23796 4196
rect 25162 4168 25912 4196
rect 20027 4165 20039 4168
rect 19981 4159 20039 4165
rect 29730 4156 29736 4208
rect 29788 4196 29794 4208
rect 29788 4168 30130 4196
rect 29788 4156 29794 4168
rect 9401 4131 9459 4137
rect 9401 4097 9413 4131
rect 9447 4128 9459 4131
rect 9858 4128 9864 4140
rect 9447 4100 9864 4128
rect 9447 4097 9459 4100
rect 9401 4091 9459 4097
rect 9858 4088 9864 4100
rect 9916 4088 9922 4140
rect 12894 4088 12900 4140
rect 12952 4088 12958 4140
rect 14277 4131 14335 4137
rect 14277 4097 14289 4131
rect 14323 4128 14335 4131
rect 15102 4128 15108 4140
rect 14323 4100 15108 4128
rect 14323 4097 14335 4100
rect 14277 4091 14335 4097
rect 15102 4088 15108 4100
rect 15160 4088 15166 4140
rect 16301 4131 16359 4137
rect 16301 4097 16313 4131
rect 16347 4097 16359 4131
rect 16301 4091 16359 4097
rect 16316 4060 16344 4091
rect 16850 4088 16856 4140
rect 16908 4128 16914 4140
rect 16945 4131 17003 4137
rect 16945 4128 16957 4131
rect 16908 4100 16957 4128
rect 16908 4088 16914 4100
rect 16945 4097 16957 4100
rect 16991 4097 17003 4131
rect 16945 4091 17003 4097
rect 17770 4088 17776 4140
rect 17828 4128 17834 4140
rect 17865 4131 17923 4137
rect 17865 4128 17877 4131
rect 17828 4100 17877 4128
rect 17828 4088 17834 4100
rect 17865 4097 17877 4100
rect 17911 4097 17923 4131
rect 17865 4091 17923 4097
rect 18601 4131 18659 4137
rect 18601 4097 18613 4131
rect 18647 4128 18659 4131
rect 19058 4128 19064 4140
rect 18647 4100 19064 4128
rect 18647 4097 18659 4100
rect 18601 4091 18659 4097
rect 19058 4088 19064 4100
rect 19116 4088 19122 4140
rect 19153 4131 19211 4137
rect 19153 4097 19165 4131
rect 19199 4128 19211 4131
rect 19794 4128 19800 4140
rect 19199 4100 19800 4128
rect 19199 4097 19211 4100
rect 19153 4091 19211 4097
rect 19794 4088 19800 4100
rect 19852 4128 19858 4140
rect 20993 4131 21051 4137
rect 20993 4128 21005 4131
rect 19852 4100 21005 4128
rect 19852 4088 19858 4100
rect 20993 4097 21005 4100
rect 21039 4128 21051 4131
rect 21039 4100 22094 4128
rect 21039 4097 21051 4100
rect 20993 4091 21051 4097
rect 21358 4060 21364 4072
rect 16316 4032 16988 4060
rect 8478 3952 8484 4004
rect 8536 3992 8542 4004
rect 16960 4001 16988 4032
rect 20180 4032 21364 4060
rect 9217 3995 9275 4001
rect 9217 3992 9229 3995
rect 8536 3964 9229 3992
rect 8536 3952 8542 3964
rect 9217 3961 9229 3964
rect 9263 3961 9275 3995
rect 9217 3955 9275 3961
rect 16945 3995 17003 4001
rect 16945 3961 16957 3995
rect 16991 3961 17003 3995
rect 16945 3955 17003 3961
rect 16117 3927 16175 3933
rect 16117 3893 16129 3927
rect 16163 3924 16175 3927
rect 16574 3924 16580 3936
rect 16163 3896 16580 3924
rect 16163 3893 16175 3896
rect 16117 3887 16175 3893
rect 16574 3884 16580 3896
rect 16632 3884 16638 3936
rect 19245 3927 19303 3933
rect 19245 3893 19257 3927
rect 19291 3924 19303 3927
rect 19610 3924 19616 3936
rect 19291 3896 19616 3924
rect 19291 3893 19303 3896
rect 19245 3887 19303 3893
rect 19610 3884 19616 3896
rect 19668 3884 19674 3936
rect 20180 3933 20208 4032
rect 21358 4020 21364 4032
rect 21416 4020 21422 4072
rect 20349 3995 20407 4001
rect 20349 3961 20361 3995
rect 20395 3992 20407 3995
rect 21818 3992 21824 4004
rect 20395 3964 21824 3992
rect 20395 3961 20407 3964
rect 20349 3955 20407 3961
rect 21818 3952 21824 3964
rect 21876 3952 21882 4004
rect 20165 3927 20223 3933
rect 20165 3893 20177 3927
rect 20211 3893 20223 3927
rect 20165 3887 20223 3893
rect 20622 3884 20628 3936
rect 20680 3924 20686 3936
rect 20809 3927 20867 3933
rect 20809 3924 20821 3927
rect 20680 3896 20821 3924
rect 20680 3884 20686 3896
rect 20809 3893 20821 3896
rect 20855 3893 20867 3927
rect 22066 3924 22094 4100
rect 23658 4088 23664 4140
rect 23716 4088 23722 4140
rect 26050 4088 26056 4140
rect 26108 4088 26114 4140
rect 27157 4131 27215 4137
rect 27157 4097 27169 4131
rect 27203 4128 27215 4131
rect 28353 4131 28411 4137
rect 28353 4128 28365 4131
rect 27203 4100 28365 4128
rect 27203 4097 27215 4100
rect 27157 4091 27215 4097
rect 28353 4097 28365 4100
rect 28399 4097 28411 4131
rect 28353 4091 28411 4097
rect 28445 4131 28503 4137
rect 28445 4097 28457 4131
rect 28491 4128 28503 4131
rect 28994 4128 29000 4140
rect 28491 4100 29000 4128
rect 28491 4097 28503 4100
rect 28445 4091 28503 4097
rect 23934 4020 23940 4072
rect 23992 4020 23998 4072
rect 25958 4060 25964 4072
rect 24964 4032 25964 4060
rect 24964 3936 24992 4032
rect 25958 4020 25964 4032
rect 26016 4060 26022 4072
rect 27172 4060 27200 4091
rect 28994 4088 29000 4100
rect 29052 4088 29058 4140
rect 29362 4088 29368 4140
rect 29420 4088 29426 4140
rect 31202 4088 31208 4140
rect 31260 4128 31266 4140
rect 31389 4131 31447 4137
rect 31389 4128 31401 4131
rect 31260 4100 31401 4128
rect 31260 4088 31266 4100
rect 31389 4097 31401 4100
rect 31435 4128 31447 4131
rect 31435 4100 31754 4128
rect 31435 4097 31447 4100
rect 31389 4091 31447 4097
rect 26016 4032 27200 4060
rect 29641 4063 29699 4069
rect 26016 4020 26022 4032
rect 29641 4029 29653 4063
rect 29687 4060 29699 4063
rect 30374 4060 30380 4072
rect 29687 4032 30380 4060
rect 29687 4029 29699 4032
rect 29641 4023 29699 4029
rect 30374 4020 30380 4032
rect 30432 4020 30438 4072
rect 31726 4060 31754 4100
rect 41414 4060 41420 4072
rect 31726 4032 41420 4060
rect 41414 4020 41420 4032
rect 41472 4020 41478 4072
rect 24946 3924 24952 3936
rect 22066 3896 24952 3924
rect 20809 3887 20867 3893
rect 24946 3884 24952 3896
rect 25004 3884 25010 3936
rect 26970 3884 26976 3936
rect 27028 3924 27034 3936
rect 27157 3927 27215 3933
rect 27157 3924 27169 3927
rect 27028 3896 27169 3924
rect 27028 3884 27034 3896
rect 27157 3893 27169 3896
rect 27203 3893 27215 3927
rect 27157 3887 27215 3893
rect 1104 3834 44896 3856
rect 1104 3782 6423 3834
rect 6475 3782 6487 3834
rect 6539 3782 6551 3834
rect 6603 3782 6615 3834
rect 6667 3782 6679 3834
rect 6731 3782 17370 3834
rect 17422 3782 17434 3834
rect 17486 3782 17498 3834
rect 17550 3782 17562 3834
rect 17614 3782 17626 3834
rect 17678 3782 28317 3834
rect 28369 3782 28381 3834
rect 28433 3782 28445 3834
rect 28497 3782 28509 3834
rect 28561 3782 28573 3834
rect 28625 3782 39264 3834
rect 39316 3782 39328 3834
rect 39380 3782 39392 3834
rect 39444 3782 39456 3834
rect 39508 3782 39520 3834
rect 39572 3782 44896 3834
rect 1104 3760 44896 3782
rect 19426 3680 19432 3732
rect 19484 3680 19490 3732
rect 20441 3723 20499 3729
rect 20441 3689 20453 3723
rect 20487 3720 20499 3723
rect 20714 3720 20720 3732
rect 20487 3692 20720 3720
rect 20487 3689 20499 3692
rect 20441 3683 20499 3689
rect 20714 3680 20720 3692
rect 20772 3680 20778 3732
rect 23845 3723 23903 3729
rect 23845 3689 23857 3723
rect 23891 3720 23903 3723
rect 23934 3720 23940 3732
rect 23891 3692 23940 3720
rect 23891 3689 23903 3692
rect 23845 3683 23903 3689
rect 23934 3680 23940 3692
rect 23992 3680 23998 3732
rect 24857 3723 24915 3729
rect 24857 3689 24869 3723
rect 24903 3720 24915 3723
rect 26050 3720 26056 3732
rect 24903 3692 26056 3720
rect 24903 3689 24915 3692
rect 24857 3683 24915 3689
rect 26050 3680 26056 3692
rect 26108 3680 26114 3732
rect 26789 3723 26847 3729
rect 26789 3689 26801 3723
rect 26835 3720 26847 3723
rect 26878 3720 26884 3732
rect 26835 3692 26884 3720
rect 26835 3689 26847 3692
rect 26789 3683 26847 3689
rect 26878 3680 26884 3692
rect 26936 3680 26942 3732
rect 30285 3655 30343 3661
rect 30285 3621 30297 3655
rect 30331 3652 30343 3655
rect 30558 3652 30564 3664
rect 30331 3624 30564 3652
rect 30331 3621 30343 3624
rect 30285 3615 30343 3621
rect 30558 3612 30564 3624
rect 30616 3612 30622 3664
rect 6270 3544 6276 3596
rect 6328 3544 6334 3596
rect 30006 3544 30012 3596
rect 30064 3544 30070 3596
rect 934 3476 940 3528
rect 992 3516 998 3528
rect 1765 3519 1823 3525
rect 1765 3516 1777 3519
rect 992 3488 1777 3516
rect 992 3476 998 3488
rect 1765 3485 1777 3488
rect 1811 3485 1823 3519
rect 1765 3479 1823 3485
rect 5626 3476 5632 3528
rect 5684 3476 5690 3528
rect 13541 3519 13599 3525
rect 13541 3485 13553 3519
rect 13587 3516 13599 3519
rect 13722 3516 13728 3528
rect 13587 3488 13728 3516
rect 13587 3485 13599 3488
rect 13541 3479 13599 3485
rect 13722 3476 13728 3488
rect 13780 3476 13786 3528
rect 14737 3519 14795 3525
rect 14737 3485 14749 3519
rect 14783 3516 14795 3519
rect 14826 3516 14832 3528
rect 14783 3488 14832 3516
rect 14783 3485 14795 3488
rect 14737 3479 14795 3485
rect 14826 3476 14832 3488
rect 14884 3476 14890 3528
rect 15378 3476 15384 3528
rect 15436 3476 15442 3528
rect 15841 3519 15899 3525
rect 15841 3485 15853 3519
rect 15887 3516 15899 3519
rect 16114 3516 16120 3528
rect 15887 3488 16120 3516
rect 15887 3485 15899 3488
rect 15841 3479 15899 3485
rect 16114 3476 16120 3488
rect 16172 3476 16178 3528
rect 16206 3476 16212 3528
rect 16264 3476 16270 3528
rect 18138 3476 18144 3528
rect 18196 3476 18202 3528
rect 19610 3476 19616 3528
rect 19668 3476 19674 3528
rect 20622 3476 20628 3528
rect 20680 3476 20686 3528
rect 24026 3476 24032 3528
rect 24084 3476 24090 3528
rect 24765 3519 24823 3525
rect 24765 3485 24777 3519
rect 24811 3516 24823 3519
rect 24946 3516 24952 3528
rect 24811 3488 24952 3516
rect 24811 3485 24823 3488
rect 24765 3479 24823 3485
rect 24946 3476 24952 3488
rect 25004 3476 25010 3528
rect 26970 3476 26976 3528
rect 27028 3476 27034 3528
rect 29917 3519 29975 3525
rect 29917 3485 29929 3519
rect 29963 3516 29975 3519
rect 31202 3516 31208 3528
rect 29963 3488 31208 3516
rect 29963 3485 29975 3488
rect 29917 3479 29975 3485
rect 31202 3476 31208 3488
rect 31260 3476 31266 3528
rect 44361 3519 44419 3525
rect 44361 3485 44373 3519
rect 44407 3516 44419 3519
rect 44634 3516 44640 3528
rect 44407 3488 44640 3516
rect 44407 3485 44419 3488
rect 44361 3479 44419 3485
rect 44634 3476 44640 3488
rect 44692 3476 44698 3528
rect 16574 3408 16580 3460
rect 16632 3408 16638 3460
rect 17635 3451 17693 3457
rect 17635 3417 17647 3451
rect 17681 3448 17693 3451
rect 18046 3448 18052 3460
rect 17681 3420 18052 3448
rect 17681 3417 17693 3420
rect 17635 3411 17693 3417
rect 18046 3408 18052 3420
rect 18104 3408 18110 3460
rect 23290 3408 23296 3460
rect 23348 3448 23354 3460
rect 33502 3448 33508 3460
rect 23348 3420 33508 3448
rect 23348 3408 23354 3420
rect 33502 3408 33508 3420
rect 33560 3408 33566 3460
rect 13630 3340 13636 3392
rect 13688 3340 13694 3392
rect 15194 3340 15200 3392
rect 15252 3340 15258 3392
rect 17770 3340 17776 3392
rect 17828 3380 17834 3392
rect 18233 3383 18291 3389
rect 18233 3380 18245 3383
rect 17828 3352 18245 3380
rect 17828 3340 17834 3352
rect 18233 3349 18245 3352
rect 18279 3349 18291 3383
rect 18233 3343 18291 3349
rect 1104 3290 45051 3312
rect 1104 3238 11896 3290
rect 11948 3238 11960 3290
rect 12012 3238 12024 3290
rect 12076 3238 12088 3290
rect 12140 3238 12152 3290
rect 12204 3238 22843 3290
rect 22895 3238 22907 3290
rect 22959 3238 22971 3290
rect 23023 3238 23035 3290
rect 23087 3238 23099 3290
rect 23151 3238 33790 3290
rect 33842 3238 33854 3290
rect 33906 3238 33918 3290
rect 33970 3238 33982 3290
rect 34034 3238 34046 3290
rect 34098 3238 44737 3290
rect 44789 3238 44801 3290
rect 44853 3238 44865 3290
rect 44917 3238 44929 3290
rect 44981 3238 44993 3290
rect 45045 3238 45051 3290
rect 1104 3216 45051 3238
rect 9306 3136 9312 3188
rect 9364 3176 9370 3188
rect 9364 3148 16068 3176
rect 9364 3136 9370 3148
rect 15194 3068 15200 3120
rect 15252 3068 15258 3120
rect 16040 3108 16068 3148
rect 16114 3136 16120 3188
rect 16172 3176 16178 3188
rect 17037 3179 17095 3185
rect 17037 3176 17049 3179
rect 16172 3148 17049 3176
rect 16172 3136 16178 3148
rect 17037 3145 17049 3148
rect 17083 3145 17095 3179
rect 17037 3139 17095 3145
rect 17144 3148 31754 3176
rect 17144 3108 17172 3148
rect 16040 3080 17172 3108
rect 7190 3000 7196 3052
rect 7248 3000 7254 3052
rect 13630 3000 13636 3052
rect 13688 3000 13694 3052
rect 14826 3000 14832 3052
rect 14884 3000 14890 3052
rect 16206 3000 16212 3052
rect 16264 3049 16270 3052
rect 16264 3043 16313 3049
rect 16264 3009 16267 3043
rect 16301 3009 16313 3043
rect 16264 3003 16313 3009
rect 16853 3043 16911 3049
rect 16853 3009 16865 3043
rect 16899 3040 16911 3043
rect 17770 3040 17776 3052
rect 16899 3012 17776 3040
rect 16899 3009 16911 3012
rect 16853 3003 16911 3009
rect 16264 3000 16270 3003
rect 17770 3000 17776 3012
rect 17828 3000 17834 3052
rect 18046 3000 18052 3052
rect 18104 3000 18110 3052
rect 8389 2975 8447 2981
rect 8389 2941 8401 2975
rect 8435 2972 8447 2975
rect 9674 2972 9680 2984
rect 8435 2944 9680 2972
rect 8435 2941 8447 2944
rect 8389 2935 8447 2941
rect 9674 2932 9680 2944
rect 9732 2932 9738 2984
rect 14461 2975 14519 2981
rect 14461 2941 14473 2975
rect 14507 2941 14519 2975
rect 14461 2935 14519 2941
rect 13817 2907 13875 2913
rect 13817 2873 13829 2907
rect 13863 2904 13875 2907
rect 14476 2904 14504 2935
rect 17126 2932 17132 2984
rect 17184 2972 17190 2984
rect 17681 2975 17739 2981
rect 17681 2972 17693 2975
rect 17184 2944 17693 2972
rect 17184 2932 17190 2944
rect 17681 2941 17693 2944
rect 17727 2941 17739 2975
rect 17681 2935 17739 2941
rect 13863 2876 14504 2904
rect 19076 2904 19104 3094
rect 19794 3068 19800 3120
rect 19852 3068 19858 3120
rect 20441 3043 20499 3049
rect 20441 3009 20453 3043
rect 20487 3009 20499 3043
rect 20441 3003 20499 3009
rect 20257 2907 20315 2913
rect 20257 2904 20269 2907
rect 19076 2876 20269 2904
rect 13863 2873 13875 2876
rect 13817 2867 13875 2873
rect 20257 2873 20269 2876
rect 20303 2873 20315 2907
rect 20257 2867 20315 2873
rect 934 2796 940 2848
rect 992 2836 998 2848
rect 1765 2839 1823 2845
rect 1765 2836 1777 2839
rect 992 2808 1777 2836
rect 992 2796 998 2808
rect 1765 2805 1777 2808
rect 1811 2805 1823 2839
rect 1765 2799 1823 2805
rect 18874 2796 18880 2848
rect 18932 2836 18938 2848
rect 20456 2836 20484 3003
rect 22646 3000 22652 3052
rect 22704 3040 22710 3052
rect 22925 3043 22983 3049
rect 22925 3040 22937 3043
rect 22704 3012 22937 3040
rect 22704 3000 22710 3012
rect 22925 3009 22937 3012
rect 22971 3009 22983 3043
rect 31726 3040 31754 3148
rect 44174 3136 44180 3188
rect 44232 3136 44238 3188
rect 34241 3043 34299 3049
rect 34241 3040 34253 3043
rect 31726 3012 34253 3040
rect 22925 3003 22983 3009
rect 34241 3009 34253 3012
rect 34287 3009 34299 3043
rect 34241 3003 34299 3009
rect 44361 3043 44419 3049
rect 44361 3009 44373 3043
rect 44407 3040 44419 3043
rect 45094 3040 45100 3052
rect 44407 3012 45100 3040
rect 44407 3009 44419 3012
rect 44361 3003 44419 3009
rect 45094 3000 45100 3012
rect 45152 3000 45158 3052
rect 22554 2932 22560 2984
rect 22612 2972 22618 2984
rect 23385 2975 23443 2981
rect 23385 2972 23397 2975
rect 22612 2944 23397 2972
rect 22612 2932 22618 2944
rect 23385 2941 23397 2944
rect 23431 2941 23443 2975
rect 23385 2935 23443 2941
rect 35434 2932 35440 2984
rect 35492 2932 35498 2984
rect 18932 2808 20484 2836
rect 18932 2796 18938 2808
rect 1104 2746 44896 2768
rect 1104 2694 6423 2746
rect 6475 2694 6487 2746
rect 6539 2694 6551 2746
rect 6603 2694 6615 2746
rect 6667 2694 6679 2746
rect 6731 2694 17370 2746
rect 17422 2694 17434 2746
rect 17486 2694 17498 2746
rect 17550 2694 17562 2746
rect 17614 2694 17626 2746
rect 17678 2694 28317 2746
rect 28369 2694 28381 2746
rect 28433 2694 28445 2746
rect 28497 2694 28509 2746
rect 28561 2694 28573 2746
rect 28625 2694 39264 2746
rect 39316 2694 39328 2746
rect 39380 2694 39392 2746
rect 39444 2694 39456 2746
rect 39508 2694 39520 2746
rect 39572 2694 44896 2746
rect 1104 2672 44896 2694
rect 12802 2592 12808 2644
rect 12860 2632 12866 2644
rect 12897 2635 12955 2641
rect 12897 2632 12909 2635
rect 12860 2604 12909 2632
rect 12860 2592 12866 2604
rect 12897 2601 12909 2604
rect 12943 2601 12955 2635
rect 12897 2595 12955 2601
rect 14829 2635 14887 2641
rect 14829 2601 14841 2635
rect 14875 2632 14887 2635
rect 15378 2632 15384 2644
rect 14875 2604 15384 2632
rect 14875 2601 14887 2604
rect 14829 2595 14887 2601
rect 15378 2592 15384 2604
rect 15436 2592 15442 2644
rect 16209 2635 16267 2641
rect 16209 2601 16221 2635
rect 16255 2632 16267 2635
rect 17126 2632 17132 2644
rect 16255 2604 17132 2632
rect 16255 2601 16267 2604
rect 16209 2595 16267 2601
rect 17126 2592 17132 2604
rect 17184 2592 17190 2644
rect 17862 2592 17868 2644
rect 17920 2632 17926 2644
rect 17920 2604 26234 2632
rect 17920 2592 17926 2604
rect 13725 2567 13783 2573
rect 13725 2533 13737 2567
rect 13771 2564 13783 2567
rect 16114 2564 16120 2576
rect 13771 2536 16120 2564
rect 13771 2533 13783 2536
rect 13725 2527 13783 2533
rect 16114 2524 16120 2536
rect 16172 2524 16178 2576
rect 16945 2567 17003 2573
rect 16945 2533 16957 2567
rect 16991 2564 17003 2567
rect 18874 2564 18880 2576
rect 16991 2536 18880 2564
rect 16991 2533 17003 2536
rect 16945 2527 17003 2533
rect 18874 2524 18880 2536
rect 18932 2524 18938 2576
rect 14 2456 20 2508
rect 72 2496 78 2508
rect 2409 2499 2467 2505
rect 2409 2496 2421 2499
rect 72 2468 2421 2496
rect 72 2456 78 2468
rect 2409 2465 2421 2468
rect 2455 2465 2467 2499
rect 18138 2496 18144 2508
rect 2409 2459 2467 2465
rect 15396 2468 18144 2496
rect 1302 2388 1308 2440
rect 1360 2428 1366 2440
rect 1765 2431 1823 2437
rect 1765 2428 1777 2431
rect 1360 2400 1777 2428
rect 1360 2388 1366 2400
rect 1765 2397 1777 2400
rect 1811 2397 1823 2431
rect 1765 2391 1823 2397
rect 4154 2388 4160 2440
rect 4212 2388 4218 2440
rect 4522 2388 4528 2440
rect 4580 2428 4586 2440
rect 4801 2431 4859 2437
rect 4801 2428 4813 2431
rect 4580 2400 4813 2428
rect 4580 2388 4586 2400
rect 4801 2397 4813 2400
rect 4847 2397 4859 2431
rect 4801 2391 4859 2397
rect 7742 2388 7748 2440
rect 7800 2428 7806 2440
rect 8021 2431 8079 2437
rect 8021 2428 8033 2431
rect 7800 2400 8033 2428
rect 7800 2388 7806 2400
rect 8021 2397 8033 2400
rect 8067 2397 8079 2431
rect 8021 2391 8079 2397
rect 11054 2388 11060 2440
rect 11112 2428 11118 2440
rect 11885 2431 11943 2437
rect 11885 2428 11897 2431
rect 11112 2400 11897 2428
rect 11112 2388 11118 2400
rect 11885 2397 11897 2400
rect 11931 2397 11943 2431
rect 11885 2391 11943 2397
rect 12894 2388 12900 2440
rect 12952 2428 12958 2440
rect 15396 2437 15424 2468
rect 18138 2456 18144 2468
rect 18196 2456 18202 2508
rect 26206 2496 26234 2604
rect 27522 2592 27528 2644
rect 27580 2592 27586 2644
rect 32490 2592 32496 2644
rect 32548 2592 32554 2644
rect 37458 2592 37464 2644
rect 37516 2592 37522 2644
rect 43898 2592 43904 2644
rect 43956 2592 43962 2644
rect 42889 2499 42947 2505
rect 42889 2496 42901 2499
rect 26206 2468 42901 2496
rect 42889 2465 42901 2468
rect 42935 2465 42947 2499
rect 42889 2459 42947 2465
rect 13081 2431 13139 2437
rect 13081 2428 13093 2431
rect 12952 2400 13093 2428
rect 12952 2388 12958 2400
rect 13081 2397 13093 2400
rect 13127 2397 13139 2431
rect 13081 2391 13139 2397
rect 14737 2431 14795 2437
rect 14737 2397 14749 2431
rect 14783 2397 14795 2431
rect 14737 2391 14795 2397
rect 15381 2431 15439 2437
rect 15381 2397 15393 2431
rect 15427 2397 15439 2431
rect 15381 2391 15439 2397
rect 15473 2431 15531 2437
rect 15473 2397 15485 2431
rect 15519 2428 15531 2431
rect 16025 2431 16083 2437
rect 16025 2428 16037 2431
rect 15519 2400 16037 2428
rect 15519 2397 15531 2400
rect 15473 2391 15531 2397
rect 16025 2397 16037 2400
rect 16071 2397 16083 2431
rect 16850 2428 16856 2440
rect 16025 2391 16083 2397
rect 16546 2400 16856 2428
rect 14752 2360 14780 2391
rect 16546 2360 16574 2400
rect 16850 2388 16856 2400
rect 16908 2388 16914 2440
rect 17402 2388 17408 2440
rect 17460 2428 17466 2440
rect 17497 2431 17555 2437
rect 17497 2428 17509 2431
rect 17460 2400 17509 2428
rect 17460 2388 17466 2400
rect 17497 2397 17509 2400
rect 17543 2397 17555 2431
rect 17497 2391 17555 2397
rect 17773 2431 17831 2437
rect 17773 2397 17785 2431
rect 17819 2397 17831 2431
rect 17773 2391 17831 2397
rect 14752 2332 16574 2360
rect 16868 2360 16896 2388
rect 17788 2360 17816 2391
rect 19334 2388 19340 2440
rect 19392 2428 19398 2440
rect 19613 2431 19671 2437
rect 19613 2428 19625 2431
rect 19392 2400 19625 2428
rect 19392 2388 19398 2400
rect 19613 2397 19625 2400
rect 19659 2397 19671 2431
rect 19613 2391 19671 2397
rect 20714 2388 20720 2440
rect 20772 2428 20778 2440
rect 20901 2431 20959 2437
rect 20901 2428 20913 2431
rect 20772 2400 20913 2428
rect 20772 2388 20778 2400
rect 20901 2397 20913 2400
rect 20947 2397 20959 2431
rect 20901 2391 20959 2397
rect 23842 2388 23848 2440
rect 23900 2428 23906 2440
rect 24765 2431 24823 2437
rect 24765 2428 24777 2431
rect 23900 2400 24777 2428
rect 23900 2388 23906 2400
rect 24765 2397 24777 2400
rect 24811 2397 24823 2431
rect 24765 2391 24823 2397
rect 25774 2388 25780 2440
rect 25832 2428 25838 2440
rect 26053 2431 26111 2437
rect 26053 2428 26065 2431
rect 25832 2400 26065 2428
rect 25832 2388 25838 2400
rect 26053 2397 26065 2400
rect 26099 2397 26111 2431
rect 26053 2391 26111 2397
rect 28994 2388 29000 2440
rect 29052 2428 29058 2440
rect 29917 2431 29975 2437
rect 29917 2428 29929 2431
rect 29052 2400 29929 2428
rect 29052 2388 29058 2400
rect 29917 2397 29929 2400
rect 29963 2397 29975 2431
rect 29917 2391 29975 2397
rect 30374 2388 30380 2440
rect 30432 2428 30438 2440
rect 30561 2431 30619 2437
rect 30561 2428 30573 2431
rect 30432 2400 30573 2428
rect 30432 2388 30438 2400
rect 30561 2397 30573 2400
rect 30607 2397 30619 2431
rect 30561 2391 30619 2397
rect 37642 2388 37648 2440
rect 37700 2388 37706 2440
rect 38654 2388 38660 2440
rect 38712 2428 38718 2440
rect 38933 2431 38991 2437
rect 38933 2428 38945 2431
rect 38712 2400 38945 2428
rect 38712 2388 38718 2400
rect 38933 2397 38945 2400
rect 38979 2397 38991 2431
rect 38933 2391 38991 2397
rect 40034 2388 40040 2440
rect 40092 2428 40098 2440
rect 40221 2431 40279 2437
rect 40221 2428 40233 2431
rect 40092 2400 40233 2428
rect 40092 2388 40098 2400
rect 40221 2397 40233 2400
rect 40267 2397 40279 2431
rect 40221 2391 40279 2397
rect 43806 2388 43812 2440
rect 43864 2428 43870 2440
rect 44085 2431 44143 2437
rect 44085 2428 44097 2431
rect 43864 2400 44097 2428
rect 43864 2388 43870 2400
rect 44085 2397 44097 2400
rect 44131 2397 44143 2431
rect 44085 2391 44143 2397
rect 16868 2332 17816 2360
rect 27062 2320 27068 2372
rect 27120 2360 27126 2372
rect 27249 2363 27307 2369
rect 27249 2360 27261 2363
rect 27120 2332 27261 2360
rect 27120 2320 27126 2332
rect 27249 2329 27261 2332
rect 27295 2329 27307 2363
rect 27249 2323 27307 2329
rect 32214 2320 32220 2372
rect 32272 2360 32278 2372
rect 32401 2363 32459 2369
rect 32401 2360 32413 2363
rect 32272 2332 32413 2360
rect 32272 2320 32278 2332
rect 32401 2329 32413 2332
rect 32447 2329 32459 2363
rect 32401 2323 32459 2329
rect 41874 2320 41880 2372
rect 41932 2360 41938 2372
rect 42705 2363 42763 2369
rect 42705 2360 42717 2363
rect 41932 2332 42717 2360
rect 41932 2320 41938 2332
rect 42705 2329 42717 2332
rect 42751 2329 42763 2363
rect 42705 2323 42763 2329
rect 25869 2295 25927 2301
rect 25869 2261 25881 2295
rect 25915 2292 25927 2295
rect 30650 2292 30656 2304
rect 25915 2264 30656 2292
rect 25915 2261 25927 2264
rect 25869 2255 25927 2261
rect 30650 2252 30656 2264
rect 30708 2252 30714 2304
rect 1104 2202 45051 2224
rect 1104 2150 11896 2202
rect 11948 2150 11960 2202
rect 12012 2150 12024 2202
rect 12076 2150 12088 2202
rect 12140 2150 12152 2202
rect 12204 2150 22843 2202
rect 22895 2150 22907 2202
rect 22959 2150 22971 2202
rect 23023 2150 23035 2202
rect 23087 2150 23099 2202
rect 23151 2150 33790 2202
rect 33842 2150 33854 2202
rect 33906 2150 33918 2202
rect 33970 2150 33982 2202
rect 34034 2150 34046 2202
rect 34098 2150 44737 2202
rect 44789 2150 44801 2202
rect 44853 2150 44865 2202
rect 44917 2150 44929 2202
rect 44981 2150 44993 2202
rect 45045 2150 45051 2202
rect 1104 2128 45051 2150
rect 3234 892 3240 944
rect 3292 932 3298 944
rect 4154 932 4160 944
rect 3292 904 4160 932
rect 3292 892 3298 904
rect 4154 892 4160 904
rect 4212 892 4218 944
rect 36722 892 36728 944
rect 36780 932 36786 944
rect 37642 932 37648 944
rect 36780 904 37648 932
rect 36780 892 36786 904
rect 37642 892 37648 904
rect 37700 892 37706 944
<< via1 >>
rect 16120 19048 16172 19100
rect 16856 19048 16908 19100
rect 34152 19048 34204 19100
rect 35072 19048 35124 19100
rect 41880 19048 41932 19100
rect 42800 19048 42852 19100
rect 43444 18028 43496 18080
rect 45008 18028 45060 18080
rect 43996 17484 44048 17536
rect 45008 17484 45060 17536
rect 11896 17382 11948 17434
rect 11960 17382 12012 17434
rect 12024 17382 12076 17434
rect 12088 17382 12140 17434
rect 12152 17382 12204 17434
rect 22843 17382 22895 17434
rect 22907 17382 22959 17434
rect 22971 17382 23023 17434
rect 23035 17382 23087 17434
rect 23099 17382 23151 17434
rect 33790 17382 33842 17434
rect 33854 17382 33906 17434
rect 33918 17382 33970 17434
rect 33982 17382 34034 17434
rect 34046 17382 34098 17434
rect 44737 17382 44789 17434
rect 44801 17382 44853 17434
rect 44865 17382 44917 17434
rect 44929 17382 44981 17434
rect 44993 17382 45045 17434
rect 940 17212 992 17264
rect 3240 17255 3292 17264
rect 3240 17221 3249 17255
rect 3249 17221 3283 17255
rect 3283 17221 3292 17255
rect 3240 17212 3292 17221
rect 11060 17212 11112 17264
rect 38660 17212 38712 17264
rect 1308 17144 1360 17196
rect 4528 17144 4580 17196
rect 6460 17144 6512 17196
rect 7748 17144 7800 17196
rect 9680 17144 9732 17196
rect 12900 17144 12952 17196
rect 14188 17144 14240 17196
rect 16856 17187 16908 17196
rect 16856 17153 16865 17187
rect 16865 17153 16899 17187
rect 16899 17153 16908 17187
rect 16856 17144 16908 17153
rect 19340 17144 19392 17196
rect 22560 17144 22612 17196
rect 23848 17144 23900 17196
rect 25780 17144 25832 17196
rect 27712 17144 27764 17196
rect 29000 17144 29052 17196
rect 30932 17144 30984 17196
rect 32220 17144 32272 17196
rect 35072 17187 35124 17196
rect 35072 17153 35081 17187
rect 35081 17153 35115 17187
rect 35115 17153 35124 17187
rect 35072 17144 35124 17153
rect 35440 17144 35492 17196
rect 37372 17144 37424 17196
rect 42800 17187 42852 17196
rect 42800 17153 42809 17187
rect 42809 17153 42843 17187
rect 42843 17153 42852 17187
rect 42800 17144 42852 17153
rect 43444 17187 43496 17196
rect 43444 17153 43453 17187
rect 43453 17153 43487 17187
rect 43487 17153 43496 17187
rect 43444 17144 43496 17153
rect 43812 17144 43864 17196
rect 10876 17076 10928 17128
rect 32588 17119 32640 17128
rect 32588 17085 32597 17119
rect 32597 17085 32631 17119
rect 32631 17085 32640 17119
rect 32588 17076 32640 17085
rect 3608 17008 3660 17060
rect 15660 17008 15712 17060
rect 1768 16983 1820 16992
rect 1768 16949 1777 16983
rect 1777 16949 1811 16983
rect 1811 16949 1820 16983
rect 1768 16940 1820 16949
rect 2504 16983 2556 16992
rect 2504 16949 2513 16983
rect 2513 16949 2547 16983
rect 2547 16949 2556 16983
rect 2504 16940 2556 16949
rect 10232 16940 10284 16992
rect 16580 16940 16632 16992
rect 23756 16940 23808 16992
rect 31300 16940 31352 16992
rect 34520 16940 34572 16992
rect 38844 16940 38896 16992
rect 6423 16838 6475 16890
rect 6487 16838 6539 16890
rect 6551 16838 6603 16890
rect 6615 16838 6667 16890
rect 6679 16838 6731 16890
rect 17370 16838 17422 16890
rect 17434 16838 17486 16890
rect 17498 16838 17550 16890
rect 17562 16838 17614 16890
rect 17626 16838 17678 16890
rect 28317 16838 28369 16890
rect 28381 16838 28433 16890
rect 28445 16838 28497 16890
rect 28509 16838 28561 16890
rect 28573 16838 28625 16890
rect 39264 16838 39316 16890
rect 39328 16838 39380 16890
rect 39392 16838 39444 16890
rect 39456 16838 39508 16890
rect 39520 16838 39572 16890
rect 45100 16736 45152 16788
rect 5172 16600 5224 16652
rect 20 16532 72 16584
rect 7012 16575 7064 16584
rect 7012 16541 7021 16575
rect 7021 16541 7055 16575
rect 7055 16541 7064 16575
rect 7012 16532 7064 16541
rect 19524 16532 19576 16584
rect 20628 16532 20680 16584
rect 17224 16464 17276 16516
rect 11896 16294 11948 16346
rect 11960 16294 12012 16346
rect 12024 16294 12076 16346
rect 12088 16294 12140 16346
rect 12152 16294 12204 16346
rect 22843 16294 22895 16346
rect 22907 16294 22959 16346
rect 22971 16294 23023 16346
rect 23035 16294 23087 16346
rect 23099 16294 23151 16346
rect 33790 16294 33842 16346
rect 33854 16294 33906 16346
rect 33918 16294 33970 16346
rect 33982 16294 34034 16346
rect 34046 16294 34098 16346
rect 44737 16294 44789 16346
rect 44801 16294 44853 16346
rect 44865 16294 44917 16346
rect 44929 16294 44981 16346
rect 44993 16294 45045 16346
rect 1032 16056 1084 16108
rect 41604 16056 41656 16108
rect 35716 15988 35768 16040
rect 36176 16031 36228 16040
rect 36176 15997 36185 16031
rect 36185 15997 36219 16031
rect 36219 15997 36228 16031
rect 36176 15988 36228 15997
rect 40592 15988 40644 16040
rect 41512 15988 41564 16040
rect 36636 15852 36688 15904
rect 44364 15895 44416 15904
rect 44364 15861 44373 15895
rect 44373 15861 44407 15895
rect 44407 15861 44416 15895
rect 44364 15852 44416 15861
rect 6423 15750 6475 15802
rect 6487 15750 6539 15802
rect 6551 15750 6603 15802
rect 6615 15750 6667 15802
rect 6679 15750 6731 15802
rect 17370 15750 17422 15802
rect 17434 15750 17486 15802
rect 17498 15750 17550 15802
rect 17562 15750 17614 15802
rect 17626 15750 17678 15802
rect 28317 15750 28369 15802
rect 28381 15750 28433 15802
rect 28445 15750 28497 15802
rect 28509 15750 28561 15802
rect 28573 15750 28625 15802
rect 39264 15750 39316 15802
rect 39328 15750 39380 15802
rect 39392 15750 39444 15802
rect 39456 15750 39508 15802
rect 39520 15750 39572 15802
rect 19524 15691 19576 15700
rect 19524 15657 19533 15691
rect 19533 15657 19567 15691
rect 19567 15657 19576 15691
rect 19524 15648 19576 15657
rect 35716 15691 35768 15700
rect 35716 15657 35725 15691
rect 35725 15657 35759 15691
rect 35759 15657 35768 15691
rect 35716 15648 35768 15657
rect 10140 15487 10192 15496
rect 10140 15453 10149 15487
rect 10149 15453 10183 15487
rect 10183 15453 10192 15487
rect 10140 15444 10192 15453
rect 10232 15444 10284 15496
rect 17132 15444 17184 15496
rect 35900 15512 35952 15564
rect 43996 15555 44048 15564
rect 43996 15521 44005 15555
rect 44005 15521 44039 15555
rect 44039 15521 44048 15555
rect 43996 15512 44048 15521
rect 17776 15487 17828 15496
rect 17776 15453 17785 15487
rect 17785 15453 17819 15487
rect 17819 15453 17828 15487
rect 17776 15444 17828 15453
rect 25228 15487 25280 15496
rect 25228 15453 25237 15487
rect 25237 15453 25271 15487
rect 25271 15453 25280 15487
rect 25228 15444 25280 15453
rect 41420 15444 41472 15496
rect 19892 15419 19944 15428
rect 19892 15385 19901 15419
rect 19901 15385 19935 15419
rect 19935 15385 19944 15419
rect 19892 15376 19944 15385
rect 36268 15376 36320 15428
rect 12624 15351 12676 15360
rect 12624 15317 12633 15351
rect 12633 15317 12667 15351
rect 12667 15317 12676 15351
rect 12624 15308 12676 15317
rect 19800 15308 19852 15360
rect 19984 15351 20036 15360
rect 19984 15317 19993 15351
rect 19993 15317 20027 15351
rect 20027 15317 20036 15351
rect 19984 15308 20036 15317
rect 25136 15308 25188 15360
rect 36176 15351 36228 15360
rect 36176 15317 36185 15351
rect 36185 15317 36219 15351
rect 36219 15317 36228 15351
rect 36176 15308 36228 15317
rect 11896 15206 11948 15258
rect 11960 15206 12012 15258
rect 12024 15206 12076 15258
rect 12088 15206 12140 15258
rect 12152 15206 12204 15258
rect 22843 15206 22895 15258
rect 22907 15206 22959 15258
rect 22971 15206 23023 15258
rect 23035 15206 23087 15258
rect 23099 15206 23151 15258
rect 33790 15206 33842 15258
rect 33854 15206 33906 15258
rect 33918 15206 33970 15258
rect 33982 15206 34034 15258
rect 34046 15206 34098 15258
rect 44737 15206 44789 15258
rect 44801 15206 44853 15258
rect 44865 15206 44917 15258
rect 44929 15206 44981 15258
rect 44993 15206 45045 15258
rect 17776 15104 17828 15156
rect 19984 15104 20036 15156
rect 5632 14968 5684 15020
rect 7380 15011 7432 15020
rect 7380 14977 7389 15011
rect 7389 14977 7423 15011
rect 7423 14977 7432 15011
rect 7380 14968 7432 14977
rect 12624 14968 12676 15020
rect 13820 14968 13872 15020
rect 15200 15011 15252 15020
rect 15200 14977 15234 15011
rect 15234 14977 15252 15011
rect 15200 14968 15252 14977
rect 19708 15036 19760 15088
rect 17224 14968 17276 15020
rect 17868 14968 17920 15020
rect 19800 14968 19852 15020
rect 22100 14968 22152 15020
rect 24860 15011 24912 15020
rect 24860 14977 24869 15011
rect 24869 14977 24903 15011
rect 24903 14977 24912 15011
rect 24860 14968 24912 14977
rect 25136 15011 25188 15020
rect 25136 14977 25170 15011
rect 25170 14977 25188 15011
rect 25136 14968 25188 14977
rect 27712 14968 27764 15020
rect 30196 14968 30248 15020
rect 31392 15011 31444 15020
rect 31392 14977 31401 15011
rect 31401 14977 31435 15011
rect 31435 14977 31444 15011
rect 31392 14968 31444 14977
rect 32036 15036 32088 15088
rect 32588 15104 32640 15156
rect 6828 14764 6880 14816
rect 7196 14807 7248 14816
rect 7196 14773 7205 14807
rect 7205 14773 7239 14807
rect 7239 14773 7248 14807
rect 7196 14764 7248 14773
rect 22376 14764 22428 14816
rect 24400 14807 24452 14816
rect 24400 14773 24409 14807
rect 24409 14773 24443 14807
rect 24443 14773 24452 14807
rect 24400 14764 24452 14773
rect 26608 14764 26660 14816
rect 29552 14900 29604 14952
rect 29644 14832 29696 14884
rect 33600 14968 33652 15020
rect 36636 15011 36688 15020
rect 36636 14977 36645 15011
rect 36645 14977 36679 15011
rect 36679 14977 36688 15011
rect 36636 14968 36688 14977
rect 40132 14968 40184 15020
rect 34520 14900 34572 14952
rect 34612 14943 34664 14952
rect 34612 14909 34621 14943
rect 34621 14909 34655 14943
rect 34655 14909 34664 14943
rect 34612 14900 34664 14909
rect 38936 14900 38988 14952
rect 28908 14764 28960 14816
rect 30012 14764 30064 14816
rect 31116 14764 31168 14816
rect 31208 14807 31260 14816
rect 31208 14773 31217 14807
rect 31217 14773 31251 14807
rect 31251 14773 31260 14807
rect 31208 14764 31260 14773
rect 36176 14832 36228 14884
rect 37096 14832 37148 14884
rect 36268 14764 36320 14816
rect 36452 14807 36504 14816
rect 36452 14773 36461 14807
rect 36461 14773 36495 14807
rect 36495 14773 36504 14807
rect 36452 14764 36504 14773
rect 39672 14764 39724 14816
rect 6423 14662 6475 14714
rect 6487 14662 6539 14714
rect 6551 14662 6603 14714
rect 6615 14662 6667 14714
rect 6679 14662 6731 14714
rect 17370 14662 17422 14714
rect 17434 14662 17486 14714
rect 17498 14662 17550 14714
rect 17562 14662 17614 14714
rect 17626 14662 17678 14714
rect 28317 14662 28369 14714
rect 28381 14662 28433 14714
rect 28445 14662 28497 14714
rect 28509 14662 28561 14714
rect 28573 14662 28625 14714
rect 39264 14662 39316 14714
rect 39328 14662 39380 14714
rect 39392 14662 39444 14714
rect 39456 14662 39508 14714
rect 39520 14662 39572 14714
rect 5632 14603 5684 14612
rect 5632 14569 5641 14603
rect 5641 14569 5675 14603
rect 5675 14569 5684 14603
rect 5632 14560 5684 14569
rect 5816 14560 5868 14612
rect 7840 14560 7892 14612
rect 17224 14560 17276 14612
rect 4712 14399 4764 14408
rect 4712 14365 4721 14399
rect 4721 14365 4755 14399
rect 4755 14365 4764 14399
rect 4712 14356 4764 14365
rect 4344 14288 4396 14340
rect 5632 14399 5684 14408
rect 5632 14365 5641 14399
rect 5641 14365 5675 14399
rect 5675 14365 5684 14399
rect 5632 14356 5684 14365
rect 5724 14356 5776 14408
rect 10140 14424 10192 14476
rect 6552 14356 6604 14408
rect 7196 14356 7248 14408
rect 12256 14356 12308 14408
rect 14280 14399 14332 14408
rect 14280 14365 14289 14399
rect 14289 14365 14323 14399
rect 14323 14365 14332 14399
rect 14280 14356 14332 14365
rect 14464 14399 14516 14408
rect 14464 14365 14473 14399
rect 14473 14365 14507 14399
rect 14507 14365 14516 14399
rect 14464 14356 14516 14365
rect 15660 14399 15712 14408
rect 15660 14365 15669 14399
rect 15669 14365 15703 14399
rect 15703 14365 15712 14399
rect 15660 14356 15712 14365
rect 4160 14220 4212 14272
rect 8208 14220 8260 14272
rect 8484 14263 8536 14272
rect 8484 14229 8493 14263
rect 8493 14229 8527 14263
rect 8527 14229 8536 14263
rect 8484 14220 8536 14229
rect 11336 14220 11388 14272
rect 15292 14288 15344 14340
rect 15476 14288 15528 14340
rect 19892 14492 19944 14544
rect 25228 14560 25280 14612
rect 19984 14424 20036 14476
rect 20996 14424 21048 14476
rect 23756 14467 23808 14476
rect 23756 14433 23765 14467
rect 23765 14433 23799 14467
rect 23799 14433 23808 14467
rect 23756 14424 23808 14433
rect 23848 14467 23900 14476
rect 23848 14433 23857 14467
rect 23857 14433 23891 14467
rect 23891 14433 23900 14467
rect 23848 14424 23900 14433
rect 25504 14424 25556 14476
rect 29644 14560 29696 14612
rect 31392 14560 31444 14612
rect 33600 14603 33652 14612
rect 33600 14569 33609 14603
rect 33609 14569 33643 14603
rect 33643 14569 33652 14603
rect 33600 14560 33652 14569
rect 26792 14467 26844 14476
rect 26792 14433 26801 14467
rect 26801 14433 26835 14467
rect 26835 14433 26844 14467
rect 26792 14424 26844 14433
rect 41604 14560 41656 14612
rect 36268 14535 36320 14544
rect 36268 14501 36277 14535
rect 36277 14501 36311 14535
rect 36311 14501 36320 14535
rect 36268 14492 36320 14501
rect 12348 14220 12400 14272
rect 13544 14220 13596 14272
rect 15660 14220 15712 14272
rect 19708 14356 19760 14408
rect 22192 14356 22244 14408
rect 20628 14288 20680 14340
rect 23664 14331 23716 14340
rect 23664 14297 23673 14331
rect 23673 14297 23707 14331
rect 23707 14297 23716 14331
rect 23664 14288 23716 14297
rect 24400 14356 24452 14408
rect 26608 14399 26660 14408
rect 26608 14365 26617 14399
rect 26617 14365 26651 14399
rect 26651 14365 26660 14399
rect 26608 14356 26660 14365
rect 27804 14399 27856 14408
rect 27804 14365 27813 14399
rect 27813 14365 27847 14399
rect 27847 14365 27856 14399
rect 27804 14356 27856 14365
rect 28908 14356 28960 14408
rect 29736 14399 29788 14408
rect 29736 14365 29745 14399
rect 29745 14365 29779 14399
rect 29779 14365 29788 14399
rect 29736 14356 29788 14365
rect 30932 14356 30984 14408
rect 31116 14356 31168 14408
rect 32404 14356 32456 14408
rect 35900 14424 35952 14476
rect 38200 14424 38252 14476
rect 18512 14263 18564 14272
rect 18512 14229 18521 14263
rect 18521 14229 18555 14263
rect 18555 14229 18564 14263
rect 18512 14220 18564 14229
rect 19892 14263 19944 14272
rect 19892 14229 19901 14263
rect 19901 14229 19935 14263
rect 19935 14229 19944 14263
rect 19892 14220 19944 14229
rect 21916 14263 21968 14272
rect 21916 14229 21925 14263
rect 21925 14229 21959 14263
rect 21959 14229 21968 14263
rect 21916 14220 21968 14229
rect 23572 14220 23624 14272
rect 26792 14220 26844 14272
rect 31116 14220 31168 14272
rect 34612 14356 34664 14408
rect 36360 14356 36412 14408
rect 37096 14399 37148 14408
rect 37096 14365 37105 14399
rect 37105 14365 37139 14399
rect 37139 14365 37148 14399
rect 37096 14356 37148 14365
rect 39672 14356 39724 14408
rect 40040 14399 40092 14408
rect 40040 14365 40049 14399
rect 40049 14365 40083 14399
rect 40083 14365 40092 14399
rect 40040 14356 40092 14365
rect 41696 14356 41748 14408
rect 36452 14288 36504 14340
rect 36084 14220 36136 14272
rect 36268 14220 36320 14272
rect 37832 14220 37884 14272
rect 45008 14288 45060 14340
rect 11896 14118 11948 14170
rect 11960 14118 12012 14170
rect 12024 14118 12076 14170
rect 12088 14118 12140 14170
rect 12152 14118 12204 14170
rect 22843 14118 22895 14170
rect 22907 14118 22959 14170
rect 22971 14118 23023 14170
rect 23035 14118 23087 14170
rect 23099 14118 23151 14170
rect 33790 14118 33842 14170
rect 33854 14118 33906 14170
rect 33918 14118 33970 14170
rect 33982 14118 34034 14170
rect 34046 14118 34098 14170
rect 44737 14118 44789 14170
rect 44801 14118 44853 14170
rect 44865 14118 44917 14170
rect 44929 14118 44981 14170
rect 44993 14118 45045 14170
rect 4712 14016 4764 14068
rect 5632 14016 5684 14068
rect 7840 14016 7892 14068
rect 9772 14016 9824 14068
rect 12256 14059 12308 14068
rect 12256 14025 12265 14059
rect 12265 14025 12299 14059
rect 12299 14025 12308 14059
rect 12256 14016 12308 14025
rect 14280 14016 14332 14068
rect 5540 13948 5592 14000
rect 6828 13991 6880 14000
rect 6828 13957 6862 13991
rect 6862 13957 6880 13991
rect 6828 13948 6880 13957
rect 8208 13948 8260 14000
rect 11244 13948 11296 14000
rect 1032 13880 1084 13932
rect 940 13812 992 13864
rect 3056 13923 3108 13932
rect 3056 13889 3065 13923
rect 3065 13889 3099 13923
rect 3099 13889 3108 13923
rect 3056 13880 3108 13889
rect 4988 13923 5040 13932
rect 4988 13889 4997 13923
rect 4997 13889 5031 13923
rect 5031 13889 5040 13923
rect 4988 13880 5040 13889
rect 5816 13880 5868 13932
rect 6552 13923 6604 13932
rect 6552 13889 6561 13923
rect 6561 13889 6595 13923
rect 6595 13889 6604 13923
rect 6552 13880 6604 13889
rect 5264 13855 5316 13864
rect 5264 13821 5273 13855
rect 5273 13821 5307 13855
rect 5307 13821 5316 13855
rect 5264 13812 5316 13821
rect 7104 13880 7156 13932
rect 8484 13880 8536 13932
rect 9404 13880 9456 13932
rect 11152 13923 11204 13932
rect 11152 13889 11161 13923
rect 11161 13889 11195 13923
rect 11195 13889 11204 13923
rect 11152 13880 11204 13889
rect 5724 13744 5776 13796
rect 11336 13812 11388 13864
rect 13636 13880 13688 13932
rect 19892 14059 19944 14068
rect 19892 14025 19901 14059
rect 19901 14025 19935 14059
rect 19935 14025 19944 14059
rect 19892 14016 19944 14025
rect 26608 14016 26660 14068
rect 30196 14059 30248 14068
rect 30196 14025 30205 14059
rect 30205 14025 30239 14059
rect 30239 14025 30248 14059
rect 30196 14016 30248 14025
rect 31392 14016 31444 14068
rect 37832 14059 37884 14068
rect 37832 14025 37841 14059
rect 37841 14025 37875 14059
rect 37875 14025 37884 14059
rect 37832 14016 37884 14025
rect 40132 14059 40184 14068
rect 40132 14025 40141 14059
rect 40141 14025 40175 14059
rect 40175 14025 40184 14059
rect 40132 14016 40184 14025
rect 41420 14016 41472 14068
rect 21916 13948 21968 14000
rect 25504 13948 25556 14000
rect 15108 13880 15160 13932
rect 15568 13923 15620 13932
rect 15568 13889 15577 13923
rect 15577 13889 15611 13923
rect 15611 13889 15620 13923
rect 15568 13880 15620 13889
rect 19340 13880 19392 13932
rect 22100 13880 22152 13932
rect 23848 13880 23900 13932
rect 29552 13880 29604 13932
rect 30012 13923 30064 13932
rect 30012 13889 30021 13923
rect 30021 13889 30055 13923
rect 30055 13889 30064 13923
rect 30012 13880 30064 13889
rect 12624 13812 12676 13864
rect 17868 13812 17920 13864
rect 20996 13855 21048 13864
rect 20996 13821 21005 13855
rect 21005 13821 21039 13855
rect 21039 13821 21048 13855
rect 20996 13812 21048 13821
rect 6000 13676 6052 13728
rect 8760 13719 8812 13728
rect 8760 13685 8769 13719
rect 8769 13685 8803 13719
rect 8803 13685 8812 13719
rect 8760 13676 8812 13685
rect 12716 13676 12768 13728
rect 20352 13719 20404 13728
rect 20352 13685 20361 13719
rect 20361 13685 20395 13719
rect 20395 13685 20404 13719
rect 20352 13676 20404 13685
rect 23020 13812 23072 13864
rect 24860 13812 24912 13864
rect 26148 13812 26200 13864
rect 27804 13812 27856 13864
rect 29000 13812 29052 13864
rect 29736 13812 29788 13864
rect 31208 13948 31260 14000
rect 30288 13880 30340 13932
rect 32404 13812 32456 13864
rect 34612 13948 34664 14000
rect 26792 13744 26844 13796
rect 38384 13880 38436 13932
rect 40040 13948 40092 14000
rect 41696 13991 41748 14000
rect 41696 13957 41705 13991
rect 41705 13957 41739 13991
rect 41739 13957 41748 13991
rect 41696 13948 41748 13957
rect 38844 13880 38896 13932
rect 36268 13812 36320 13864
rect 36452 13855 36504 13864
rect 36452 13821 36461 13855
rect 36461 13821 36495 13855
rect 36495 13821 36504 13855
rect 36452 13812 36504 13821
rect 37924 13855 37976 13864
rect 37924 13821 37933 13855
rect 37933 13821 37967 13855
rect 37967 13821 37976 13855
rect 37924 13812 37976 13821
rect 38200 13812 38252 13864
rect 41788 13855 41840 13864
rect 41788 13821 41797 13855
rect 41797 13821 41831 13855
rect 41831 13821 41840 13855
rect 41788 13812 41840 13821
rect 36636 13676 36688 13728
rect 38936 13676 38988 13728
rect 41972 13744 42024 13796
rect 6423 13574 6475 13626
rect 6487 13574 6539 13626
rect 6551 13574 6603 13626
rect 6615 13574 6667 13626
rect 6679 13574 6731 13626
rect 17370 13574 17422 13626
rect 17434 13574 17486 13626
rect 17498 13574 17550 13626
rect 17562 13574 17614 13626
rect 17626 13574 17678 13626
rect 28317 13574 28369 13626
rect 28381 13574 28433 13626
rect 28445 13574 28497 13626
rect 28509 13574 28561 13626
rect 28573 13574 28625 13626
rect 39264 13574 39316 13626
rect 39328 13574 39380 13626
rect 39392 13574 39444 13626
rect 39456 13574 39508 13626
rect 39520 13574 39572 13626
rect 4160 13472 4212 13524
rect 4988 13472 5040 13524
rect 6828 13472 6880 13524
rect 8760 13472 8812 13524
rect 11060 13472 11112 13524
rect 12624 13472 12676 13524
rect 15568 13472 15620 13524
rect 18512 13472 18564 13524
rect 19340 13472 19392 13524
rect 22192 13472 22244 13524
rect 7380 13404 7432 13456
rect 11244 13447 11296 13456
rect 11244 13413 11253 13447
rect 11253 13413 11287 13447
rect 11287 13413 11296 13447
rect 11244 13404 11296 13413
rect 4068 13268 4120 13320
rect 11152 13336 11204 13388
rect 12348 13404 12400 13456
rect 25504 13472 25556 13524
rect 36360 13472 36412 13524
rect 5816 13243 5868 13252
rect 5816 13209 5825 13243
rect 5825 13209 5859 13243
rect 5859 13209 5868 13243
rect 5816 13200 5868 13209
rect 6000 13243 6052 13252
rect 6000 13209 6025 13243
rect 6025 13209 6052 13243
rect 6000 13200 6052 13209
rect 7104 13200 7156 13252
rect 8208 13268 8260 13320
rect 11336 13268 11388 13320
rect 11520 13336 11572 13388
rect 19984 13379 20036 13388
rect 19984 13345 19993 13379
rect 19993 13345 20027 13379
rect 20027 13345 20036 13379
rect 19984 13336 20036 13345
rect 24676 13336 24728 13388
rect 12716 13268 12768 13320
rect 12808 13311 12860 13320
rect 12808 13277 12817 13311
rect 12817 13277 12851 13311
rect 12851 13277 12860 13311
rect 12808 13268 12860 13277
rect 8484 13200 8536 13252
rect 12532 13243 12584 13252
rect 12532 13209 12541 13243
rect 12541 13209 12575 13243
rect 12575 13209 12584 13243
rect 12532 13200 12584 13209
rect 4344 13132 4396 13184
rect 6552 13132 6604 13184
rect 13084 13200 13136 13252
rect 14280 13311 14332 13320
rect 14280 13277 14289 13311
rect 14289 13277 14323 13311
rect 14323 13277 14332 13311
rect 14280 13268 14332 13277
rect 14464 13311 14516 13320
rect 14464 13277 14473 13311
rect 14473 13277 14507 13311
rect 14507 13277 14516 13311
rect 14464 13268 14516 13277
rect 20352 13268 20404 13320
rect 23020 13268 23072 13320
rect 23572 13268 23624 13320
rect 24860 13268 24912 13320
rect 27896 13311 27948 13320
rect 15108 13243 15160 13252
rect 15108 13209 15117 13243
rect 15117 13209 15151 13243
rect 15151 13209 15160 13243
rect 15108 13200 15160 13209
rect 15292 13243 15344 13252
rect 15292 13209 15317 13243
rect 15317 13209 15344 13243
rect 15292 13200 15344 13209
rect 17776 13243 17828 13252
rect 17776 13209 17810 13243
rect 17810 13209 17828 13243
rect 17776 13200 17828 13209
rect 17868 13200 17920 13252
rect 27896 13277 27905 13311
rect 27905 13277 27939 13311
rect 27939 13277 27948 13311
rect 27896 13268 27948 13277
rect 28172 13311 28224 13320
rect 28172 13277 28181 13311
rect 28181 13277 28215 13311
rect 28215 13277 28224 13311
rect 28172 13268 28224 13277
rect 28908 13268 28960 13320
rect 30840 13268 30892 13320
rect 32772 13311 32824 13320
rect 32772 13277 32781 13311
rect 32781 13277 32815 13311
rect 32815 13277 32824 13311
rect 32772 13268 32824 13277
rect 37832 13472 37884 13524
rect 38384 13404 38436 13456
rect 36636 13311 36688 13320
rect 36636 13277 36659 13311
rect 36659 13277 36688 13311
rect 36636 13268 36688 13277
rect 12992 13175 13044 13184
rect 12992 13141 13001 13175
rect 13001 13141 13035 13175
rect 13035 13141 13044 13175
rect 12992 13132 13044 13141
rect 18880 13132 18932 13184
rect 22008 13175 22060 13184
rect 22008 13141 22017 13175
rect 22017 13141 22051 13175
rect 22051 13141 22060 13175
rect 22008 13132 22060 13141
rect 22652 13132 22704 13184
rect 28080 13175 28132 13184
rect 28080 13141 28089 13175
rect 28089 13141 28123 13175
rect 28123 13141 28132 13175
rect 28080 13132 28132 13141
rect 28264 13132 28316 13184
rect 31484 13132 31536 13184
rect 37096 13200 37148 13252
rect 38108 13132 38160 13184
rect 11896 13030 11948 13082
rect 11960 13030 12012 13082
rect 12024 13030 12076 13082
rect 12088 13030 12140 13082
rect 12152 13030 12204 13082
rect 22843 13030 22895 13082
rect 22907 13030 22959 13082
rect 22971 13030 23023 13082
rect 23035 13030 23087 13082
rect 23099 13030 23151 13082
rect 33790 13030 33842 13082
rect 33854 13030 33906 13082
rect 33918 13030 33970 13082
rect 33982 13030 34034 13082
rect 34046 13030 34098 13082
rect 44737 13030 44789 13082
rect 44801 13030 44853 13082
rect 44865 13030 44917 13082
rect 44929 13030 44981 13082
rect 44993 13030 45045 13082
rect 3056 12928 3108 12980
rect 4528 12971 4580 12980
rect 4528 12937 4537 12971
rect 4537 12937 4571 12971
rect 4571 12937 4580 12971
rect 4528 12928 4580 12937
rect 5724 12928 5776 12980
rect 11060 12971 11112 12980
rect 11060 12937 11069 12971
rect 11069 12937 11103 12971
rect 11103 12937 11112 12971
rect 11060 12928 11112 12937
rect 4896 12860 4948 12912
rect 5264 12860 5316 12912
rect 11336 12860 11388 12912
rect 12808 12928 12860 12980
rect 14464 12928 14516 12980
rect 18880 12971 18932 12980
rect 18880 12937 18889 12971
rect 18889 12937 18923 12971
rect 18923 12937 18932 12971
rect 18880 12928 18932 12937
rect 12440 12860 12492 12912
rect 3424 12792 3476 12844
rect 4344 12835 4396 12844
rect 4344 12801 4353 12835
rect 4353 12801 4387 12835
rect 4387 12801 4396 12835
rect 4344 12792 4396 12801
rect 4436 12724 4488 12776
rect 6552 12835 6604 12844
rect 6552 12801 6561 12835
rect 6561 12801 6595 12835
rect 6595 12801 6604 12835
rect 6552 12792 6604 12801
rect 5724 12588 5776 12640
rect 5816 12631 5868 12640
rect 5816 12597 5825 12631
rect 5825 12597 5859 12631
rect 5859 12597 5868 12631
rect 5816 12588 5868 12597
rect 6828 12792 6880 12844
rect 9404 12835 9456 12844
rect 9404 12801 9413 12835
rect 9413 12801 9447 12835
rect 9447 12801 9456 12835
rect 9404 12792 9456 12801
rect 11060 12792 11112 12844
rect 11152 12835 11204 12844
rect 11152 12801 11161 12835
rect 11161 12801 11195 12835
rect 11195 12801 11204 12835
rect 11152 12792 11204 12801
rect 11244 12792 11296 12844
rect 12348 12835 12400 12844
rect 13728 12860 13780 12912
rect 12348 12801 12362 12835
rect 12362 12801 12396 12835
rect 12396 12801 12400 12835
rect 12348 12792 12400 12801
rect 13084 12792 13136 12844
rect 14280 12792 14332 12844
rect 17868 12860 17920 12912
rect 18052 12792 18104 12844
rect 20720 12860 20772 12912
rect 19432 12792 19484 12844
rect 22744 12835 22796 12844
rect 22744 12801 22753 12835
rect 22753 12801 22787 12835
rect 22787 12801 22796 12835
rect 22744 12792 22796 12801
rect 24860 12928 24912 12980
rect 24584 12792 24636 12844
rect 10784 12656 10836 12708
rect 22008 12656 22060 12708
rect 27160 12835 27212 12844
rect 27160 12801 27169 12835
rect 27169 12801 27203 12835
rect 27203 12801 27212 12835
rect 27160 12792 27212 12801
rect 28908 12928 28960 12980
rect 28264 12903 28316 12912
rect 28264 12869 28273 12903
rect 28273 12869 28307 12903
rect 28307 12869 28316 12903
rect 28264 12860 28316 12869
rect 31484 12971 31536 12980
rect 31484 12937 31493 12971
rect 31493 12937 31527 12971
rect 31527 12937 31536 12971
rect 31484 12928 31536 12937
rect 38200 12928 38252 12980
rect 32036 12860 32088 12912
rect 30380 12835 30432 12844
rect 30380 12801 30389 12835
rect 30389 12801 30423 12835
rect 30423 12801 30432 12835
rect 30380 12792 30432 12801
rect 31208 12792 31260 12844
rect 31484 12724 31536 12776
rect 32312 12767 32364 12776
rect 32312 12733 32321 12767
rect 32321 12733 32355 12767
rect 32355 12733 32364 12767
rect 32312 12724 32364 12733
rect 6920 12588 6972 12640
rect 14832 12588 14884 12640
rect 24952 12631 25004 12640
rect 24952 12597 24961 12631
rect 24961 12597 24995 12631
rect 24995 12597 25004 12631
rect 24952 12588 25004 12597
rect 26884 12588 26936 12640
rect 28080 12588 28132 12640
rect 31024 12631 31076 12640
rect 31024 12597 31033 12631
rect 31033 12597 31067 12631
rect 31067 12597 31076 12631
rect 31024 12588 31076 12597
rect 31484 12588 31536 12640
rect 38936 12860 38988 12912
rect 40040 12860 40092 12912
rect 33324 12835 33376 12844
rect 33324 12801 33333 12835
rect 33333 12801 33367 12835
rect 33367 12801 33376 12835
rect 33324 12792 33376 12801
rect 36084 12835 36136 12844
rect 36084 12801 36093 12835
rect 36093 12801 36127 12835
rect 36127 12801 36136 12835
rect 36084 12792 36136 12801
rect 37648 12835 37700 12844
rect 37648 12801 37657 12835
rect 37657 12801 37691 12835
rect 37691 12801 37700 12835
rect 37648 12792 37700 12801
rect 38384 12835 38436 12844
rect 38384 12801 38393 12835
rect 38393 12801 38427 12835
rect 38427 12801 38436 12835
rect 38384 12792 38436 12801
rect 41052 12835 41104 12844
rect 41052 12801 41061 12835
rect 41061 12801 41095 12835
rect 41095 12801 41104 12835
rect 41052 12792 41104 12801
rect 38660 12767 38712 12776
rect 38660 12733 38669 12767
rect 38669 12733 38703 12767
rect 38703 12733 38712 12767
rect 38660 12724 38712 12733
rect 34336 12656 34388 12708
rect 33140 12631 33192 12640
rect 33140 12597 33149 12631
rect 33149 12597 33183 12631
rect 33183 12597 33192 12631
rect 33140 12588 33192 12597
rect 36544 12588 36596 12640
rect 37464 12631 37516 12640
rect 37464 12597 37473 12631
rect 37473 12597 37507 12631
rect 37507 12597 37516 12631
rect 37464 12588 37516 12597
rect 40960 12588 41012 12640
rect 45008 12588 45060 12640
rect 6423 12486 6475 12538
rect 6487 12486 6539 12538
rect 6551 12486 6603 12538
rect 6615 12486 6667 12538
rect 6679 12486 6731 12538
rect 17370 12486 17422 12538
rect 17434 12486 17486 12538
rect 17498 12486 17550 12538
rect 17562 12486 17614 12538
rect 17626 12486 17678 12538
rect 28317 12486 28369 12538
rect 28381 12486 28433 12538
rect 28445 12486 28497 12538
rect 28509 12486 28561 12538
rect 28573 12486 28625 12538
rect 39264 12486 39316 12538
rect 39328 12486 39380 12538
rect 39392 12486 39444 12538
rect 39456 12486 39508 12538
rect 39520 12486 39572 12538
rect 6920 12427 6972 12436
rect 6920 12393 6929 12427
rect 6929 12393 6963 12427
rect 6963 12393 6972 12427
rect 6920 12384 6972 12393
rect 11520 12384 11572 12436
rect 12532 12384 12584 12436
rect 12992 12384 13044 12436
rect 13360 12384 13412 12436
rect 15108 12384 15160 12436
rect 17776 12384 17828 12436
rect 20628 12384 20680 12436
rect 22468 12384 22520 12436
rect 22744 12384 22796 12436
rect 24584 12427 24636 12436
rect 24584 12393 24593 12427
rect 24593 12393 24627 12427
rect 24627 12393 24636 12427
rect 24584 12384 24636 12393
rect 4528 12316 4580 12368
rect 14832 12359 14884 12368
rect 4068 12248 4120 12300
rect 9864 12291 9916 12300
rect 9864 12257 9873 12291
rect 9873 12257 9907 12291
rect 9907 12257 9916 12291
rect 9864 12248 9916 12257
rect 10784 12291 10836 12300
rect 10784 12257 10793 12291
rect 10793 12257 10827 12291
rect 10827 12257 10836 12291
rect 10784 12248 10836 12257
rect 10968 12248 11020 12300
rect 4344 12180 4396 12232
rect 4896 12180 4948 12232
rect 4988 12223 5040 12232
rect 4988 12189 4997 12223
rect 4997 12189 5031 12223
rect 5031 12189 5040 12223
rect 4988 12180 5040 12189
rect 3884 12044 3936 12096
rect 5540 12223 5592 12232
rect 5540 12189 5549 12223
rect 5549 12189 5583 12223
rect 5583 12189 5592 12223
rect 5540 12180 5592 12189
rect 5724 12112 5776 12164
rect 6920 12180 6972 12232
rect 9772 12223 9824 12232
rect 9772 12189 9781 12223
rect 9781 12189 9815 12223
rect 9815 12189 9824 12223
rect 9772 12180 9824 12189
rect 11336 12180 11388 12232
rect 11428 12180 11480 12232
rect 14832 12325 14841 12359
rect 14841 12325 14875 12359
rect 14875 12325 14884 12359
rect 14832 12316 14884 12325
rect 27896 12427 27948 12436
rect 27896 12393 27905 12427
rect 27905 12393 27939 12427
rect 27939 12393 27948 12427
rect 27896 12384 27948 12393
rect 28080 12384 28132 12436
rect 28264 12384 28316 12436
rect 28724 12384 28776 12436
rect 30288 12427 30340 12436
rect 30288 12393 30297 12427
rect 30297 12393 30331 12427
rect 30331 12393 30340 12427
rect 30288 12384 30340 12393
rect 33324 12384 33376 12436
rect 38660 12384 38712 12436
rect 40040 12427 40092 12436
rect 40040 12393 40049 12427
rect 40049 12393 40083 12427
rect 40083 12393 40092 12427
rect 40040 12384 40092 12393
rect 28356 12316 28408 12368
rect 28540 12316 28592 12368
rect 13452 12248 13504 12300
rect 5908 12112 5960 12164
rect 11152 12155 11204 12164
rect 11152 12121 11161 12155
rect 11161 12121 11195 12155
rect 11195 12121 11204 12155
rect 11152 12112 11204 12121
rect 7748 12087 7800 12096
rect 7748 12053 7757 12087
rect 7757 12053 7791 12087
rect 7791 12053 7800 12087
rect 7748 12044 7800 12053
rect 11060 12044 11112 12096
rect 11520 12112 11572 12164
rect 12624 12180 12676 12232
rect 12716 12180 12768 12232
rect 12256 12112 12308 12164
rect 11796 12044 11848 12096
rect 13360 12044 13412 12096
rect 13636 12180 13688 12232
rect 23848 12291 23900 12300
rect 23848 12257 23857 12291
rect 23857 12257 23891 12291
rect 23891 12257 23900 12291
rect 23848 12248 23900 12257
rect 16948 12180 17000 12232
rect 17776 12180 17828 12232
rect 21364 12180 21416 12232
rect 21456 12223 21508 12232
rect 21456 12189 21465 12223
rect 21465 12189 21499 12223
rect 21499 12189 21508 12223
rect 21456 12180 21508 12189
rect 26148 12291 26200 12300
rect 26148 12257 26157 12291
rect 26157 12257 26191 12291
rect 26191 12257 26200 12291
rect 26148 12248 26200 12257
rect 27436 12248 27488 12300
rect 25228 12223 25280 12232
rect 25228 12189 25237 12223
rect 25237 12189 25271 12223
rect 25271 12189 25280 12223
rect 25228 12180 25280 12189
rect 14464 12087 14516 12096
rect 14464 12053 14473 12087
rect 14473 12053 14507 12087
rect 14507 12053 14516 12087
rect 14464 12044 14516 12053
rect 19524 12044 19576 12096
rect 20996 12044 21048 12096
rect 22100 12044 22152 12096
rect 24952 12044 25004 12096
rect 26424 12155 26476 12164
rect 26424 12121 26433 12155
rect 26433 12121 26467 12155
rect 26467 12121 26476 12155
rect 26424 12112 26476 12121
rect 26884 12112 26936 12164
rect 28540 12223 28592 12232
rect 28540 12189 28549 12223
rect 28549 12189 28583 12223
rect 28583 12189 28592 12223
rect 28540 12180 28592 12189
rect 28632 12223 28684 12232
rect 28632 12189 28641 12223
rect 28641 12189 28675 12223
rect 28675 12189 28684 12223
rect 28632 12180 28684 12189
rect 30564 12248 30616 12300
rect 30472 12223 30524 12232
rect 30472 12189 30481 12223
rect 30481 12189 30515 12223
rect 30515 12189 30524 12223
rect 30472 12180 30524 12189
rect 31852 12248 31904 12300
rect 38200 12248 38252 12300
rect 41512 12291 41564 12300
rect 41512 12257 41521 12291
rect 41521 12257 41555 12291
rect 41555 12257 41564 12291
rect 41512 12248 41564 12257
rect 28908 12112 28960 12164
rect 30932 12180 30984 12232
rect 33600 12223 33652 12232
rect 33600 12189 33609 12223
rect 33609 12189 33643 12223
rect 33643 12189 33652 12223
rect 33600 12180 33652 12189
rect 34336 12223 34388 12232
rect 34336 12189 34345 12223
rect 34345 12189 34379 12223
rect 34379 12189 34388 12223
rect 34336 12180 34388 12189
rect 34888 12223 34940 12232
rect 34888 12189 34897 12223
rect 34897 12189 34931 12223
rect 34931 12189 34940 12223
rect 34888 12180 34940 12189
rect 40224 12223 40276 12232
rect 40224 12189 40233 12223
rect 40233 12189 40267 12223
rect 40267 12189 40276 12223
rect 40224 12180 40276 12189
rect 41420 12180 41472 12232
rect 28632 12044 28684 12096
rect 31392 12112 31444 12164
rect 33140 12112 33192 12164
rect 32496 12044 32548 12096
rect 36544 12112 36596 12164
rect 37464 12155 37516 12164
rect 37464 12121 37473 12155
rect 37473 12121 37507 12155
rect 37507 12121 37516 12155
rect 37464 12112 37516 12121
rect 38108 12112 38160 12164
rect 36636 12087 36688 12096
rect 36636 12053 36645 12087
rect 36645 12053 36679 12087
rect 36679 12053 36688 12087
rect 36636 12044 36688 12053
rect 39120 12044 39172 12096
rect 11896 11942 11948 11994
rect 11960 11942 12012 11994
rect 12024 11942 12076 11994
rect 12088 11942 12140 11994
rect 12152 11942 12204 11994
rect 22843 11942 22895 11994
rect 22907 11942 22959 11994
rect 22971 11942 23023 11994
rect 23035 11942 23087 11994
rect 23099 11942 23151 11994
rect 33790 11942 33842 11994
rect 33854 11942 33906 11994
rect 33918 11942 33970 11994
rect 33982 11942 34034 11994
rect 34046 11942 34098 11994
rect 44737 11942 44789 11994
rect 44801 11942 44853 11994
rect 44865 11942 44917 11994
rect 44929 11942 44981 11994
rect 44993 11942 45045 11994
rect 4068 11840 4120 11892
rect 4988 11840 5040 11892
rect 11244 11840 11296 11892
rect 12716 11883 12768 11892
rect 12716 11849 12725 11883
rect 12725 11849 12759 11883
rect 12759 11849 12768 11883
rect 12716 11840 12768 11849
rect 14464 11840 14516 11892
rect 18052 11883 18104 11892
rect 18052 11849 18061 11883
rect 18061 11849 18095 11883
rect 18095 11849 18104 11883
rect 18052 11840 18104 11849
rect 19432 11840 19484 11892
rect 19524 11840 19576 11892
rect 20904 11840 20956 11892
rect 21088 11883 21140 11892
rect 21088 11849 21097 11883
rect 21097 11849 21131 11883
rect 21131 11849 21140 11883
rect 21088 11840 21140 11849
rect 21364 11840 21416 11892
rect 22468 11883 22520 11892
rect 22468 11849 22477 11883
rect 22477 11849 22511 11883
rect 22511 11849 22520 11883
rect 22468 11840 22520 11849
rect 26424 11883 26476 11892
rect 26424 11849 26433 11883
rect 26433 11849 26467 11883
rect 26467 11849 26476 11883
rect 26424 11840 26476 11849
rect 2136 11747 2188 11756
rect 2136 11713 2145 11747
rect 2145 11713 2179 11747
rect 2179 11713 2188 11747
rect 2136 11704 2188 11713
rect 3332 11704 3384 11756
rect 3884 11704 3936 11756
rect 4344 11704 4396 11756
rect 5908 11772 5960 11824
rect 16948 11772 17000 11824
rect 23848 11772 23900 11824
rect 24952 11772 25004 11824
rect 2780 11679 2832 11688
rect 2780 11645 2789 11679
rect 2789 11645 2823 11679
rect 2823 11645 2832 11679
rect 2780 11636 2832 11645
rect 5816 11747 5868 11756
rect 5816 11713 5825 11747
rect 5825 11713 5859 11747
rect 5859 11713 5868 11747
rect 5816 11704 5868 11713
rect 6920 11747 6972 11756
rect 6920 11713 6929 11747
rect 6929 11713 6963 11747
rect 6963 11713 6972 11747
rect 6920 11704 6972 11713
rect 7656 11704 7708 11756
rect 7748 11704 7800 11756
rect 7104 11679 7156 11688
rect 7104 11645 7113 11679
rect 7113 11645 7147 11679
rect 7147 11645 7156 11679
rect 7104 11636 7156 11645
rect 10876 11747 10928 11756
rect 10876 11713 10885 11747
rect 10885 11713 10919 11747
rect 10919 11713 10928 11747
rect 10876 11704 10928 11713
rect 11428 11704 11480 11756
rect 11796 11704 11848 11756
rect 12072 11704 12124 11756
rect 12348 11747 12400 11756
rect 12348 11713 12357 11747
rect 12357 11713 12391 11747
rect 12391 11713 12400 11747
rect 12348 11704 12400 11713
rect 12440 11704 12492 11756
rect 17224 11747 17276 11756
rect 7932 11500 7984 11552
rect 11244 11500 11296 11552
rect 17224 11713 17233 11747
rect 17233 11713 17267 11747
rect 17267 11713 17276 11747
rect 17224 11704 17276 11713
rect 13728 11679 13780 11688
rect 13728 11645 13737 11679
rect 13737 11645 13771 11679
rect 13771 11645 13780 11679
rect 13728 11636 13780 11645
rect 18236 11747 18288 11756
rect 18236 11713 18245 11747
rect 18245 11713 18279 11747
rect 18279 11713 18288 11747
rect 18236 11704 18288 11713
rect 18880 11747 18932 11756
rect 18880 11713 18889 11747
rect 18889 11713 18923 11747
rect 18923 11713 18932 11747
rect 18880 11704 18932 11713
rect 22008 11704 22060 11756
rect 20904 11636 20956 11688
rect 21180 11679 21232 11688
rect 21180 11645 21189 11679
rect 21189 11645 21223 11679
rect 21223 11645 21232 11679
rect 21180 11636 21232 11645
rect 22744 11636 22796 11688
rect 30380 11772 30432 11824
rect 32772 11840 32824 11892
rect 37648 11840 37700 11892
rect 37096 11772 37148 11824
rect 37188 11772 37240 11824
rect 40960 11815 41012 11824
rect 27436 11747 27488 11756
rect 27436 11713 27445 11747
rect 27445 11713 27479 11747
rect 27479 11713 27488 11747
rect 27436 11704 27488 11713
rect 27620 11747 27672 11756
rect 27620 11713 27629 11747
rect 27629 11713 27663 11747
rect 27663 11713 27672 11747
rect 27620 11704 27672 11713
rect 29000 11747 29052 11756
rect 29000 11713 29009 11747
rect 29009 11713 29043 11747
rect 29043 11713 29052 11747
rect 29000 11704 29052 11713
rect 28172 11636 28224 11688
rect 28908 11636 28960 11688
rect 30656 11747 30708 11756
rect 30656 11713 30665 11747
rect 30665 11713 30699 11747
rect 30699 11713 30708 11747
rect 30656 11704 30708 11713
rect 30840 11747 30892 11756
rect 30840 11713 30849 11747
rect 30849 11713 30883 11747
rect 30883 11713 30892 11747
rect 30840 11704 30892 11713
rect 31024 11747 31076 11756
rect 31024 11713 31033 11747
rect 31033 11713 31067 11747
rect 31067 11713 31076 11747
rect 31024 11704 31076 11713
rect 31208 11704 31260 11756
rect 32312 11747 32364 11756
rect 32312 11713 32321 11747
rect 32321 11713 32355 11747
rect 32355 11713 32364 11747
rect 32312 11704 32364 11713
rect 32496 11747 32548 11756
rect 32496 11713 32505 11747
rect 32505 11713 32539 11747
rect 32539 11713 32548 11747
rect 32496 11704 32548 11713
rect 33600 11704 33652 11756
rect 35900 11704 35952 11756
rect 36360 11747 36412 11756
rect 36360 11713 36369 11747
rect 36369 11713 36403 11747
rect 36403 11713 36412 11747
rect 36360 11704 36412 11713
rect 37280 11704 37332 11756
rect 38200 11704 38252 11756
rect 40960 11781 40994 11815
rect 40994 11781 41012 11815
rect 40960 11772 41012 11781
rect 38660 11747 38712 11756
rect 38660 11713 38694 11747
rect 38694 11713 38712 11747
rect 38660 11704 38712 11713
rect 40684 11747 40736 11756
rect 40684 11713 40693 11747
rect 40693 11713 40727 11747
rect 40727 11713 40736 11747
rect 40684 11704 40736 11713
rect 35992 11636 36044 11688
rect 36452 11679 36504 11688
rect 36452 11645 36461 11679
rect 36461 11645 36495 11679
rect 36495 11645 36504 11679
rect 36452 11636 36504 11645
rect 25596 11568 25648 11620
rect 27620 11568 27672 11620
rect 20076 11500 20128 11552
rect 20812 11500 20864 11552
rect 20904 11500 20956 11552
rect 21456 11500 21508 11552
rect 22284 11500 22336 11552
rect 23388 11500 23440 11552
rect 27160 11500 27212 11552
rect 30472 11568 30524 11620
rect 31024 11500 31076 11552
rect 32220 11500 32272 11552
rect 36636 11500 36688 11552
rect 37464 11500 37516 11552
rect 37924 11500 37976 11552
rect 41880 11500 41932 11552
rect 6423 11398 6475 11450
rect 6487 11398 6539 11450
rect 6551 11398 6603 11450
rect 6615 11398 6667 11450
rect 6679 11398 6731 11450
rect 17370 11398 17422 11450
rect 17434 11398 17486 11450
rect 17498 11398 17550 11450
rect 17562 11398 17614 11450
rect 17626 11398 17678 11450
rect 28317 11398 28369 11450
rect 28381 11398 28433 11450
rect 28445 11398 28497 11450
rect 28509 11398 28561 11450
rect 28573 11398 28625 11450
rect 39264 11398 39316 11450
rect 39328 11398 39380 11450
rect 39392 11398 39444 11450
rect 39456 11398 39508 11450
rect 39520 11398 39572 11450
rect 3424 11339 3476 11348
rect 3424 11305 3433 11339
rect 3433 11305 3467 11339
rect 3467 11305 3476 11339
rect 3424 11296 3476 11305
rect 4436 11296 4488 11348
rect 5356 11339 5408 11348
rect 5356 11305 5365 11339
rect 5365 11305 5399 11339
rect 5399 11305 5408 11339
rect 5356 11296 5408 11305
rect 6920 11296 6972 11348
rect 9864 11296 9916 11348
rect 12072 11296 12124 11348
rect 13452 11339 13504 11348
rect 13452 11305 13461 11339
rect 13461 11305 13495 11339
rect 13495 11305 13504 11339
rect 13452 11296 13504 11305
rect 17776 11296 17828 11348
rect 20076 11339 20128 11348
rect 20076 11305 20085 11339
rect 20085 11305 20119 11339
rect 20119 11305 20128 11339
rect 20076 11296 20128 11305
rect 4620 11203 4672 11212
rect 4620 11169 4629 11203
rect 4629 11169 4663 11203
rect 4663 11169 4672 11203
rect 4620 11160 4672 11169
rect 3332 11092 3384 11144
rect 3424 11092 3476 11144
rect 5172 11135 5224 11144
rect 5172 11101 5181 11135
rect 5181 11101 5215 11135
rect 5215 11101 5224 11135
rect 5172 11092 5224 11101
rect 5540 11092 5592 11144
rect 11244 11203 11296 11212
rect 11244 11169 11253 11203
rect 11253 11169 11287 11203
rect 11287 11169 11296 11203
rect 11244 11160 11296 11169
rect 12440 11160 12492 11212
rect 13728 11228 13780 11280
rect 18236 11228 18288 11280
rect 20260 11228 20312 11280
rect 25596 11296 25648 11348
rect 22008 11228 22060 11280
rect 7932 11135 7984 11144
rect 7932 11101 7941 11135
rect 7941 11101 7975 11135
rect 7975 11101 7984 11135
rect 7932 11092 7984 11101
rect 9956 11135 10008 11144
rect 9956 11101 9965 11135
rect 9965 11101 9999 11135
rect 9999 11101 10008 11135
rect 9956 11092 10008 11101
rect 14464 11160 14516 11212
rect 13636 11135 13688 11144
rect 13636 11101 13645 11135
rect 13645 11101 13679 11135
rect 13679 11101 13688 11135
rect 13636 11092 13688 11101
rect 15384 11092 15436 11144
rect 17132 11160 17184 11212
rect 18328 11160 18380 11212
rect 19984 11160 20036 11212
rect 20628 11160 20680 11212
rect 20720 11203 20772 11212
rect 20720 11169 20729 11203
rect 20729 11169 20763 11203
rect 20763 11169 20772 11203
rect 20720 11160 20772 11169
rect 20996 11203 21048 11212
rect 20996 11169 21005 11203
rect 21005 11169 21039 11203
rect 21039 11169 21048 11203
rect 20996 11160 21048 11169
rect 24860 11160 24912 11212
rect 26792 11160 26844 11212
rect 26884 11203 26936 11212
rect 26884 11169 26893 11203
rect 26893 11169 26927 11203
rect 26927 11169 26936 11203
rect 26884 11160 26936 11169
rect 27160 11228 27212 11280
rect 27896 11228 27948 11280
rect 28540 11160 28592 11212
rect 2872 11024 2924 11076
rect 3884 11024 3936 11076
rect 13176 11024 13228 11076
rect 16304 11024 16356 11076
rect 18236 11092 18288 11144
rect 22100 11092 22152 11144
rect 23388 11135 23440 11144
rect 23388 11101 23397 11135
rect 23397 11101 23431 11135
rect 23431 11101 23440 11135
rect 23388 11092 23440 11101
rect 27620 11092 27672 11144
rect 30380 11296 30432 11348
rect 30564 11296 30616 11348
rect 31576 11296 31628 11348
rect 38660 11296 38712 11348
rect 41052 11296 41104 11348
rect 41420 11339 41472 11348
rect 41420 11305 41429 11339
rect 41429 11305 41463 11339
rect 41463 11305 41472 11339
rect 41420 11296 41472 11305
rect 28724 11228 28776 11280
rect 35808 11228 35860 11280
rect 37556 11228 37608 11280
rect 32220 11160 32272 11212
rect 20720 11024 20772 11076
rect 26424 11024 26476 11076
rect 27436 11024 27488 11076
rect 28908 11135 28960 11144
rect 28908 11101 28943 11135
rect 28943 11101 28960 11135
rect 28908 11092 28960 11101
rect 30472 11135 30524 11144
rect 30472 11101 30481 11135
rect 30481 11101 30515 11135
rect 30515 11101 30524 11135
rect 30472 11092 30524 11101
rect 30932 11135 30984 11144
rect 30932 11101 30941 11135
rect 30941 11101 30975 11135
rect 30975 11101 30984 11135
rect 30932 11092 30984 11101
rect 32312 11092 32364 11144
rect 36084 11160 36136 11212
rect 40224 11228 40276 11280
rect 33600 11092 33652 11144
rect 35072 11135 35124 11144
rect 35072 11101 35081 11135
rect 35081 11101 35115 11135
rect 35115 11101 35124 11135
rect 35072 11092 35124 11101
rect 35992 11135 36044 11144
rect 35992 11101 36001 11135
rect 36001 11101 36035 11135
rect 36035 11101 36044 11135
rect 35992 11092 36044 11101
rect 36176 11092 36228 11144
rect 37188 11135 37240 11144
rect 37188 11101 37197 11135
rect 37197 11101 37231 11135
rect 37231 11101 37240 11135
rect 37188 11092 37240 11101
rect 37280 11092 37332 11144
rect 41880 11203 41932 11212
rect 41880 11169 41889 11203
rect 41889 11169 41923 11203
rect 41923 11169 41932 11203
rect 41880 11160 41932 11169
rect 41972 11203 42024 11212
rect 41972 11169 41981 11203
rect 41981 11169 42015 11203
rect 42015 11169 42024 11203
rect 41972 11160 42024 11169
rect 39120 11092 39172 11144
rect 45008 11092 45060 11144
rect 3976 10999 4028 11008
rect 3976 10965 3985 10999
rect 3985 10965 4019 10999
rect 4019 10965 4028 10999
rect 3976 10956 4028 10965
rect 10692 10956 10744 11008
rect 11152 10999 11204 11008
rect 11152 10965 11161 10999
rect 11161 10965 11195 10999
rect 11195 10965 11204 10999
rect 11152 10956 11204 10965
rect 12256 10956 12308 11008
rect 16028 10956 16080 11008
rect 20904 10956 20956 11008
rect 20996 10956 21048 11008
rect 26700 10956 26752 11008
rect 27620 10956 27672 11008
rect 30656 11024 30708 11076
rect 34796 11024 34848 11076
rect 35808 11067 35860 11076
rect 35808 11033 35817 11067
rect 35817 11033 35851 11067
rect 35851 11033 35860 11067
rect 35808 11024 35860 11033
rect 37372 11067 37424 11076
rect 37372 11033 37381 11067
rect 37381 11033 37415 11067
rect 37415 11033 37424 11067
rect 37372 11024 37424 11033
rect 37464 11067 37516 11076
rect 37464 11033 37473 11067
rect 37473 11033 37507 11067
rect 37507 11033 37516 11067
rect 37464 11024 37516 11033
rect 39764 11024 39816 11076
rect 41788 11067 41840 11076
rect 41788 11033 41797 11067
rect 41797 11033 41831 11067
rect 41831 11033 41840 11067
rect 41788 11024 41840 11033
rect 30288 10956 30340 11008
rect 33140 10999 33192 11008
rect 33140 10965 33149 10999
rect 33149 10965 33183 10999
rect 33183 10965 33192 10999
rect 33140 10956 33192 10965
rect 33508 10956 33560 11008
rect 34520 10956 34572 11008
rect 36820 10956 36872 11008
rect 38108 10956 38160 11008
rect 11896 10854 11948 10906
rect 11960 10854 12012 10906
rect 12024 10854 12076 10906
rect 12088 10854 12140 10906
rect 12152 10854 12204 10906
rect 22843 10854 22895 10906
rect 22907 10854 22959 10906
rect 22971 10854 23023 10906
rect 23035 10854 23087 10906
rect 23099 10854 23151 10906
rect 33790 10854 33842 10906
rect 33854 10854 33906 10906
rect 33918 10854 33970 10906
rect 33982 10854 34034 10906
rect 34046 10854 34098 10906
rect 44737 10854 44789 10906
rect 44801 10854 44853 10906
rect 44865 10854 44917 10906
rect 44929 10854 44981 10906
rect 44993 10854 45045 10906
rect 7012 10752 7064 10804
rect 9956 10752 10008 10804
rect 11244 10752 11296 10804
rect 11336 10752 11388 10804
rect 12256 10752 12308 10804
rect 13820 10752 13872 10804
rect 5172 10684 5224 10736
rect 3240 10616 3292 10668
rect 3332 10659 3384 10668
rect 3332 10625 3341 10659
rect 3341 10625 3375 10659
rect 3375 10625 3384 10659
rect 3332 10616 3384 10625
rect 4988 10616 5040 10668
rect 5356 10659 5408 10668
rect 5356 10625 5365 10659
rect 5365 10625 5399 10659
rect 5399 10625 5408 10659
rect 5356 10616 5408 10625
rect 4344 10480 4396 10532
rect 17224 10752 17276 10804
rect 19248 10752 19300 10804
rect 20996 10752 21048 10804
rect 21180 10752 21232 10804
rect 25596 10795 25648 10804
rect 25596 10761 25605 10795
rect 25605 10761 25639 10795
rect 25639 10761 25648 10795
rect 25596 10752 25648 10761
rect 26700 10752 26752 10804
rect 11152 10616 11204 10668
rect 12900 10616 12952 10668
rect 13268 10616 13320 10668
rect 10876 10591 10928 10600
rect 10876 10557 10885 10591
rect 10885 10557 10919 10591
rect 10919 10557 10928 10591
rect 10876 10548 10928 10557
rect 10968 10591 11020 10600
rect 10968 10557 10977 10591
rect 10977 10557 11011 10591
rect 11011 10557 11020 10591
rect 10968 10548 11020 10557
rect 12440 10591 12492 10600
rect 12440 10557 12449 10591
rect 12449 10557 12483 10591
rect 12483 10557 12492 10591
rect 12440 10548 12492 10557
rect 16028 10659 16080 10668
rect 16028 10625 16037 10659
rect 16037 10625 16071 10659
rect 16071 10625 16080 10659
rect 16028 10616 16080 10625
rect 20260 10659 20312 10668
rect 20260 10625 20269 10659
rect 20269 10625 20303 10659
rect 20303 10625 20312 10659
rect 20260 10616 20312 10625
rect 23204 10684 23256 10736
rect 22560 10659 22612 10668
rect 22560 10625 22594 10659
rect 22594 10625 22612 10659
rect 22560 10616 22612 10625
rect 16488 10548 16540 10600
rect 940 10412 992 10464
rect 2780 10412 2832 10464
rect 5540 10412 5592 10464
rect 10140 10412 10192 10464
rect 10324 10412 10376 10464
rect 10876 10412 10928 10464
rect 15200 10412 15252 10464
rect 15660 10412 15712 10464
rect 19708 10480 19760 10532
rect 21272 10480 21324 10532
rect 18604 10412 18656 10464
rect 22192 10548 22244 10600
rect 26884 10684 26936 10736
rect 28172 10684 28224 10736
rect 30932 10795 30984 10804
rect 30932 10761 30941 10795
rect 30941 10761 30975 10795
rect 30975 10761 30984 10795
rect 30932 10752 30984 10761
rect 31484 10684 31536 10736
rect 25228 10616 25280 10668
rect 26056 10616 26108 10668
rect 29644 10659 29696 10668
rect 29644 10625 29653 10659
rect 29653 10625 29687 10659
rect 29687 10625 29696 10659
rect 33508 10684 33560 10736
rect 37280 10752 37332 10804
rect 38108 10752 38160 10804
rect 39672 10684 39724 10736
rect 29644 10616 29696 10625
rect 37556 10616 37608 10668
rect 27160 10591 27212 10600
rect 27160 10557 27169 10591
rect 27169 10557 27203 10591
rect 27203 10557 27212 10591
rect 27160 10548 27212 10557
rect 27436 10591 27488 10600
rect 27436 10557 27445 10591
rect 27445 10557 27479 10591
rect 27479 10557 27488 10591
rect 27436 10548 27488 10557
rect 29092 10548 29144 10600
rect 23664 10455 23716 10464
rect 23664 10421 23673 10455
rect 23673 10421 23707 10455
rect 23707 10421 23716 10455
rect 23664 10412 23716 10421
rect 26332 10455 26384 10464
rect 26332 10421 26341 10455
rect 26341 10421 26375 10455
rect 26375 10421 26384 10455
rect 26332 10412 26384 10421
rect 29000 10412 29052 10464
rect 32404 10412 32456 10464
rect 33140 10548 33192 10600
rect 37280 10548 37332 10600
rect 39948 10616 40000 10668
rect 40684 10659 40736 10668
rect 40684 10625 40693 10659
rect 40693 10625 40727 10659
rect 40727 10625 40736 10659
rect 40684 10616 40736 10625
rect 42800 10659 42852 10668
rect 42800 10625 42809 10659
rect 42809 10625 42843 10659
rect 42843 10625 42852 10659
rect 42800 10616 42852 10625
rect 34888 10480 34940 10532
rect 35164 10412 35216 10464
rect 39856 10412 39908 10464
rect 40592 10480 40644 10532
rect 40408 10412 40460 10464
rect 6423 10310 6475 10362
rect 6487 10310 6539 10362
rect 6551 10310 6603 10362
rect 6615 10310 6667 10362
rect 6679 10310 6731 10362
rect 17370 10310 17422 10362
rect 17434 10310 17486 10362
rect 17498 10310 17550 10362
rect 17562 10310 17614 10362
rect 17626 10310 17678 10362
rect 28317 10310 28369 10362
rect 28381 10310 28433 10362
rect 28445 10310 28497 10362
rect 28509 10310 28561 10362
rect 28573 10310 28625 10362
rect 39264 10310 39316 10362
rect 39328 10310 39380 10362
rect 39392 10310 39444 10362
rect 39456 10310 39508 10362
rect 39520 10310 39572 10362
rect 2872 10251 2924 10260
rect 2872 10217 2881 10251
rect 2881 10217 2915 10251
rect 2915 10217 2924 10251
rect 2872 10208 2924 10217
rect 3240 10208 3292 10260
rect 11244 10208 11296 10260
rect 14280 10208 14332 10260
rect 16028 10208 16080 10260
rect 16488 10251 16540 10260
rect 16488 10217 16497 10251
rect 16497 10217 16531 10251
rect 16531 10217 16540 10251
rect 16488 10208 16540 10217
rect 18880 10208 18932 10260
rect 20904 10208 20956 10260
rect 26424 10208 26476 10260
rect 26792 10251 26844 10260
rect 26792 10217 26801 10251
rect 26801 10217 26835 10251
rect 26835 10217 26844 10251
rect 26792 10208 26844 10217
rect 28172 10208 28224 10260
rect 30840 10208 30892 10260
rect 11520 10140 11572 10192
rect 4620 10115 4672 10124
rect 4620 10081 4629 10115
rect 4629 10081 4663 10115
rect 4663 10081 4672 10115
rect 4620 10072 4672 10081
rect 5816 10072 5868 10124
rect 10324 10115 10376 10124
rect 10324 10081 10333 10115
rect 10333 10081 10367 10115
rect 10367 10081 10376 10115
rect 10324 10072 10376 10081
rect 10692 10115 10744 10124
rect 10692 10081 10701 10115
rect 10701 10081 10735 10115
rect 10735 10081 10744 10115
rect 10692 10072 10744 10081
rect 14832 10140 14884 10192
rect 18604 10140 18656 10192
rect 21732 10140 21784 10192
rect 22744 10140 22796 10192
rect 3976 10004 4028 10056
rect 4344 10047 4396 10056
rect 4344 10013 4353 10047
rect 4353 10013 4387 10047
rect 4387 10013 4396 10047
rect 4344 10004 4396 10013
rect 6276 10004 6328 10056
rect 16580 10072 16632 10124
rect 17776 10115 17828 10124
rect 17776 10081 17785 10115
rect 17785 10081 17819 10115
rect 17819 10081 17828 10115
rect 17776 10072 17828 10081
rect 12440 10004 12492 10056
rect 13176 10047 13228 10056
rect 13176 10013 13185 10047
rect 13185 10013 13219 10047
rect 13219 10013 13228 10047
rect 13176 10004 13228 10013
rect 13452 10004 13504 10056
rect 14280 10047 14332 10056
rect 14280 10013 14289 10047
rect 14289 10013 14323 10047
rect 14323 10013 14332 10047
rect 14280 10004 14332 10013
rect 4436 9911 4488 9920
rect 4436 9877 4445 9911
rect 4445 9877 4479 9911
rect 4479 9877 4488 9911
rect 4436 9868 4488 9877
rect 7932 9911 7984 9920
rect 7932 9877 7941 9911
rect 7941 9877 7975 9911
rect 7975 9877 7984 9911
rect 7932 9868 7984 9877
rect 12348 9868 12400 9920
rect 14832 9868 14884 9920
rect 17224 10004 17276 10056
rect 17960 10004 18012 10056
rect 18328 10047 18380 10056
rect 18328 10013 18337 10047
rect 18337 10013 18371 10047
rect 18371 10013 18380 10047
rect 18328 10004 18380 10013
rect 18512 10047 18564 10056
rect 18512 10013 18521 10047
rect 18521 10013 18555 10047
rect 18555 10013 18564 10047
rect 18512 10004 18564 10013
rect 19708 10047 19760 10056
rect 19708 10013 19717 10047
rect 19717 10013 19751 10047
rect 19751 10013 19760 10047
rect 19708 10004 19760 10013
rect 19248 9868 19300 9920
rect 22192 10072 22244 10124
rect 30472 10140 30524 10192
rect 20812 10004 20864 10056
rect 23204 10047 23256 10056
rect 23204 10013 23213 10047
rect 23213 10013 23247 10047
rect 23247 10013 23256 10047
rect 23204 10004 23256 10013
rect 26332 10047 26384 10056
rect 26332 10013 26341 10047
rect 26341 10013 26375 10047
rect 26375 10013 26384 10047
rect 26332 10004 26384 10013
rect 27620 10072 27672 10124
rect 27896 10072 27948 10124
rect 28172 10072 28224 10124
rect 29000 10004 29052 10056
rect 30380 10004 30432 10056
rect 21272 9936 21324 9988
rect 30288 9936 30340 9988
rect 31300 10047 31352 10056
rect 31300 10013 31309 10047
rect 31309 10013 31343 10047
rect 31343 10013 31352 10047
rect 31300 10004 31352 10013
rect 33600 10251 33652 10260
rect 33600 10217 33609 10251
rect 33609 10217 33643 10251
rect 33643 10217 33652 10251
rect 33600 10208 33652 10217
rect 36360 10208 36412 10260
rect 39764 10208 39816 10260
rect 39948 10208 40000 10260
rect 40316 10208 40368 10260
rect 31852 10072 31904 10124
rect 32220 10072 32272 10124
rect 34888 10115 34940 10124
rect 34888 10081 34897 10115
rect 34897 10081 34931 10115
rect 34931 10081 34940 10115
rect 34888 10072 34940 10081
rect 35164 10115 35216 10124
rect 35164 10081 35173 10115
rect 35173 10081 35207 10115
rect 35207 10081 35216 10115
rect 35164 10072 35216 10081
rect 35900 10072 35952 10124
rect 37188 10115 37240 10124
rect 37188 10081 37197 10115
rect 37197 10081 37231 10115
rect 37231 10081 37240 10115
rect 37188 10072 37240 10081
rect 37556 10115 37608 10124
rect 37556 10081 37565 10115
rect 37565 10081 37599 10115
rect 37599 10081 37608 10115
rect 37556 10072 37608 10081
rect 40500 10140 40552 10192
rect 42800 10251 42852 10260
rect 42800 10217 42809 10251
rect 42809 10217 42843 10251
rect 42843 10217 42852 10251
rect 42800 10208 42852 10217
rect 39856 10072 39908 10124
rect 20996 9868 21048 9920
rect 21180 9868 21232 9920
rect 23480 9868 23532 9920
rect 29552 9868 29604 9920
rect 31116 9936 31168 9988
rect 31576 9979 31628 9988
rect 31576 9945 31611 9979
rect 31611 9945 31628 9979
rect 32404 10047 32456 10056
rect 32404 10013 32413 10047
rect 32413 10013 32447 10047
rect 32447 10013 32456 10047
rect 32404 10004 32456 10013
rect 33692 10004 33744 10056
rect 34520 10004 34572 10056
rect 36728 10004 36780 10056
rect 37648 10047 37700 10056
rect 37648 10013 37657 10047
rect 37657 10013 37691 10047
rect 37691 10013 37700 10047
rect 37648 10004 37700 10013
rect 38108 10047 38160 10056
rect 38108 10013 38117 10047
rect 38117 10013 38151 10047
rect 38151 10013 38160 10047
rect 38108 10004 38160 10013
rect 31576 9936 31628 9945
rect 34796 9936 34848 9988
rect 40224 10047 40276 10056
rect 40224 10013 40233 10047
rect 40233 10013 40267 10047
rect 40267 10013 40276 10047
rect 40224 10004 40276 10013
rect 40408 10047 40460 10056
rect 40408 10013 40417 10047
rect 40417 10013 40451 10047
rect 40451 10013 40460 10047
rect 40408 10004 40460 10013
rect 40500 10047 40552 10056
rect 40500 10013 40509 10047
rect 40509 10013 40543 10047
rect 40543 10013 40552 10047
rect 40500 10004 40552 10013
rect 40684 10072 40736 10124
rect 42892 10047 42944 10056
rect 42892 10013 42901 10047
rect 42901 10013 42935 10047
rect 42935 10013 42944 10047
rect 42892 10004 42944 10013
rect 32956 9868 33008 9920
rect 35992 9868 36044 9920
rect 40040 9868 40092 9920
rect 40500 9868 40552 9920
rect 40960 9868 41012 9920
rect 11896 9766 11948 9818
rect 11960 9766 12012 9818
rect 12024 9766 12076 9818
rect 12088 9766 12140 9818
rect 12152 9766 12204 9818
rect 22843 9766 22895 9818
rect 22907 9766 22959 9818
rect 22971 9766 23023 9818
rect 23035 9766 23087 9818
rect 23099 9766 23151 9818
rect 33790 9766 33842 9818
rect 33854 9766 33906 9818
rect 33918 9766 33970 9818
rect 33982 9766 34034 9818
rect 34046 9766 34098 9818
rect 44737 9766 44789 9818
rect 44801 9766 44853 9818
rect 44865 9766 44917 9818
rect 44929 9766 44981 9818
rect 44993 9766 45045 9818
rect 13452 9707 13504 9716
rect 13452 9673 13461 9707
rect 13461 9673 13495 9707
rect 13495 9673 13504 9707
rect 13452 9664 13504 9673
rect 13544 9664 13596 9716
rect 17776 9664 17828 9716
rect 2504 9596 2556 9648
rect 3148 9528 3200 9580
rect 7932 9596 7984 9648
rect 12256 9596 12308 9648
rect 13268 9596 13320 9648
rect 5632 9571 5684 9580
rect 5632 9537 5641 9571
rect 5641 9537 5675 9571
rect 5675 9537 5684 9571
rect 5632 9528 5684 9537
rect 10692 9528 10744 9580
rect 13084 9528 13136 9580
rect 13360 9528 13412 9580
rect 5816 9503 5868 9512
rect 5816 9469 5825 9503
rect 5825 9469 5859 9503
rect 5859 9469 5868 9503
rect 5816 9460 5868 9469
rect 6276 9460 6328 9512
rect 10876 9503 10928 9512
rect 10876 9469 10885 9503
rect 10885 9469 10919 9503
rect 10919 9469 10928 9503
rect 10876 9460 10928 9469
rect 10968 9503 11020 9512
rect 10968 9469 10977 9503
rect 10977 9469 11011 9503
rect 11011 9469 11020 9503
rect 10968 9460 11020 9469
rect 14096 9571 14148 9580
rect 14096 9537 14105 9571
rect 14105 9537 14139 9571
rect 14139 9537 14148 9571
rect 14096 9528 14148 9537
rect 17132 9571 17184 9580
rect 17132 9537 17166 9571
rect 17166 9537 17184 9571
rect 17132 9528 17184 9537
rect 3884 9435 3936 9444
rect 3884 9401 3893 9435
rect 3893 9401 3927 9435
rect 3927 9401 3936 9435
rect 3884 9392 3936 9401
rect 7656 9392 7708 9444
rect 2780 9324 2832 9376
rect 6184 9324 6236 9376
rect 11152 9324 11204 9376
rect 12992 9392 13044 9444
rect 13360 9392 13412 9444
rect 13820 9324 13872 9376
rect 14924 9503 14976 9512
rect 14924 9469 14933 9503
rect 14933 9469 14967 9503
rect 14967 9469 14976 9503
rect 14924 9460 14976 9469
rect 16856 9503 16908 9512
rect 16856 9469 16865 9503
rect 16865 9469 16899 9503
rect 16899 9469 16908 9503
rect 16856 9460 16908 9469
rect 14004 9392 14056 9444
rect 16304 9435 16356 9444
rect 16304 9401 16313 9435
rect 16313 9401 16347 9435
rect 16347 9401 16356 9435
rect 16304 9392 16356 9401
rect 22008 9664 22060 9716
rect 20812 9596 20864 9648
rect 23848 9596 23900 9648
rect 27436 9664 27488 9716
rect 31300 9664 31352 9716
rect 31668 9664 31720 9716
rect 35900 9664 35952 9716
rect 36360 9664 36412 9716
rect 21088 9571 21140 9580
rect 21088 9537 21097 9571
rect 21097 9537 21131 9571
rect 21131 9537 21140 9571
rect 21088 9528 21140 9537
rect 21180 9571 21232 9580
rect 21180 9537 21189 9571
rect 21189 9537 21223 9571
rect 21223 9537 21232 9571
rect 21180 9528 21232 9537
rect 22100 9528 22152 9580
rect 23296 9528 23348 9580
rect 20904 9460 20956 9512
rect 20996 9460 21048 9512
rect 21732 9460 21784 9512
rect 29644 9596 29696 9648
rect 32864 9639 32916 9648
rect 32864 9605 32873 9639
rect 32873 9605 32907 9639
rect 32907 9605 32916 9639
rect 32864 9596 32916 9605
rect 25228 9571 25280 9580
rect 25228 9537 25237 9571
rect 25237 9537 25271 9571
rect 25271 9537 25280 9571
rect 25228 9528 25280 9537
rect 26332 9528 26384 9580
rect 27344 9571 27396 9580
rect 27344 9537 27353 9571
rect 27353 9537 27387 9571
rect 27387 9537 27396 9571
rect 27344 9528 27396 9537
rect 27988 9571 28040 9580
rect 27988 9537 27997 9571
rect 27997 9537 28031 9571
rect 28031 9537 28040 9571
rect 27988 9528 28040 9537
rect 28080 9528 28132 9580
rect 29184 9528 29236 9580
rect 29552 9571 29604 9580
rect 29552 9537 29586 9571
rect 29586 9537 29604 9571
rect 29552 9528 29604 9537
rect 31116 9571 31168 9580
rect 31116 9537 31125 9571
rect 31125 9537 31159 9571
rect 31159 9537 31168 9571
rect 31116 9528 31168 9537
rect 31300 9571 31352 9580
rect 31300 9537 31309 9571
rect 31309 9537 31343 9571
rect 31343 9537 31352 9571
rect 31300 9528 31352 9537
rect 32220 9528 32272 9580
rect 32956 9528 33008 9580
rect 33416 9571 33468 9580
rect 33416 9537 33425 9571
rect 33425 9537 33459 9571
rect 33459 9537 33468 9571
rect 33416 9528 33468 9537
rect 35164 9596 35216 9648
rect 39672 9664 39724 9716
rect 39948 9664 40000 9716
rect 40500 9664 40552 9716
rect 29000 9460 29052 9512
rect 29276 9503 29328 9512
rect 29276 9469 29285 9503
rect 29285 9469 29319 9503
rect 29319 9469 29328 9503
rect 29276 9460 29328 9469
rect 36360 9460 36412 9512
rect 18236 9367 18288 9376
rect 18236 9333 18245 9367
rect 18245 9333 18279 9367
rect 18279 9333 18288 9367
rect 18236 9324 18288 9333
rect 19340 9367 19392 9376
rect 19340 9333 19349 9367
rect 19349 9333 19383 9367
rect 19383 9333 19392 9367
rect 19340 9324 19392 9333
rect 20352 9324 20404 9376
rect 20720 9367 20772 9376
rect 20720 9333 20729 9367
rect 20729 9333 20763 9367
rect 20763 9333 20772 9367
rect 20720 9324 20772 9333
rect 22100 9324 22152 9376
rect 27712 9392 27764 9444
rect 25320 9324 25372 9376
rect 27068 9324 27120 9376
rect 27804 9367 27856 9376
rect 27804 9333 27813 9367
rect 27813 9333 27847 9367
rect 27847 9333 27856 9367
rect 27804 9324 27856 9333
rect 27896 9324 27948 9376
rect 32220 9392 32272 9444
rect 32312 9392 32364 9444
rect 36728 9571 36780 9580
rect 36728 9537 36737 9571
rect 36737 9537 36771 9571
rect 36771 9537 36780 9571
rect 36728 9528 36780 9537
rect 36820 9571 36872 9580
rect 36820 9537 36829 9571
rect 36829 9537 36863 9571
rect 36863 9537 36872 9571
rect 36820 9528 36872 9537
rect 37464 9571 37516 9580
rect 37464 9537 37473 9571
rect 37473 9537 37507 9571
rect 37507 9537 37516 9571
rect 37464 9528 37516 9537
rect 37556 9460 37608 9512
rect 37648 9392 37700 9444
rect 42892 9596 42944 9648
rect 39764 9528 39816 9580
rect 39948 9528 40000 9580
rect 40408 9528 40460 9580
rect 40132 9503 40184 9512
rect 40132 9469 40141 9503
rect 40141 9469 40175 9503
rect 40175 9469 40184 9503
rect 40132 9460 40184 9469
rect 41604 9571 41656 9580
rect 41604 9537 41613 9571
rect 41613 9537 41647 9571
rect 41647 9537 41656 9571
rect 41604 9528 41656 9537
rect 40592 9503 40644 9512
rect 40592 9469 40626 9503
rect 40626 9469 40644 9503
rect 40592 9460 40644 9469
rect 41052 9460 41104 9512
rect 41972 9460 42024 9512
rect 39672 9392 39724 9444
rect 40040 9392 40092 9444
rect 30564 9324 30616 9376
rect 30748 9324 30800 9376
rect 37004 9324 37056 9376
rect 37556 9324 37608 9376
rect 41788 9392 41840 9444
rect 42616 9571 42668 9580
rect 42616 9537 42625 9571
rect 42625 9537 42659 9571
rect 42659 9537 42668 9571
rect 42616 9528 42668 9537
rect 42708 9528 42760 9580
rect 44180 9392 44232 9444
rect 41328 9324 41380 9376
rect 42616 9324 42668 9376
rect 42892 9324 42944 9376
rect 6423 9222 6475 9274
rect 6487 9222 6539 9274
rect 6551 9222 6603 9274
rect 6615 9222 6667 9274
rect 6679 9222 6731 9274
rect 17370 9222 17422 9274
rect 17434 9222 17486 9274
rect 17498 9222 17550 9274
rect 17562 9222 17614 9274
rect 17626 9222 17678 9274
rect 28317 9222 28369 9274
rect 28381 9222 28433 9274
rect 28445 9222 28497 9274
rect 28509 9222 28561 9274
rect 28573 9222 28625 9274
rect 39264 9222 39316 9274
rect 39328 9222 39380 9274
rect 39392 9222 39444 9274
rect 39456 9222 39508 9274
rect 39520 9222 39572 9274
rect 5816 9120 5868 9172
rect 7104 9120 7156 9172
rect 10876 9120 10928 9172
rect 7564 9095 7616 9104
rect 7564 9061 7573 9095
rect 7573 9061 7607 9095
rect 7607 9061 7616 9095
rect 7564 9052 7616 9061
rect 12256 9120 12308 9172
rect 12992 9120 13044 9172
rect 13084 9120 13136 9172
rect 14096 9052 14148 9104
rect 10692 8984 10744 9036
rect 4160 8916 4212 8968
rect 5632 8916 5684 8968
rect 6276 8848 6328 8900
rect 9956 8959 10008 8968
rect 9956 8925 9965 8959
rect 9965 8925 9999 8959
rect 9999 8925 10008 8959
rect 9956 8916 10008 8925
rect 10232 8848 10284 8900
rect 10600 8848 10652 8900
rect 10968 8848 11020 8900
rect 5540 8780 5592 8832
rect 8024 8823 8076 8832
rect 8024 8789 8033 8823
rect 8033 8789 8067 8823
rect 8067 8789 8076 8823
rect 8024 8780 8076 8789
rect 9772 8823 9824 8832
rect 9772 8789 9781 8823
rect 9781 8789 9815 8823
rect 9815 8789 9824 8823
rect 9772 8780 9824 8789
rect 10324 8780 10376 8832
rect 13544 8984 13596 9036
rect 17224 9120 17276 9172
rect 18512 9120 18564 9172
rect 23480 9120 23532 9172
rect 23756 9120 23808 9172
rect 19340 9052 19392 9104
rect 13452 8916 13504 8968
rect 14464 8959 14516 8968
rect 14464 8925 14473 8959
rect 14473 8925 14507 8959
rect 14507 8925 14516 8959
rect 14464 8916 14516 8925
rect 19892 8984 19944 9036
rect 22560 9052 22612 9104
rect 26332 9163 26384 9172
rect 26332 9129 26341 9163
rect 26341 9129 26375 9163
rect 26375 9129 26384 9163
rect 26332 9120 26384 9129
rect 28080 9120 28132 9172
rect 29184 9163 29236 9172
rect 29184 9129 29193 9163
rect 29193 9129 29227 9163
rect 29227 9129 29236 9163
rect 29184 9120 29236 9129
rect 35164 9163 35216 9172
rect 35164 9129 35173 9163
rect 35173 9129 35207 9163
rect 35207 9129 35216 9163
rect 35164 9120 35216 9129
rect 40224 9120 40276 9172
rect 31392 9052 31444 9104
rect 23664 8984 23716 9036
rect 14924 8916 14976 8968
rect 16856 8916 16908 8968
rect 18236 8959 18288 8968
rect 18236 8925 18245 8959
rect 18245 8925 18279 8959
rect 18279 8925 18288 8959
rect 18236 8916 18288 8925
rect 20168 8916 20220 8968
rect 20352 8959 20404 8968
rect 20352 8925 20361 8959
rect 20361 8925 20395 8959
rect 20395 8925 20404 8959
rect 20352 8916 20404 8925
rect 24492 8916 24544 8968
rect 15568 8848 15620 8900
rect 20812 8848 20864 8900
rect 18052 8823 18104 8832
rect 18052 8789 18061 8823
rect 18061 8789 18095 8823
rect 18095 8789 18104 8823
rect 18052 8780 18104 8789
rect 19524 8823 19576 8832
rect 19524 8789 19533 8823
rect 19533 8789 19567 8823
rect 19567 8789 19576 8823
rect 19524 8780 19576 8789
rect 24860 8891 24912 8900
rect 24860 8857 24869 8891
rect 24869 8857 24903 8891
rect 24903 8857 24912 8891
rect 24860 8848 24912 8857
rect 25320 8848 25372 8900
rect 23204 8780 23256 8832
rect 23480 8823 23532 8832
rect 23480 8789 23489 8823
rect 23489 8789 23523 8823
rect 23523 8789 23532 8823
rect 23480 8780 23532 8789
rect 25136 8780 25188 8832
rect 27068 8916 27120 8968
rect 27528 8916 27580 8968
rect 32220 8984 32272 9036
rect 35256 8984 35308 9036
rect 35808 9052 35860 9104
rect 39856 9052 39908 9104
rect 41604 9120 41656 9172
rect 30564 8959 30616 8968
rect 30564 8925 30573 8959
rect 30573 8925 30607 8959
rect 30607 8925 30616 8959
rect 30564 8916 30616 8925
rect 31484 8916 31536 8968
rect 34152 8916 34204 8968
rect 37280 8984 37332 9036
rect 37372 8984 37424 9036
rect 26240 8780 26292 8832
rect 27896 8780 27948 8832
rect 28080 8891 28132 8900
rect 28080 8857 28114 8891
rect 28114 8857 28132 8891
rect 28080 8848 28132 8857
rect 30104 8848 30156 8900
rect 35624 8916 35676 8968
rect 29092 8780 29144 8832
rect 35072 8848 35124 8900
rect 37004 8916 37056 8968
rect 39396 8916 39448 8968
rect 39764 8916 39816 8968
rect 40040 8959 40092 8968
rect 40040 8925 40049 8959
rect 40049 8925 40083 8959
rect 40083 8925 40092 8959
rect 40040 8916 40092 8925
rect 40316 8916 40368 8968
rect 40500 8916 40552 8968
rect 31208 8780 31260 8832
rect 35624 8780 35676 8832
rect 35716 8823 35768 8832
rect 35716 8789 35725 8823
rect 35725 8789 35759 8823
rect 35759 8789 35768 8823
rect 35716 8780 35768 8789
rect 38936 8848 38988 8900
rect 39212 8891 39264 8900
rect 39212 8857 39221 8891
rect 39221 8857 39255 8891
rect 39255 8857 39264 8891
rect 39212 8848 39264 8857
rect 38476 8780 38528 8832
rect 42800 8891 42852 8900
rect 42800 8857 42834 8891
rect 42834 8857 42852 8891
rect 42800 8848 42852 8857
rect 39672 8780 39724 8832
rect 41052 8780 41104 8832
rect 42708 8780 42760 8832
rect 11896 8678 11948 8730
rect 11960 8678 12012 8730
rect 12024 8678 12076 8730
rect 12088 8678 12140 8730
rect 12152 8678 12204 8730
rect 22843 8678 22895 8730
rect 22907 8678 22959 8730
rect 22971 8678 23023 8730
rect 23035 8678 23087 8730
rect 23099 8678 23151 8730
rect 33790 8678 33842 8730
rect 33854 8678 33906 8730
rect 33918 8678 33970 8730
rect 33982 8678 34034 8730
rect 34046 8678 34098 8730
rect 44737 8678 44789 8730
rect 44801 8678 44853 8730
rect 44865 8678 44917 8730
rect 44929 8678 44981 8730
rect 44993 8678 45045 8730
rect 2780 8576 2832 8628
rect 3792 8576 3844 8628
rect 3976 8483 4028 8492
rect 3976 8449 3985 8483
rect 3985 8449 4019 8483
rect 4019 8449 4028 8483
rect 3976 8440 4028 8449
rect 4436 8508 4488 8560
rect 7656 8576 7708 8628
rect 8024 8576 8076 8628
rect 10324 8619 10376 8628
rect 10324 8585 10333 8619
rect 10333 8585 10367 8619
rect 10367 8585 10376 8619
rect 10324 8576 10376 8585
rect 10968 8619 11020 8628
rect 10968 8585 10977 8619
rect 10977 8585 11011 8619
rect 11011 8585 11020 8619
rect 10968 8576 11020 8585
rect 11612 8576 11664 8628
rect 7012 8508 7064 8560
rect 10232 8508 10284 8560
rect 11520 8508 11572 8560
rect 11888 8508 11940 8560
rect 12900 8576 12952 8628
rect 6276 8372 6328 8424
rect 8208 8440 8260 8492
rect 7932 8347 7984 8356
rect 7932 8313 7941 8347
rect 7941 8313 7975 8347
rect 7975 8313 7984 8347
rect 7932 8304 7984 8313
rect 10508 8483 10560 8492
rect 10508 8449 10517 8483
rect 10517 8449 10551 8483
rect 10551 8449 10560 8483
rect 10508 8440 10560 8449
rect 11152 8483 11204 8492
rect 11152 8449 11161 8483
rect 11161 8449 11195 8483
rect 11195 8449 11204 8483
rect 11152 8440 11204 8449
rect 10600 8372 10652 8424
rect 15660 8508 15712 8560
rect 16856 8508 16908 8560
rect 20168 8576 20220 8628
rect 21180 8576 21232 8628
rect 25136 8576 25188 8628
rect 25228 8576 25280 8628
rect 31300 8619 31352 8628
rect 31300 8585 31309 8619
rect 31309 8585 31343 8619
rect 31343 8585 31352 8619
rect 31300 8576 31352 8585
rect 16212 8440 16264 8492
rect 18052 8440 18104 8492
rect 19708 8440 19760 8492
rect 20904 8440 20956 8492
rect 21272 8440 21324 8492
rect 15384 8372 15436 8424
rect 15660 8415 15712 8424
rect 15660 8381 15669 8415
rect 15669 8381 15703 8415
rect 15703 8381 15712 8415
rect 15660 8372 15712 8381
rect 19984 8372 20036 8424
rect 20076 8415 20128 8424
rect 20076 8381 20085 8415
rect 20085 8381 20119 8415
rect 20119 8381 20128 8415
rect 20076 8372 20128 8381
rect 22468 8483 22520 8492
rect 22468 8449 22502 8483
rect 22502 8449 22520 8483
rect 22468 8440 22520 8449
rect 22192 8415 22244 8424
rect 22192 8381 22201 8415
rect 22201 8381 22235 8415
rect 22235 8381 22244 8415
rect 22192 8372 22244 8381
rect 5356 8279 5408 8288
rect 5356 8245 5365 8279
rect 5365 8245 5399 8279
rect 5399 8245 5408 8279
rect 5356 8236 5408 8245
rect 7748 8236 7800 8288
rect 11520 8236 11572 8288
rect 16856 8304 16908 8356
rect 21916 8304 21968 8356
rect 26056 8508 26108 8560
rect 27436 8508 27488 8560
rect 28172 8508 28224 8560
rect 31852 8508 31904 8560
rect 35624 8619 35676 8628
rect 35624 8585 35633 8619
rect 35633 8585 35667 8619
rect 35667 8585 35676 8619
rect 35624 8576 35676 8585
rect 37464 8576 37516 8628
rect 39396 8619 39448 8628
rect 39396 8585 39405 8619
rect 39405 8585 39439 8619
rect 39439 8585 39448 8619
rect 39396 8576 39448 8585
rect 35716 8508 35768 8560
rect 36084 8508 36136 8560
rect 37372 8508 37424 8560
rect 38752 8508 38804 8560
rect 40684 8576 40736 8628
rect 41696 8576 41748 8628
rect 25964 8440 26016 8492
rect 29644 8440 29696 8492
rect 30472 8440 30524 8492
rect 23848 8304 23900 8356
rect 27160 8304 27212 8356
rect 27528 8304 27580 8356
rect 29276 8304 29328 8356
rect 31576 8440 31628 8492
rect 31484 8372 31536 8424
rect 31668 8372 31720 8424
rect 34520 8415 34572 8424
rect 34520 8381 34529 8415
rect 34529 8381 34563 8415
rect 34563 8381 34572 8415
rect 34520 8372 34572 8381
rect 35440 8483 35492 8492
rect 35440 8449 35449 8483
rect 35449 8449 35483 8483
rect 35483 8449 35492 8483
rect 35440 8440 35492 8449
rect 35808 8483 35860 8492
rect 35808 8449 35817 8483
rect 35817 8449 35851 8483
rect 35851 8449 35860 8483
rect 35808 8440 35860 8449
rect 36360 8440 36412 8492
rect 35992 8372 36044 8424
rect 36544 8372 36596 8424
rect 31760 8304 31812 8356
rect 34152 8304 34204 8356
rect 36268 8304 36320 8356
rect 38016 8304 38068 8356
rect 38568 8483 38620 8492
rect 38568 8449 38577 8483
rect 38577 8449 38611 8483
rect 38611 8449 38620 8483
rect 38568 8440 38620 8449
rect 39764 8483 39816 8492
rect 39764 8449 39773 8483
rect 39773 8449 39807 8483
rect 39807 8449 39816 8483
rect 39764 8440 39816 8449
rect 40132 8508 40184 8560
rect 42708 8576 42760 8628
rect 42892 8619 42944 8628
rect 42892 8585 42901 8619
rect 42901 8585 42935 8619
rect 42935 8585 42944 8619
rect 42892 8576 42944 8585
rect 44180 8619 44232 8628
rect 44180 8585 44189 8619
rect 44189 8585 44223 8619
rect 44223 8585 44232 8619
rect 44180 8576 44232 8585
rect 39948 8440 40000 8492
rect 40960 8483 41012 8492
rect 40960 8449 40969 8483
rect 40969 8449 41003 8483
rect 41003 8449 41012 8483
rect 40960 8440 41012 8449
rect 41328 8440 41380 8492
rect 41696 8440 41748 8492
rect 44364 8483 44416 8492
rect 44364 8449 44373 8483
rect 44373 8449 44407 8483
rect 44407 8449 44416 8483
rect 44364 8440 44416 8449
rect 41052 8372 41104 8424
rect 18604 8279 18656 8288
rect 18604 8245 18613 8279
rect 18613 8245 18647 8279
rect 18647 8245 18656 8279
rect 18604 8236 18656 8245
rect 29184 8236 29236 8288
rect 36176 8236 36228 8288
rect 36452 8279 36504 8288
rect 36452 8245 36461 8279
rect 36461 8245 36495 8279
rect 36495 8245 36504 8279
rect 36452 8236 36504 8245
rect 38660 8279 38712 8288
rect 38660 8245 38669 8279
rect 38669 8245 38703 8279
rect 38703 8245 38712 8279
rect 38660 8236 38712 8245
rect 40408 8236 40460 8288
rect 41052 8236 41104 8288
rect 43168 8279 43220 8288
rect 43168 8245 43177 8279
rect 43177 8245 43211 8279
rect 43211 8245 43220 8279
rect 43168 8236 43220 8245
rect 6423 8134 6475 8186
rect 6487 8134 6539 8186
rect 6551 8134 6603 8186
rect 6615 8134 6667 8186
rect 6679 8134 6731 8186
rect 17370 8134 17422 8186
rect 17434 8134 17486 8186
rect 17498 8134 17550 8186
rect 17562 8134 17614 8186
rect 17626 8134 17678 8186
rect 28317 8134 28369 8186
rect 28381 8134 28433 8186
rect 28445 8134 28497 8186
rect 28509 8134 28561 8186
rect 28573 8134 28625 8186
rect 39264 8134 39316 8186
rect 39328 8134 39380 8186
rect 39392 8134 39444 8186
rect 39456 8134 39508 8186
rect 39520 8134 39572 8186
rect 6276 8032 6328 8084
rect 3148 7939 3200 7948
rect 3148 7905 3157 7939
rect 3157 7905 3191 7939
rect 3191 7905 3200 7939
rect 3148 7896 3200 7905
rect 940 7828 992 7880
rect 5540 7828 5592 7880
rect 5816 7828 5868 7880
rect 8208 7964 8260 8016
rect 7932 7896 7984 7948
rect 5448 7760 5500 7812
rect 9128 7760 9180 7812
rect 2964 7692 3016 7744
rect 5264 7692 5316 7744
rect 7288 7692 7340 7744
rect 10508 8032 10560 8084
rect 10876 8032 10928 8084
rect 16212 8075 16264 8084
rect 16212 8041 16221 8075
rect 16221 8041 16255 8075
rect 16255 8041 16264 8075
rect 16212 8032 16264 8041
rect 18236 8032 18288 8084
rect 13544 7896 13596 7948
rect 20076 8032 20128 8084
rect 22468 8032 22520 8084
rect 27988 8032 28040 8084
rect 31576 7964 31628 8016
rect 32956 8032 33008 8084
rect 36452 8032 36504 8084
rect 36544 8075 36596 8084
rect 36544 8041 36553 8075
rect 36553 8041 36587 8075
rect 36587 8041 36596 8075
rect 36544 8032 36596 8041
rect 37004 8075 37056 8084
rect 37004 8041 37013 8075
rect 37013 8041 37047 8075
rect 37047 8041 37056 8075
rect 37004 8032 37056 8041
rect 37372 8075 37424 8084
rect 37372 8041 37381 8075
rect 37381 8041 37415 8075
rect 37415 8041 37424 8075
rect 37372 8032 37424 8041
rect 39396 8032 39448 8084
rect 42800 8032 42852 8084
rect 36176 7964 36228 8016
rect 9864 7828 9916 7880
rect 10600 7828 10652 7880
rect 12900 7828 12952 7880
rect 14924 7828 14976 7880
rect 9772 7760 9824 7812
rect 15476 7828 15528 7880
rect 15660 7828 15712 7880
rect 19892 7939 19944 7948
rect 19892 7905 19901 7939
rect 19901 7905 19935 7939
rect 19935 7905 19944 7939
rect 19892 7896 19944 7905
rect 16856 7871 16908 7880
rect 16856 7837 16865 7871
rect 16865 7837 16899 7871
rect 16899 7837 16908 7871
rect 16856 7828 16908 7837
rect 18604 7828 18656 7880
rect 19524 7828 19576 7880
rect 21916 7871 21968 7880
rect 21916 7837 21925 7871
rect 21925 7837 21959 7871
rect 21959 7837 21968 7871
rect 21916 7828 21968 7837
rect 23388 7828 23440 7880
rect 23572 7828 23624 7880
rect 26148 7896 26200 7948
rect 27160 7896 27212 7948
rect 27896 7896 27948 7948
rect 28908 7896 28960 7948
rect 12256 7692 12308 7744
rect 12900 7735 12952 7744
rect 12900 7701 12909 7735
rect 12909 7701 12943 7735
rect 12943 7701 12952 7735
rect 12900 7692 12952 7701
rect 17960 7760 18012 7812
rect 27436 7828 27488 7880
rect 29644 7828 29696 7880
rect 29736 7828 29788 7880
rect 32588 7828 32640 7880
rect 34336 7939 34388 7948
rect 34336 7905 34345 7939
rect 34345 7905 34379 7939
rect 34379 7905 34388 7939
rect 34336 7896 34388 7905
rect 21272 7735 21324 7744
rect 21272 7701 21281 7735
rect 21281 7701 21315 7735
rect 21315 7701 21324 7735
rect 21272 7692 21324 7701
rect 21732 7735 21784 7744
rect 21732 7701 21741 7735
rect 21741 7701 21775 7735
rect 21775 7701 21784 7735
rect 21732 7692 21784 7701
rect 23388 7692 23440 7744
rect 27804 7760 27856 7812
rect 30564 7803 30616 7812
rect 30564 7769 30598 7803
rect 30598 7769 30616 7803
rect 30564 7760 30616 7769
rect 31944 7760 31996 7812
rect 35072 7828 35124 7880
rect 35164 7871 35216 7880
rect 35164 7837 35173 7871
rect 35173 7837 35207 7871
rect 35207 7837 35216 7871
rect 35164 7828 35216 7837
rect 38660 7896 38712 7948
rect 37096 7871 37148 7880
rect 37096 7837 37105 7871
rect 37105 7837 37139 7871
rect 37139 7837 37148 7871
rect 37096 7828 37148 7837
rect 37188 7828 37240 7880
rect 38016 7871 38068 7880
rect 38016 7837 38025 7871
rect 38025 7837 38059 7871
rect 38059 7837 38068 7871
rect 38016 7828 38068 7837
rect 38752 7828 38804 7880
rect 39304 7871 39356 7880
rect 39304 7837 39313 7871
rect 39313 7837 39347 7871
rect 39347 7837 39356 7871
rect 39304 7828 39356 7837
rect 40500 7939 40552 7948
rect 40500 7905 40509 7939
rect 40509 7905 40543 7939
rect 40543 7905 40552 7939
rect 40500 7896 40552 7905
rect 41052 7828 41104 7880
rect 43168 7828 43220 7880
rect 44364 7871 44416 7880
rect 44364 7837 44373 7871
rect 44373 7837 44407 7871
rect 44407 7837 44416 7871
rect 44364 7828 44416 7837
rect 34428 7692 34480 7744
rect 36268 7692 36320 7744
rect 37188 7692 37240 7744
rect 39580 7760 39632 7812
rect 41420 7760 41472 7812
rect 41604 7692 41656 7744
rect 43444 7692 43496 7744
rect 11896 7590 11948 7642
rect 11960 7590 12012 7642
rect 12024 7590 12076 7642
rect 12088 7590 12140 7642
rect 12152 7590 12204 7642
rect 22843 7590 22895 7642
rect 22907 7590 22959 7642
rect 22971 7590 23023 7642
rect 23035 7590 23087 7642
rect 23099 7590 23151 7642
rect 33790 7590 33842 7642
rect 33854 7590 33906 7642
rect 33918 7590 33970 7642
rect 33982 7590 34034 7642
rect 34046 7590 34098 7642
rect 44737 7590 44789 7642
rect 44801 7590 44853 7642
rect 44865 7590 44917 7642
rect 44929 7590 44981 7642
rect 44993 7590 45045 7642
rect 3976 7488 4028 7540
rect 5356 7488 5408 7540
rect 9128 7531 9180 7540
rect 9128 7497 9137 7531
rect 9137 7497 9171 7531
rect 9171 7497 9180 7531
rect 9128 7488 9180 7497
rect 11796 7488 11848 7540
rect 14464 7488 14516 7540
rect 31116 7488 31168 7540
rect 31392 7531 31444 7540
rect 31392 7497 31401 7531
rect 31401 7497 31435 7531
rect 31435 7497 31444 7531
rect 31392 7488 31444 7497
rect 5540 7420 5592 7472
rect 6920 7420 6972 7472
rect 5172 7395 5224 7404
rect 5172 7361 5181 7395
rect 5181 7361 5215 7395
rect 5215 7361 5224 7395
rect 5172 7352 5224 7361
rect 7288 7395 7340 7404
rect 7288 7361 7297 7395
rect 7297 7361 7331 7395
rect 7331 7361 7340 7395
rect 7288 7352 7340 7361
rect 7748 7395 7800 7404
rect 7748 7361 7757 7395
rect 7757 7361 7791 7395
rect 7791 7361 7800 7395
rect 7748 7352 7800 7361
rect 5080 7284 5132 7336
rect 5448 7327 5500 7336
rect 5448 7293 5457 7327
rect 5457 7293 5491 7327
rect 5491 7293 5500 7327
rect 5448 7284 5500 7293
rect 9864 7395 9916 7404
rect 9864 7361 9873 7395
rect 9873 7361 9907 7395
rect 9907 7361 9916 7395
rect 9864 7352 9916 7361
rect 12256 7352 12308 7404
rect 12624 7352 12676 7404
rect 14924 7420 14976 7472
rect 21732 7420 21784 7472
rect 23388 7463 23440 7472
rect 23388 7429 23422 7463
rect 23422 7429 23440 7463
rect 23388 7420 23440 7429
rect 27896 7420 27948 7472
rect 28908 7420 28960 7472
rect 13360 7352 13412 7404
rect 15476 7395 15528 7404
rect 15476 7361 15485 7395
rect 15485 7361 15519 7395
rect 15519 7361 15528 7395
rect 15476 7352 15528 7361
rect 16212 7352 16264 7404
rect 19892 7395 19944 7404
rect 19892 7361 19901 7395
rect 19901 7361 19935 7395
rect 19935 7361 19944 7395
rect 19892 7352 19944 7361
rect 25964 7395 26016 7404
rect 25964 7361 25973 7395
rect 25973 7361 26007 7395
rect 26007 7361 26016 7395
rect 25964 7352 26016 7361
rect 29184 7395 29236 7404
rect 29184 7361 29193 7395
rect 29193 7361 29227 7395
rect 29227 7361 29236 7395
rect 29184 7352 29236 7361
rect 29644 7395 29696 7404
rect 29644 7361 29653 7395
rect 29653 7361 29687 7395
rect 29687 7361 29696 7395
rect 29644 7352 29696 7361
rect 30656 7420 30708 7472
rect 32956 7488 33008 7540
rect 34336 7488 34388 7540
rect 37096 7488 37148 7540
rect 31852 7420 31904 7472
rect 31944 7420 31996 7472
rect 31392 7352 31444 7404
rect 31760 7352 31812 7404
rect 32220 7352 32272 7404
rect 32588 7395 32640 7404
rect 32588 7361 32597 7395
rect 32597 7361 32631 7395
rect 32631 7361 32640 7395
rect 32588 7352 32640 7361
rect 32680 7395 32732 7404
rect 32680 7361 32689 7395
rect 32689 7361 32723 7395
rect 32723 7361 32732 7395
rect 32680 7352 32732 7361
rect 32772 7395 32824 7404
rect 32772 7361 32781 7395
rect 32781 7361 32815 7395
rect 32815 7361 32824 7395
rect 32772 7352 32824 7361
rect 32956 7395 33008 7404
rect 32956 7361 32965 7395
rect 32965 7361 32999 7395
rect 32999 7361 33008 7395
rect 32956 7352 33008 7361
rect 33048 7352 33100 7404
rect 33784 7420 33836 7472
rect 33692 7352 33744 7404
rect 34336 7352 34388 7404
rect 35348 7352 35400 7404
rect 35992 7395 36044 7404
rect 35992 7361 36001 7395
rect 36001 7361 36035 7395
rect 36035 7361 36044 7395
rect 35992 7352 36044 7361
rect 15568 7327 15620 7336
rect 4252 7148 4304 7200
rect 4988 7148 5040 7200
rect 5448 7148 5500 7200
rect 10968 7148 11020 7200
rect 11060 7191 11112 7200
rect 11060 7157 11069 7191
rect 11069 7157 11103 7191
rect 11103 7157 11112 7191
rect 11060 7148 11112 7157
rect 12900 7148 12952 7200
rect 15568 7293 15577 7327
rect 15577 7293 15611 7327
rect 15611 7293 15620 7327
rect 15568 7284 15620 7293
rect 15660 7327 15712 7336
rect 15660 7293 15669 7327
rect 15669 7293 15703 7327
rect 15703 7293 15712 7327
rect 15660 7284 15712 7293
rect 22192 7284 22244 7336
rect 20904 7216 20956 7268
rect 21824 7216 21876 7268
rect 15016 7148 15068 7200
rect 15108 7191 15160 7200
rect 15108 7157 15117 7191
rect 15117 7157 15151 7191
rect 15151 7157 15160 7191
rect 15108 7148 15160 7157
rect 17960 7148 18012 7200
rect 26240 7327 26292 7336
rect 26240 7293 26249 7327
rect 26249 7293 26283 7327
rect 26283 7293 26292 7327
rect 26240 7284 26292 7293
rect 27160 7327 27212 7336
rect 27160 7293 27169 7327
rect 27169 7293 27203 7327
rect 27203 7293 27212 7327
rect 27160 7284 27212 7293
rect 28724 7284 28776 7336
rect 31576 7284 31628 7336
rect 32404 7284 32456 7336
rect 35256 7284 35308 7336
rect 35624 7284 35676 7336
rect 36268 7327 36320 7336
rect 36268 7293 36277 7327
rect 36277 7293 36311 7327
rect 36311 7293 36320 7327
rect 36268 7284 36320 7293
rect 31852 7216 31904 7268
rect 32588 7216 32640 7268
rect 34244 7216 34296 7268
rect 35072 7216 35124 7268
rect 36728 7284 36780 7336
rect 37188 7284 37240 7336
rect 38568 7531 38620 7540
rect 38568 7497 38577 7531
rect 38577 7497 38611 7531
rect 38611 7497 38620 7531
rect 38568 7488 38620 7497
rect 39304 7488 39356 7540
rect 39580 7531 39632 7540
rect 39580 7497 39589 7531
rect 39589 7497 39623 7531
rect 39623 7497 39632 7531
rect 39580 7488 39632 7497
rect 41420 7531 41472 7540
rect 41420 7497 41429 7531
rect 41429 7497 41463 7531
rect 41463 7497 41472 7531
rect 41420 7488 41472 7497
rect 41604 7395 41656 7404
rect 41604 7361 41613 7395
rect 41613 7361 41647 7395
rect 41647 7361 41656 7395
rect 41604 7352 41656 7361
rect 39396 7327 39448 7336
rect 39396 7293 39405 7327
rect 39405 7293 39439 7327
rect 39439 7293 39448 7327
rect 39396 7284 39448 7293
rect 39764 7327 39816 7336
rect 39764 7293 39773 7327
rect 39773 7293 39807 7327
rect 39807 7293 39816 7327
rect 39764 7284 39816 7293
rect 23388 7148 23440 7200
rect 24400 7148 24452 7200
rect 27620 7148 27672 7200
rect 30656 7148 30708 7200
rect 31484 7148 31536 7200
rect 32036 7148 32088 7200
rect 32312 7191 32364 7200
rect 32312 7157 32321 7191
rect 32321 7157 32355 7191
rect 32355 7157 32364 7191
rect 32312 7148 32364 7157
rect 32404 7148 32456 7200
rect 33784 7191 33836 7200
rect 33784 7157 33793 7191
rect 33793 7157 33827 7191
rect 33827 7157 33836 7191
rect 33784 7148 33836 7157
rect 34796 7148 34848 7200
rect 36636 7191 36688 7200
rect 36636 7157 36645 7191
rect 36645 7157 36679 7191
rect 36679 7157 36688 7191
rect 36636 7148 36688 7157
rect 40224 7216 40276 7268
rect 40316 7216 40368 7268
rect 40776 7284 40828 7336
rect 40868 7327 40920 7336
rect 40868 7293 40877 7327
rect 40877 7293 40911 7327
rect 40911 7293 40920 7327
rect 40868 7284 40920 7293
rect 41420 7284 41472 7336
rect 40132 7148 40184 7200
rect 6423 7046 6475 7098
rect 6487 7046 6539 7098
rect 6551 7046 6603 7098
rect 6615 7046 6667 7098
rect 6679 7046 6731 7098
rect 17370 7046 17422 7098
rect 17434 7046 17486 7098
rect 17498 7046 17550 7098
rect 17562 7046 17614 7098
rect 17626 7046 17678 7098
rect 28317 7046 28369 7098
rect 28381 7046 28433 7098
rect 28445 7046 28497 7098
rect 28509 7046 28561 7098
rect 28573 7046 28625 7098
rect 39264 7046 39316 7098
rect 39328 7046 39380 7098
rect 39392 7046 39444 7098
rect 39456 7046 39508 7098
rect 39520 7046 39572 7098
rect 3148 6944 3200 6996
rect 10140 6944 10192 6996
rect 10600 6944 10652 6996
rect 11796 6944 11848 6996
rect 13360 6944 13412 6996
rect 15660 6944 15712 6996
rect 6920 6808 6972 6860
rect 9404 6808 9456 6860
rect 10600 6808 10652 6860
rect 3884 6740 3936 6792
rect 5356 6740 5408 6792
rect 6184 6740 6236 6792
rect 7564 6740 7616 6792
rect 11060 6740 11112 6792
rect 13452 6851 13504 6860
rect 13452 6817 13461 6851
rect 13461 6817 13495 6851
rect 13495 6817 13504 6851
rect 13452 6808 13504 6817
rect 14924 6808 14976 6860
rect 20996 6944 21048 6996
rect 21456 6944 21508 6996
rect 32772 6944 32824 6996
rect 37004 6944 37056 6996
rect 40224 6944 40276 6996
rect 40776 6944 40828 6996
rect 18604 6851 18656 6860
rect 18604 6817 18613 6851
rect 18613 6817 18647 6851
rect 18647 6817 18656 6851
rect 18604 6808 18656 6817
rect 20444 6876 20496 6928
rect 20904 6876 20956 6928
rect 21272 6876 21324 6928
rect 21640 6876 21692 6928
rect 4436 6672 4488 6724
rect 10692 6672 10744 6724
rect 6828 6604 6880 6656
rect 14188 6672 14240 6724
rect 15108 6740 15160 6792
rect 18512 6783 18564 6792
rect 18512 6749 18521 6783
rect 18521 6749 18555 6783
rect 18555 6749 18564 6783
rect 18512 6740 18564 6749
rect 15016 6672 15068 6724
rect 15568 6715 15620 6724
rect 15568 6681 15602 6715
rect 15602 6681 15620 6715
rect 15568 6672 15620 6681
rect 10876 6647 10928 6656
rect 10876 6613 10885 6647
rect 10885 6613 10919 6647
rect 10919 6613 10928 6647
rect 10876 6604 10928 6613
rect 11612 6604 11664 6656
rect 14556 6604 14608 6656
rect 17776 6672 17828 6724
rect 18144 6672 18196 6724
rect 17132 6647 17184 6656
rect 17132 6613 17141 6647
rect 17141 6613 17175 6647
rect 17175 6613 17184 6647
rect 17132 6604 17184 6613
rect 17224 6604 17276 6656
rect 17868 6604 17920 6656
rect 20444 6783 20496 6792
rect 20444 6749 20456 6783
rect 20456 6749 20490 6783
rect 20490 6749 20496 6783
rect 20444 6740 20496 6749
rect 21456 6783 21508 6792
rect 21456 6749 21466 6783
rect 21466 6749 21500 6783
rect 21500 6749 21508 6783
rect 21456 6740 21508 6749
rect 21640 6783 21692 6792
rect 21640 6749 21649 6783
rect 21649 6749 21683 6783
rect 21683 6749 21692 6783
rect 21640 6740 21692 6749
rect 21824 6783 21876 6792
rect 21824 6749 21838 6783
rect 21838 6749 21872 6783
rect 21872 6749 21876 6783
rect 21824 6740 21876 6749
rect 21732 6715 21784 6724
rect 21732 6681 21741 6715
rect 21741 6681 21775 6715
rect 21775 6681 21784 6715
rect 21732 6672 21784 6681
rect 23756 6851 23808 6860
rect 23756 6817 23765 6851
rect 23765 6817 23799 6851
rect 23799 6817 23808 6851
rect 23756 6808 23808 6817
rect 23848 6851 23900 6860
rect 23848 6817 23857 6851
rect 23857 6817 23891 6851
rect 23891 6817 23900 6851
rect 23848 6808 23900 6817
rect 24400 6740 24452 6792
rect 25044 6740 25096 6792
rect 26056 6740 26108 6792
rect 27620 6808 27672 6860
rect 32404 6876 32456 6928
rect 32588 6876 32640 6928
rect 32220 6851 32272 6860
rect 32220 6817 32229 6851
rect 32229 6817 32263 6851
rect 32263 6817 32272 6851
rect 32220 6808 32272 6817
rect 33048 6808 33100 6860
rect 27252 6783 27304 6792
rect 27252 6749 27261 6783
rect 27261 6749 27295 6783
rect 27295 6749 27304 6783
rect 27252 6740 27304 6749
rect 29736 6783 29788 6792
rect 29736 6749 29745 6783
rect 29745 6749 29779 6783
rect 29779 6749 29788 6783
rect 29736 6740 29788 6749
rect 28724 6672 28776 6724
rect 31024 6672 31076 6724
rect 32588 6740 32640 6792
rect 33784 6740 33836 6792
rect 39764 6876 39816 6928
rect 40868 6876 40920 6928
rect 35164 6808 35216 6860
rect 40408 6808 40460 6860
rect 20720 6604 20772 6656
rect 22008 6647 22060 6656
rect 22008 6613 22017 6647
rect 22017 6613 22051 6647
rect 22051 6613 22060 6647
rect 22008 6604 22060 6613
rect 23572 6604 23624 6656
rect 25872 6604 25924 6656
rect 27896 6604 27948 6656
rect 30380 6604 30432 6656
rect 31944 6672 31996 6724
rect 34888 6740 34940 6792
rect 32036 6647 32088 6656
rect 32036 6613 32045 6647
rect 32045 6613 32079 6647
rect 32079 6613 32088 6647
rect 32036 6604 32088 6613
rect 32680 6604 32732 6656
rect 35532 6672 35584 6724
rect 35808 6740 35860 6792
rect 35992 6672 36044 6724
rect 36360 6715 36412 6724
rect 36360 6681 36369 6715
rect 36369 6681 36403 6715
rect 36403 6681 36412 6715
rect 36360 6672 36412 6681
rect 34152 6604 34204 6656
rect 35348 6604 35400 6656
rect 36268 6604 36320 6656
rect 36544 6783 36596 6792
rect 36544 6749 36553 6783
rect 36553 6749 36587 6783
rect 36587 6749 36596 6783
rect 36544 6740 36596 6749
rect 36636 6740 36688 6792
rect 36912 6783 36964 6792
rect 36912 6749 36921 6783
rect 36921 6749 36955 6783
rect 36955 6749 36964 6783
rect 36912 6740 36964 6749
rect 40132 6740 40184 6792
rect 40224 6783 40276 6792
rect 40224 6749 40233 6783
rect 40233 6749 40267 6783
rect 40267 6749 40276 6783
rect 40224 6740 40276 6749
rect 40500 6783 40552 6792
rect 40500 6749 40509 6783
rect 40509 6749 40543 6783
rect 40543 6749 40552 6783
rect 40500 6740 40552 6749
rect 40684 6783 40736 6792
rect 40684 6749 40693 6783
rect 40693 6749 40727 6783
rect 40727 6749 40736 6783
rect 40684 6740 40736 6749
rect 40776 6740 40828 6792
rect 43444 6851 43496 6860
rect 43444 6817 43453 6851
rect 43453 6817 43487 6851
rect 43487 6817 43496 6851
rect 43444 6808 43496 6817
rect 37372 6604 37424 6656
rect 37648 6604 37700 6656
rect 41420 6604 41472 6656
rect 43720 6647 43772 6656
rect 43720 6613 43729 6647
rect 43729 6613 43763 6647
rect 43763 6613 43772 6647
rect 43720 6604 43772 6613
rect 11896 6502 11948 6554
rect 11960 6502 12012 6554
rect 12024 6502 12076 6554
rect 12088 6502 12140 6554
rect 12152 6502 12204 6554
rect 22843 6502 22895 6554
rect 22907 6502 22959 6554
rect 22971 6502 23023 6554
rect 23035 6502 23087 6554
rect 23099 6502 23151 6554
rect 33790 6502 33842 6554
rect 33854 6502 33906 6554
rect 33918 6502 33970 6554
rect 33982 6502 34034 6554
rect 34046 6502 34098 6554
rect 44737 6502 44789 6554
rect 44801 6502 44853 6554
rect 44865 6502 44917 6554
rect 44929 6502 44981 6554
rect 44993 6502 45045 6554
rect 4344 6400 4396 6452
rect 5172 6400 5224 6452
rect 6000 6400 6052 6452
rect 9956 6400 10008 6452
rect 10692 6400 10744 6452
rect 15568 6443 15620 6452
rect 15568 6409 15577 6443
rect 15577 6409 15611 6443
rect 15611 6409 15620 6443
rect 15568 6400 15620 6409
rect 17960 6443 18012 6452
rect 17960 6409 17969 6443
rect 17969 6409 18003 6443
rect 18003 6409 18012 6443
rect 17960 6400 18012 6409
rect 4252 6375 4304 6384
rect 4252 6341 4286 6375
rect 4286 6341 4304 6375
rect 4252 6332 4304 6341
rect 10876 6332 10928 6384
rect 12532 6332 12584 6384
rect 13268 6332 13320 6384
rect 14924 6332 14976 6384
rect 15016 6332 15068 6384
rect 19248 6400 19300 6452
rect 21732 6400 21784 6452
rect 27252 6443 27304 6452
rect 27252 6409 27261 6443
rect 27261 6409 27295 6443
rect 27295 6409 27304 6443
rect 27252 6400 27304 6409
rect 30564 6400 30616 6452
rect 30656 6400 30708 6452
rect 31024 6400 31076 6452
rect 31392 6400 31444 6452
rect 33876 6400 33928 6452
rect 34428 6400 34480 6452
rect 18604 6332 18656 6384
rect 4528 6264 4580 6316
rect 8484 6307 8536 6316
rect 8484 6273 8493 6307
rect 8493 6273 8527 6307
rect 8527 6273 8536 6307
rect 8484 6264 8536 6273
rect 9036 6264 9088 6316
rect 10968 6307 11020 6316
rect 10968 6273 10977 6307
rect 10977 6273 11011 6307
rect 11011 6273 11020 6307
rect 10968 6264 11020 6273
rect 17132 6264 17184 6316
rect 18236 6264 18288 6316
rect 19156 6307 19208 6316
rect 19156 6273 19165 6307
rect 19165 6273 19199 6307
rect 19199 6273 19208 6307
rect 19156 6264 19208 6273
rect 19248 6307 19300 6316
rect 19248 6273 19257 6307
rect 19257 6273 19291 6307
rect 19291 6273 19300 6307
rect 19248 6264 19300 6273
rect 19340 6307 19392 6316
rect 19340 6273 19349 6307
rect 19349 6273 19383 6307
rect 19383 6273 19392 6307
rect 19340 6264 19392 6273
rect 3976 6239 4028 6248
rect 3976 6205 3985 6239
rect 3985 6205 4019 6239
rect 4019 6205 4028 6239
rect 3976 6196 4028 6205
rect 8944 6239 8996 6248
rect 8944 6205 8953 6239
rect 8953 6205 8987 6239
rect 8987 6205 8996 6239
rect 8944 6196 8996 6205
rect 15476 6196 15528 6248
rect 19432 6196 19484 6248
rect 10140 6128 10192 6180
rect 10876 6128 10928 6180
rect 20352 6264 20404 6316
rect 23756 6375 23808 6384
rect 23756 6341 23765 6375
rect 23765 6341 23799 6375
rect 23799 6341 23808 6375
rect 23756 6332 23808 6341
rect 24584 6332 24636 6384
rect 25872 6332 25924 6384
rect 22744 6264 22796 6316
rect 23112 6307 23164 6316
rect 23112 6273 23121 6307
rect 23121 6273 23155 6307
rect 23155 6273 23164 6307
rect 23112 6264 23164 6273
rect 27068 6264 27120 6316
rect 35072 6332 35124 6384
rect 27620 6264 27672 6316
rect 29276 6307 29328 6316
rect 29276 6273 29285 6307
rect 29285 6273 29319 6307
rect 29319 6273 29328 6307
rect 29276 6264 29328 6273
rect 20168 6239 20220 6248
rect 20168 6205 20177 6239
rect 20177 6205 20211 6239
rect 20211 6205 20220 6239
rect 20168 6196 20220 6205
rect 20812 6239 20864 6248
rect 20812 6205 20821 6239
rect 20821 6205 20855 6239
rect 20855 6205 20864 6239
rect 20812 6196 20864 6205
rect 23480 6196 23532 6248
rect 24492 6196 24544 6248
rect 22560 6128 22612 6180
rect 23020 6128 23072 6180
rect 29184 6196 29236 6248
rect 30748 6264 30800 6316
rect 32312 6264 32364 6316
rect 30012 6239 30064 6248
rect 30012 6205 30021 6239
rect 30021 6205 30055 6239
rect 30055 6205 30064 6239
rect 30012 6196 30064 6205
rect 33876 6307 33928 6316
rect 33876 6273 33885 6307
rect 33885 6273 33919 6307
rect 33919 6273 33928 6307
rect 33876 6264 33928 6273
rect 34060 6264 34112 6316
rect 33692 6196 33744 6248
rect 35348 6264 35400 6316
rect 35440 6307 35492 6316
rect 35440 6273 35449 6307
rect 35449 6273 35483 6307
rect 35483 6273 35492 6307
rect 35440 6264 35492 6273
rect 35992 6264 36044 6316
rect 36452 6400 36504 6452
rect 37556 6400 37608 6452
rect 36268 6332 36320 6384
rect 34520 6196 34572 6248
rect 37372 6264 37424 6316
rect 37648 6307 37700 6316
rect 37648 6273 37657 6307
rect 37657 6273 37691 6307
rect 37691 6273 37700 6307
rect 37648 6264 37700 6273
rect 43720 6400 43772 6452
rect 38660 6307 38712 6316
rect 38660 6273 38669 6307
rect 38669 6273 38703 6307
rect 38703 6273 38712 6307
rect 38660 6264 38712 6273
rect 39028 6307 39080 6316
rect 39028 6273 39037 6307
rect 39037 6273 39071 6307
rect 39071 6273 39080 6307
rect 39028 6264 39080 6273
rect 37280 6196 37332 6248
rect 8300 6103 8352 6112
rect 8300 6069 8309 6103
rect 8309 6069 8343 6103
rect 8343 6069 8352 6103
rect 8300 6060 8352 6069
rect 9312 6103 9364 6112
rect 9312 6069 9321 6103
rect 9321 6069 9355 6103
rect 9355 6069 9364 6103
rect 9312 6060 9364 6069
rect 18328 6103 18380 6112
rect 18328 6069 18337 6103
rect 18337 6069 18371 6103
rect 18371 6069 18380 6103
rect 18328 6060 18380 6069
rect 20628 6060 20680 6112
rect 22468 6060 22520 6112
rect 24124 6103 24176 6112
rect 24124 6069 24133 6103
rect 24133 6069 24167 6103
rect 24167 6069 24176 6103
rect 24124 6060 24176 6069
rect 24860 6060 24912 6112
rect 29000 6060 29052 6112
rect 29092 6103 29144 6112
rect 29092 6069 29101 6103
rect 29101 6069 29135 6103
rect 29135 6069 29144 6103
rect 29092 6060 29144 6069
rect 29828 6103 29880 6112
rect 29828 6069 29837 6103
rect 29837 6069 29871 6103
rect 29871 6069 29880 6103
rect 29828 6060 29880 6069
rect 29920 6103 29972 6112
rect 29920 6069 29929 6103
rect 29929 6069 29963 6103
rect 29963 6069 29972 6103
rect 29920 6060 29972 6069
rect 33416 6060 33468 6112
rect 35624 6128 35676 6180
rect 34980 6060 35032 6112
rect 35348 6060 35400 6112
rect 35440 6060 35492 6112
rect 38568 6128 38620 6180
rect 40684 6239 40736 6248
rect 40684 6205 40693 6239
rect 40693 6205 40727 6239
rect 40727 6205 40736 6239
rect 41512 6307 41564 6316
rect 41512 6273 41521 6307
rect 41521 6273 41555 6307
rect 41555 6273 41564 6307
rect 41512 6264 41564 6273
rect 40684 6196 40736 6205
rect 40960 6196 41012 6248
rect 41512 6128 41564 6180
rect 36268 6103 36320 6112
rect 36268 6069 36277 6103
rect 36277 6069 36311 6103
rect 36311 6069 36320 6103
rect 36268 6060 36320 6069
rect 36912 6060 36964 6112
rect 38752 6060 38804 6112
rect 42616 6103 42668 6112
rect 42616 6069 42625 6103
rect 42625 6069 42659 6103
rect 42659 6069 42668 6103
rect 42616 6060 42668 6069
rect 6423 5958 6475 6010
rect 6487 5958 6539 6010
rect 6551 5958 6603 6010
rect 6615 5958 6667 6010
rect 6679 5958 6731 6010
rect 17370 5958 17422 6010
rect 17434 5958 17486 6010
rect 17498 5958 17550 6010
rect 17562 5958 17614 6010
rect 17626 5958 17678 6010
rect 28317 5958 28369 6010
rect 28381 5958 28433 6010
rect 28445 5958 28497 6010
rect 28509 5958 28561 6010
rect 28573 5958 28625 6010
rect 39264 5958 39316 6010
rect 39328 5958 39380 6010
rect 39392 5958 39444 6010
rect 39456 5958 39508 6010
rect 39520 5958 39572 6010
rect 940 5856 992 5908
rect 5264 5856 5316 5908
rect 11796 5856 11848 5908
rect 2964 5695 3016 5704
rect 2964 5661 2973 5695
rect 2973 5661 3007 5695
rect 3007 5661 3016 5695
rect 2964 5652 3016 5661
rect 3976 5695 4028 5704
rect 3976 5661 3985 5695
rect 3985 5661 4019 5695
rect 4019 5661 4028 5695
rect 3976 5652 4028 5661
rect 4712 5652 4764 5704
rect 5448 5652 5500 5704
rect 8944 5788 8996 5840
rect 15476 5856 15528 5908
rect 18144 5856 18196 5908
rect 19340 5856 19392 5908
rect 20168 5856 20220 5908
rect 20352 5856 20404 5908
rect 23020 5899 23072 5908
rect 23020 5865 23029 5899
rect 23029 5865 23063 5899
rect 23063 5865 23072 5899
rect 23020 5856 23072 5865
rect 23112 5856 23164 5908
rect 16120 5788 16172 5840
rect 17960 5788 18012 5840
rect 19156 5788 19208 5840
rect 15752 5720 15804 5772
rect 18236 5720 18288 5772
rect 6000 5695 6052 5704
rect 6000 5661 6009 5695
rect 6009 5661 6043 5695
rect 6043 5661 6052 5695
rect 6000 5652 6052 5661
rect 8392 5695 8444 5704
rect 8392 5661 8401 5695
rect 8401 5661 8435 5695
rect 8435 5661 8444 5695
rect 8392 5652 8444 5661
rect 12532 5652 12584 5704
rect 12624 5695 12676 5704
rect 12624 5661 12633 5695
rect 12633 5661 12667 5695
rect 12667 5661 12676 5695
rect 12624 5652 12676 5661
rect 13360 5652 13412 5704
rect 13544 5695 13596 5704
rect 13544 5661 13553 5695
rect 13553 5661 13587 5695
rect 13587 5661 13596 5695
rect 13544 5652 13596 5661
rect 13820 5652 13872 5704
rect 14924 5652 14976 5704
rect 16304 5695 16356 5704
rect 16304 5661 16313 5695
rect 16313 5661 16347 5695
rect 16347 5661 16356 5695
rect 16304 5652 16356 5661
rect 17684 5695 17736 5704
rect 17684 5661 17693 5695
rect 17693 5661 17727 5695
rect 17727 5661 17736 5695
rect 17684 5652 17736 5661
rect 17776 5652 17828 5704
rect 6920 5584 6972 5636
rect 14556 5627 14608 5636
rect 6184 5559 6236 5568
rect 6184 5525 6193 5559
rect 6193 5525 6227 5559
rect 6227 5525 6236 5559
rect 6184 5516 6236 5525
rect 7196 5516 7248 5568
rect 12716 5559 12768 5568
rect 12716 5525 12725 5559
rect 12725 5525 12759 5559
rect 12759 5525 12768 5559
rect 12716 5516 12768 5525
rect 12808 5516 12860 5568
rect 14556 5593 14590 5627
rect 14590 5593 14608 5627
rect 14556 5584 14608 5593
rect 16580 5584 16632 5636
rect 14464 5516 14516 5568
rect 15844 5516 15896 5568
rect 18604 5695 18656 5704
rect 18604 5661 18613 5695
rect 18613 5661 18647 5695
rect 18647 5661 18656 5695
rect 18604 5652 18656 5661
rect 23388 5788 23440 5840
rect 24584 5899 24636 5908
rect 24584 5865 24593 5899
rect 24593 5865 24627 5899
rect 24627 5865 24636 5899
rect 24584 5856 24636 5865
rect 26056 5899 26108 5908
rect 26056 5865 26065 5899
rect 26065 5865 26099 5899
rect 26099 5865 26108 5899
rect 26056 5856 26108 5865
rect 27620 5899 27672 5908
rect 27620 5865 27629 5899
rect 27629 5865 27663 5899
rect 27663 5865 27672 5899
rect 27620 5856 27672 5865
rect 29276 5856 29328 5908
rect 34244 5856 34296 5908
rect 34336 5899 34388 5908
rect 34336 5865 34345 5899
rect 34345 5865 34379 5899
rect 34379 5865 34388 5899
rect 34336 5856 34388 5865
rect 19524 5720 19576 5772
rect 22008 5720 22060 5772
rect 18328 5584 18380 5636
rect 19616 5627 19668 5636
rect 19616 5593 19625 5627
rect 19625 5593 19659 5627
rect 19659 5593 19668 5627
rect 19616 5584 19668 5593
rect 20628 5695 20680 5704
rect 20628 5661 20637 5695
rect 20637 5661 20671 5695
rect 20671 5661 20680 5695
rect 20628 5652 20680 5661
rect 20720 5695 20772 5704
rect 20720 5661 20729 5695
rect 20729 5661 20763 5695
rect 20763 5661 20772 5695
rect 20720 5652 20772 5661
rect 21180 5652 21232 5704
rect 20812 5516 20864 5568
rect 20904 5516 20956 5568
rect 24124 5652 24176 5704
rect 29736 5788 29788 5840
rect 24860 5652 24912 5704
rect 25044 5695 25096 5704
rect 25044 5661 25053 5695
rect 25053 5661 25087 5695
rect 25087 5661 25096 5695
rect 25044 5652 25096 5661
rect 25872 5695 25924 5704
rect 25872 5661 25881 5695
rect 25881 5661 25915 5695
rect 25915 5661 25924 5695
rect 25872 5652 25924 5661
rect 26240 5652 26292 5704
rect 29920 5720 29972 5772
rect 30656 5720 30708 5772
rect 35164 5856 35216 5908
rect 35532 5856 35584 5908
rect 36544 5856 36596 5908
rect 37188 5856 37240 5908
rect 37280 5856 37332 5908
rect 40316 5856 40368 5908
rect 40500 5788 40552 5840
rect 37648 5720 37700 5772
rect 29828 5652 29880 5704
rect 30380 5695 30432 5704
rect 30380 5661 30389 5695
rect 30389 5661 30423 5695
rect 30423 5661 30432 5695
rect 30380 5652 30432 5661
rect 30472 5652 30524 5704
rect 34060 5695 34112 5704
rect 34060 5661 34069 5695
rect 34069 5661 34103 5695
rect 34103 5661 34112 5695
rect 34060 5652 34112 5661
rect 34428 5652 34480 5704
rect 34796 5652 34848 5704
rect 38016 5695 38068 5704
rect 38016 5661 38025 5695
rect 38025 5661 38059 5695
rect 38059 5661 38068 5695
rect 38016 5652 38068 5661
rect 39028 5720 39080 5772
rect 40776 5763 40828 5772
rect 40776 5729 40785 5763
rect 40785 5729 40819 5763
rect 40819 5729 40828 5763
rect 40776 5720 40828 5729
rect 22468 5559 22520 5568
rect 22468 5525 22477 5559
rect 22477 5525 22511 5559
rect 22511 5525 22520 5559
rect 22468 5516 22520 5525
rect 34888 5584 34940 5636
rect 35348 5584 35400 5636
rect 36728 5627 36780 5636
rect 36728 5593 36737 5627
rect 36737 5593 36771 5627
rect 36771 5593 36780 5627
rect 36728 5584 36780 5593
rect 36912 5627 36964 5636
rect 36912 5593 36937 5627
rect 36937 5593 36964 5627
rect 36912 5584 36964 5593
rect 37372 5584 37424 5636
rect 38568 5652 38620 5704
rect 38660 5652 38712 5704
rect 42616 5652 42668 5704
rect 24308 5516 24360 5568
rect 25228 5516 25280 5568
rect 29184 5516 29236 5568
rect 30748 5559 30800 5568
rect 30748 5525 30757 5559
rect 30757 5525 30791 5559
rect 30791 5525 30800 5559
rect 30748 5516 30800 5525
rect 37096 5559 37148 5568
rect 37096 5525 37105 5559
rect 37105 5525 37139 5559
rect 37139 5525 37148 5559
rect 37096 5516 37148 5525
rect 43904 5584 43956 5636
rect 38660 5559 38712 5568
rect 38660 5525 38669 5559
rect 38669 5525 38703 5559
rect 38703 5525 38712 5559
rect 38660 5516 38712 5525
rect 41696 5516 41748 5568
rect 11896 5414 11948 5466
rect 11960 5414 12012 5466
rect 12024 5414 12076 5466
rect 12088 5414 12140 5466
rect 12152 5414 12204 5466
rect 22843 5414 22895 5466
rect 22907 5414 22959 5466
rect 22971 5414 23023 5466
rect 23035 5414 23087 5466
rect 23099 5414 23151 5466
rect 33790 5414 33842 5466
rect 33854 5414 33906 5466
rect 33918 5414 33970 5466
rect 33982 5414 34034 5466
rect 34046 5414 34098 5466
rect 44737 5414 44789 5466
rect 44801 5414 44853 5466
rect 44865 5414 44917 5466
rect 44929 5414 44981 5466
rect 44993 5414 45045 5466
rect 4344 5355 4396 5364
rect 4344 5321 4353 5355
rect 4353 5321 4387 5355
rect 4387 5321 4396 5355
rect 4344 5312 4396 5321
rect 4436 5355 4488 5364
rect 4436 5321 4445 5355
rect 4445 5321 4479 5355
rect 4479 5321 4488 5355
rect 4436 5312 4488 5321
rect 10876 5355 10928 5364
rect 10876 5321 10885 5355
rect 10885 5321 10919 5355
rect 10919 5321 10928 5355
rect 10876 5312 10928 5321
rect 13268 5312 13320 5364
rect 7196 5287 7248 5296
rect 7196 5253 7205 5287
rect 7205 5253 7239 5287
rect 7239 5253 7248 5287
rect 7196 5244 7248 5253
rect 4712 5176 4764 5228
rect 5264 5176 5316 5228
rect 940 5108 992 5160
rect 1860 5151 1912 5160
rect 1860 5117 1869 5151
rect 1869 5117 1903 5151
rect 1903 5117 1912 5151
rect 1860 5108 1912 5117
rect 5080 5108 5132 5160
rect 8300 5176 8352 5228
rect 9404 5244 9456 5296
rect 10416 5244 10468 5296
rect 12808 5287 12860 5296
rect 12808 5253 12817 5287
rect 12817 5253 12851 5287
rect 12851 5253 12860 5287
rect 12808 5244 12860 5253
rect 12716 5176 12768 5228
rect 13452 5176 13504 5228
rect 13728 5244 13780 5296
rect 15844 5244 15896 5296
rect 15752 5219 15804 5228
rect 15752 5185 15761 5219
rect 15761 5185 15795 5219
rect 15795 5185 15804 5219
rect 15752 5176 15804 5185
rect 13820 5151 13872 5160
rect 13820 5117 13829 5151
rect 13829 5117 13863 5151
rect 13863 5117 13872 5151
rect 13820 5108 13872 5117
rect 17960 5312 18012 5364
rect 20536 5312 20588 5364
rect 16948 5287 17000 5296
rect 16948 5253 16957 5287
rect 16957 5253 16991 5287
rect 16991 5253 17000 5287
rect 16948 5244 17000 5253
rect 17684 5176 17736 5228
rect 18512 5244 18564 5296
rect 18236 5219 18288 5228
rect 18236 5185 18245 5219
rect 18245 5185 18279 5219
rect 18279 5185 18288 5219
rect 18236 5176 18288 5185
rect 18880 5176 18932 5228
rect 15844 5151 15896 5160
rect 15844 5117 15853 5151
rect 15853 5117 15887 5151
rect 15887 5117 15896 5151
rect 15844 5108 15896 5117
rect 15936 5108 15988 5160
rect 16120 5108 16172 5160
rect 16948 5108 17000 5160
rect 17960 5151 18012 5160
rect 17960 5117 17969 5151
rect 17969 5117 18003 5151
rect 18003 5117 18012 5151
rect 17960 5108 18012 5117
rect 18420 5108 18472 5160
rect 19708 5244 19760 5296
rect 20444 5244 20496 5296
rect 4528 5040 4580 5092
rect 7196 4972 7248 5024
rect 12164 5015 12216 5024
rect 12164 4981 12173 5015
rect 12173 4981 12207 5015
rect 12207 4981 12216 5015
rect 12164 4972 12216 4981
rect 12900 4972 12952 5024
rect 18604 5040 18656 5092
rect 17776 4972 17828 5024
rect 18512 4972 18564 5024
rect 19064 4972 19116 5024
rect 22468 5312 22520 5364
rect 22744 5355 22796 5364
rect 22744 5321 22753 5355
rect 22753 5321 22787 5355
rect 22787 5321 22796 5355
rect 22744 5312 22796 5321
rect 20904 5244 20956 5296
rect 24032 5312 24084 5364
rect 28724 5312 28776 5364
rect 20996 5176 21048 5228
rect 23388 5244 23440 5296
rect 21180 5108 21232 5160
rect 23940 5219 23992 5228
rect 23940 5185 23949 5219
rect 23949 5185 23983 5219
rect 23983 5185 23992 5219
rect 23940 5176 23992 5185
rect 29000 5244 29052 5296
rect 24308 5219 24360 5228
rect 24308 5185 24317 5219
rect 24317 5185 24351 5219
rect 24351 5185 24360 5219
rect 24308 5176 24360 5185
rect 25228 5219 25280 5228
rect 25228 5185 25237 5219
rect 25237 5185 25271 5219
rect 25271 5185 25280 5219
rect 25228 5176 25280 5185
rect 25320 5219 25372 5228
rect 25320 5185 25329 5219
rect 25329 5185 25363 5219
rect 25363 5185 25372 5219
rect 25320 5176 25372 5185
rect 19800 5040 19852 5092
rect 20168 5015 20220 5024
rect 20168 4981 20177 5015
rect 20177 4981 20211 5015
rect 20211 4981 20220 5015
rect 20168 4972 20220 4981
rect 21364 5015 21416 5024
rect 21364 4981 21373 5015
rect 21373 4981 21407 5015
rect 21407 4981 21416 5015
rect 22560 5040 22612 5092
rect 27344 5176 27396 5228
rect 33416 5176 33468 5228
rect 37556 5287 37608 5296
rect 37556 5253 37565 5287
rect 37565 5253 37599 5287
rect 37599 5253 37608 5287
rect 37556 5244 37608 5253
rect 27160 5108 27212 5160
rect 21364 4972 21416 4981
rect 23940 4972 23992 5024
rect 25872 4972 25924 5024
rect 29092 5108 29144 5160
rect 29828 5151 29880 5160
rect 29828 5117 29837 5151
rect 29837 5117 29871 5151
rect 29871 5117 29880 5151
rect 29828 5108 29880 5117
rect 35164 5176 35216 5228
rect 35532 5176 35584 5228
rect 37188 5176 37240 5228
rect 38660 5244 38712 5296
rect 38752 5287 38804 5296
rect 38752 5253 38786 5287
rect 38786 5253 38804 5287
rect 38752 5244 38804 5253
rect 41512 5312 41564 5364
rect 41420 5176 41472 5228
rect 41696 5219 41748 5228
rect 41696 5185 41705 5219
rect 41705 5185 41739 5219
rect 41739 5185 41748 5219
rect 41696 5176 41748 5185
rect 42800 5219 42852 5228
rect 42800 5185 42809 5219
rect 42809 5185 42843 5219
rect 42843 5185 42852 5219
rect 42800 5176 42852 5185
rect 38568 5151 38620 5160
rect 38568 5117 38577 5151
rect 38577 5117 38611 5151
rect 38611 5117 38620 5151
rect 38568 5108 38620 5117
rect 44640 5108 44692 5160
rect 29368 4972 29420 5024
rect 30748 4972 30800 5024
rect 34980 5015 35032 5024
rect 34980 4981 34989 5015
rect 34989 4981 35023 5015
rect 35023 4981 35032 5015
rect 34980 4972 35032 4981
rect 38936 5083 38988 5092
rect 38936 5049 38945 5083
rect 38945 5049 38979 5083
rect 38979 5049 38988 5083
rect 38936 5040 38988 5049
rect 37188 4972 37240 5024
rect 6423 4870 6475 4922
rect 6487 4870 6539 4922
rect 6551 4870 6603 4922
rect 6615 4870 6667 4922
rect 6679 4870 6731 4922
rect 17370 4870 17422 4922
rect 17434 4870 17486 4922
rect 17498 4870 17550 4922
rect 17562 4870 17614 4922
rect 17626 4870 17678 4922
rect 28317 4870 28369 4922
rect 28381 4870 28433 4922
rect 28445 4870 28497 4922
rect 28509 4870 28561 4922
rect 28573 4870 28625 4922
rect 39264 4870 39316 4922
rect 39328 4870 39380 4922
rect 39392 4870 39444 4922
rect 39456 4870 39508 4922
rect 39520 4870 39572 4922
rect 10416 4811 10468 4820
rect 10416 4777 10425 4811
rect 10425 4777 10459 4811
rect 10459 4777 10468 4811
rect 10416 4768 10468 4777
rect 1860 4700 1912 4752
rect 13360 4768 13412 4820
rect 16304 4768 16356 4820
rect 13268 4700 13320 4752
rect 4344 4632 4396 4684
rect 4712 4607 4764 4616
rect 4712 4573 4721 4607
rect 4721 4573 4755 4607
rect 4755 4573 4764 4607
rect 4712 4564 4764 4573
rect 11796 4675 11848 4684
rect 11796 4641 11805 4675
rect 11805 4641 11839 4675
rect 11839 4641 11848 4675
rect 11796 4632 11848 4641
rect 12716 4632 12768 4684
rect 9864 4607 9916 4616
rect 9864 4573 9873 4607
rect 9873 4573 9907 4607
rect 9907 4573 9916 4607
rect 9864 4564 9916 4573
rect 14464 4607 14516 4616
rect 14464 4573 14473 4607
rect 14473 4573 14507 4607
rect 14507 4573 14516 4607
rect 14464 4564 14516 4573
rect 15936 4632 15988 4684
rect 18420 4768 18472 4820
rect 18880 4811 18932 4820
rect 18880 4777 18889 4811
rect 18889 4777 18923 4811
rect 18923 4777 18932 4811
rect 18880 4768 18932 4777
rect 21180 4811 21232 4820
rect 21180 4777 21189 4811
rect 21189 4777 21223 4811
rect 21223 4777 21232 4811
rect 21180 4768 21232 4777
rect 23756 4768 23808 4820
rect 24584 4768 24636 4820
rect 25320 4768 25372 4820
rect 16580 4632 16632 4684
rect 18144 4632 18196 4684
rect 23940 4743 23992 4752
rect 23940 4709 23949 4743
rect 23949 4709 23983 4743
rect 23983 4709 23992 4743
rect 27344 4811 27396 4820
rect 27344 4777 27353 4811
rect 27353 4777 27387 4811
rect 27387 4777 27396 4811
rect 27344 4768 27396 4777
rect 35532 4768 35584 4820
rect 38016 4768 38068 4820
rect 38568 4768 38620 4820
rect 23940 4700 23992 4709
rect 23664 4632 23716 4684
rect 24492 4632 24544 4684
rect 12164 4496 12216 4548
rect 13544 4496 13596 4548
rect 21824 4607 21876 4616
rect 21824 4573 21833 4607
rect 21833 4573 21867 4607
rect 21867 4573 21876 4607
rect 21824 4564 21876 4573
rect 17408 4539 17460 4548
rect 17408 4505 17417 4539
rect 17417 4505 17451 4539
rect 17451 4505 17460 4539
rect 17408 4496 17460 4505
rect 19432 4496 19484 4548
rect 20720 4496 20772 4548
rect 24032 4607 24084 4616
rect 24032 4573 24041 4607
rect 24041 4573 24075 4607
rect 24075 4573 24084 4607
rect 24032 4564 24084 4573
rect 24584 4607 24636 4616
rect 24584 4573 24593 4607
rect 24593 4573 24627 4607
rect 24627 4573 24636 4607
rect 24584 4564 24636 4573
rect 30012 4700 30064 4752
rect 29368 4632 29420 4684
rect 29000 4564 29052 4616
rect 30564 4607 30616 4616
rect 30564 4573 30573 4607
rect 30573 4573 30607 4607
rect 30607 4573 30616 4607
rect 30564 4564 30616 4573
rect 36268 4564 36320 4616
rect 36728 4607 36780 4616
rect 36728 4573 36737 4607
rect 36737 4573 36771 4607
rect 36771 4573 36780 4607
rect 36728 4564 36780 4573
rect 37188 4632 37240 4684
rect 37464 4564 37516 4616
rect 44180 4632 44232 4684
rect 25872 4539 25924 4548
rect 25872 4505 25881 4539
rect 25881 4505 25915 4539
rect 25915 4505 25924 4539
rect 25872 4496 25924 4505
rect 26884 4496 26936 4548
rect 5632 4428 5684 4480
rect 15108 4471 15160 4480
rect 15108 4437 15117 4471
rect 15117 4437 15151 4471
rect 15151 4437 15160 4471
rect 15108 4428 15160 4437
rect 24032 4428 24084 4480
rect 24124 4428 24176 4480
rect 25412 4428 25464 4480
rect 29736 4471 29788 4480
rect 29736 4437 29745 4471
rect 29745 4437 29779 4471
rect 29779 4437 29788 4471
rect 29736 4428 29788 4437
rect 30380 4471 30432 4480
rect 30380 4437 30389 4471
rect 30389 4437 30423 4471
rect 30423 4437 30432 4471
rect 30380 4428 30432 4437
rect 11896 4326 11948 4378
rect 11960 4326 12012 4378
rect 12024 4326 12076 4378
rect 12088 4326 12140 4378
rect 12152 4326 12204 4378
rect 22843 4326 22895 4378
rect 22907 4326 22959 4378
rect 22971 4326 23023 4378
rect 23035 4326 23087 4378
rect 23099 4326 23151 4378
rect 33790 4326 33842 4378
rect 33854 4326 33906 4378
rect 33918 4326 33970 4378
rect 33982 4326 34034 4378
rect 34046 4326 34098 4378
rect 44737 4326 44789 4378
rect 44801 4326 44853 4378
rect 44865 4326 44917 4378
rect 44929 4326 44981 4378
rect 44993 4326 45045 4378
rect 12716 4267 12768 4276
rect 12716 4233 12725 4267
rect 12725 4233 12759 4267
rect 12759 4233 12768 4267
rect 12716 4224 12768 4233
rect 13820 4224 13872 4276
rect 16948 4224 17000 4276
rect 17408 4224 17460 4276
rect 18604 4267 18656 4276
rect 18604 4233 18613 4267
rect 18613 4233 18647 4267
rect 18647 4233 18656 4267
rect 18604 4224 18656 4233
rect 20168 4267 20220 4276
rect 20168 4233 20198 4267
rect 20198 4233 20220 4267
rect 20168 4224 20220 4233
rect 23756 4224 23808 4276
rect 25412 4267 25464 4276
rect 25412 4233 25421 4267
rect 25421 4233 25455 4267
rect 25455 4233 25464 4267
rect 25412 4224 25464 4233
rect 29736 4156 29788 4208
rect 9864 4088 9916 4140
rect 12900 4131 12952 4140
rect 12900 4097 12909 4131
rect 12909 4097 12943 4131
rect 12943 4097 12952 4131
rect 12900 4088 12952 4097
rect 15108 4088 15160 4140
rect 16856 4088 16908 4140
rect 17776 4088 17828 4140
rect 19064 4088 19116 4140
rect 19800 4088 19852 4140
rect 8484 3952 8536 4004
rect 16580 3884 16632 3936
rect 19616 3884 19668 3936
rect 21364 4020 21416 4072
rect 21824 3952 21876 4004
rect 20628 3884 20680 3936
rect 23664 4131 23716 4140
rect 23664 4097 23673 4131
rect 23673 4097 23707 4131
rect 23707 4097 23716 4131
rect 23664 4088 23716 4097
rect 26056 4131 26108 4140
rect 26056 4097 26065 4131
rect 26065 4097 26099 4131
rect 26099 4097 26108 4131
rect 26056 4088 26108 4097
rect 23940 4063 23992 4072
rect 23940 4029 23949 4063
rect 23949 4029 23983 4063
rect 23983 4029 23992 4063
rect 23940 4020 23992 4029
rect 25964 4020 26016 4072
rect 29000 4088 29052 4140
rect 29368 4131 29420 4140
rect 29368 4097 29377 4131
rect 29377 4097 29411 4131
rect 29411 4097 29420 4131
rect 29368 4088 29420 4097
rect 31208 4088 31260 4140
rect 30380 4020 30432 4072
rect 41420 4020 41472 4072
rect 24952 3884 25004 3936
rect 26976 3884 27028 3936
rect 6423 3782 6475 3834
rect 6487 3782 6539 3834
rect 6551 3782 6603 3834
rect 6615 3782 6667 3834
rect 6679 3782 6731 3834
rect 17370 3782 17422 3834
rect 17434 3782 17486 3834
rect 17498 3782 17550 3834
rect 17562 3782 17614 3834
rect 17626 3782 17678 3834
rect 28317 3782 28369 3834
rect 28381 3782 28433 3834
rect 28445 3782 28497 3834
rect 28509 3782 28561 3834
rect 28573 3782 28625 3834
rect 39264 3782 39316 3834
rect 39328 3782 39380 3834
rect 39392 3782 39444 3834
rect 39456 3782 39508 3834
rect 39520 3782 39572 3834
rect 19432 3723 19484 3732
rect 19432 3689 19441 3723
rect 19441 3689 19475 3723
rect 19475 3689 19484 3723
rect 19432 3680 19484 3689
rect 20720 3680 20772 3732
rect 23940 3680 23992 3732
rect 26056 3680 26108 3732
rect 26884 3680 26936 3732
rect 30564 3612 30616 3664
rect 6276 3587 6328 3596
rect 6276 3553 6285 3587
rect 6285 3553 6319 3587
rect 6319 3553 6328 3587
rect 6276 3544 6328 3553
rect 30012 3587 30064 3596
rect 30012 3553 30021 3587
rect 30021 3553 30055 3587
rect 30055 3553 30064 3587
rect 30012 3544 30064 3553
rect 940 3476 992 3528
rect 5632 3519 5684 3528
rect 5632 3485 5641 3519
rect 5641 3485 5675 3519
rect 5675 3485 5684 3519
rect 5632 3476 5684 3485
rect 13728 3476 13780 3528
rect 14832 3476 14884 3528
rect 15384 3519 15436 3528
rect 15384 3485 15393 3519
rect 15393 3485 15427 3519
rect 15427 3485 15436 3519
rect 15384 3476 15436 3485
rect 16120 3476 16172 3528
rect 16212 3519 16264 3528
rect 16212 3485 16221 3519
rect 16221 3485 16255 3519
rect 16255 3485 16264 3519
rect 16212 3476 16264 3485
rect 18144 3519 18196 3528
rect 18144 3485 18153 3519
rect 18153 3485 18187 3519
rect 18187 3485 18196 3519
rect 18144 3476 18196 3485
rect 19616 3519 19668 3528
rect 19616 3485 19625 3519
rect 19625 3485 19659 3519
rect 19659 3485 19668 3519
rect 19616 3476 19668 3485
rect 20628 3519 20680 3528
rect 20628 3485 20637 3519
rect 20637 3485 20671 3519
rect 20671 3485 20680 3519
rect 20628 3476 20680 3485
rect 24032 3519 24084 3528
rect 24032 3485 24041 3519
rect 24041 3485 24075 3519
rect 24075 3485 24084 3519
rect 24032 3476 24084 3485
rect 24952 3476 25004 3528
rect 26976 3519 27028 3528
rect 26976 3485 26985 3519
rect 26985 3485 27019 3519
rect 27019 3485 27028 3519
rect 26976 3476 27028 3485
rect 31208 3476 31260 3528
rect 44640 3476 44692 3528
rect 16580 3408 16632 3460
rect 18052 3408 18104 3460
rect 23296 3408 23348 3460
rect 33508 3408 33560 3460
rect 13636 3383 13688 3392
rect 13636 3349 13645 3383
rect 13645 3349 13679 3383
rect 13679 3349 13688 3383
rect 13636 3340 13688 3349
rect 15200 3383 15252 3392
rect 15200 3349 15209 3383
rect 15209 3349 15243 3383
rect 15243 3349 15252 3383
rect 15200 3340 15252 3349
rect 17776 3340 17828 3392
rect 11896 3238 11948 3290
rect 11960 3238 12012 3290
rect 12024 3238 12076 3290
rect 12088 3238 12140 3290
rect 12152 3238 12204 3290
rect 22843 3238 22895 3290
rect 22907 3238 22959 3290
rect 22971 3238 23023 3290
rect 23035 3238 23087 3290
rect 23099 3238 23151 3290
rect 33790 3238 33842 3290
rect 33854 3238 33906 3290
rect 33918 3238 33970 3290
rect 33982 3238 34034 3290
rect 34046 3238 34098 3290
rect 44737 3238 44789 3290
rect 44801 3238 44853 3290
rect 44865 3238 44917 3290
rect 44929 3238 44981 3290
rect 44993 3238 45045 3290
rect 9312 3136 9364 3188
rect 15200 3068 15252 3120
rect 16120 3136 16172 3188
rect 7196 3043 7248 3052
rect 7196 3009 7205 3043
rect 7205 3009 7239 3043
rect 7239 3009 7248 3043
rect 7196 3000 7248 3009
rect 13636 3043 13688 3052
rect 13636 3009 13645 3043
rect 13645 3009 13679 3043
rect 13679 3009 13688 3043
rect 13636 3000 13688 3009
rect 14832 3043 14884 3052
rect 14832 3009 14841 3043
rect 14841 3009 14875 3043
rect 14875 3009 14884 3043
rect 14832 3000 14884 3009
rect 16212 3000 16264 3052
rect 17776 3000 17828 3052
rect 18052 3043 18104 3052
rect 18052 3009 18061 3043
rect 18061 3009 18095 3043
rect 18095 3009 18104 3043
rect 18052 3000 18104 3009
rect 9680 2932 9732 2984
rect 17132 2932 17184 2984
rect 19800 3111 19852 3120
rect 19800 3077 19809 3111
rect 19809 3077 19843 3111
rect 19843 3077 19852 3111
rect 19800 3068 19852 3077
rect 940 2796 992 2848
rect 18880 2796 18932 2848
rect 22652 3000 22704 3052
rect 44180 3179 44232 3188
rect 44180 3145 44189 3179
rect 44189 3145 44223 3179
rect 44223 3145 44232 3179
rect 44180 3136 44232 3145
rect 45100 3000 45152 3052
rect 22560 2932 22612 2984
rect 35440 2975 35492 2984
rect 35440 2941 35449 2975
rect 35449 2941 35483 2975
rect 35483 2941 35492 2975
rect 35440 2932 35492 2941
rect 6423 2694 6475 2746
rect 6487 2694 6539 2746
rect 6551 2694 6603 2746
rect 6615 2694 6667 2746
rect 6679 2694 6731 2746
rect 17370 2694 17422 2746
rect 17434 2694 17486 2746
rect 17498 2694 17550 2746
rect 17562 2694 17614 2746
rect 17626 2694 17678 2746
rect 28317 2694 28369 2746
rect 28381 2694 28433 2746
rect 28445 2694 28497 2746
rect 28509 2694 28561 2746
rect 28573 2694 28625 2746
rect 39264 2694 39316 2746
rect 39328 2694 39380 2746
rect 39392 2694 39444 2746
rect 39456 2694 39508 2746
rect 39520 2694 39572 2746
rect 12808 2592 12860 2644
rect 15384 2592 15436 2644
rect 17132 2592 17184 2644
rect 17868 2592 17920 2644
rect 16120 2524 16172 2576
rect 18880 2524 18932 2576
rect 20 2456 72 2508
rect 1308 2388 1360 2440
rect 4160 2431 4212 2440
rect 4160 2397 4169 2431
rect 4169 2397 4203 2431
rect 4203 2397 4212 2431
rect 4160 2388 4212 2397
rect 4528 2388 4580 2440
rect 7748 2388 7800 2440
rect 11060 2388 11112 2440
rect 12900 2388 12952 2440
rect 18144 2456 18196 2508
rect 27528 2635 27580 2644
rect 27528 2601 27537 2635
rect 27537 2601 27571 2635
rect 27571 2601 27580 2635
rect 27528 2592 27580 2601
rect 32496 2635 32548 2644
rect 32496 2601 32505 2635
rect 32505 2601 32539 2635
rect 32539 2601 32548 2635
rect 32496 2592 32548 2601
rect 37464 2635 37516 2644
rect 37464 2601 37473 2635
rect 37473 2601 37507 2635
rect 37507 2601 37516 2635
rect 37464 2592 37516 2601
rect 43904 2635 43956 2644
rect 43904 2601 43913 2635
rect 43913 2601 43947 2635
rect 43947 2601 43956 2635
rect 43904 2592 43956 2601
rect 16856 2431 16908 2440
rect 16856 2397 16865 2431
rect 16865 2397 16899 2431
rect 16899 2397 16908 2431
rect 16856 2388 16908 2397
rect 17408 2388 17460 2440
rect 19340 2388 19392 2440
rect 20720 2388 20772 2440
rect 23848 2388 23900 2440
rect 25780 2388 25832 2440
rect 29000 2388 29052 2440
rect 30380 2388 30432 2440
rect 37648 2431 37700 2440
rect 37648 2397 37657 2431
rect 37657 2397 37691 2431
rect 37691 2397 37700 2431
rect 37648 2388 37700 2397
rect 38660 2388 38712 2440
rect 40040 2388 40092 2440
rect 43812 2388 43864 2440
rect 27068 2320 27120 2372
rect 32220 2320 32272 2372
rect 41880 2320 41932 2372
rect 30656 2252 30708 2304
rect 11896 2150 11948 2202
rect 11960 2150 12012 2202
rect 12024 2150 12076 2202
rect 12088 2150 12140 2202
rect 12152 2150 12204 2202
rect 22843 2150 22895 2202
rect 22907 2150 22959 2202
rect 22971 2150 23023 2202
rect 23035 2150 23087 2202
rect 23099 2150 23151 2202
rect 33790 2150 33842 2202
rect 33854 2150 33906 2202
rect 33918 2150 33970 2202
rect 33982 2150 34034 2202
rect 34046 2150 34098 2202
rect 44737 2150 44789 2202
rect 44801 2150 44853 2202
rect 44865 2150 44917 2202
rect 44929 2150 44981 2202
rect 44993 2150 45045 2202
rect 3240 892 3292 944
rect 4160 892 4212 944
rect 36728 892 36780 944
rect 37648 892 37700 944
<< metal2 >>
rect -10 19200 102 20000
rect 1278 19200 1390 20000
rect 3210 19200 3322 20000
rect 4498 19200 4610 20000
rect 6430 19200 6542 20000
rect 7718 19200 7830 20000
rect 9650 19200 9762 20000
rect 10938 19200 11050 20000
rect 12870 19200 12982 20000
rect 14158 19200 14270 20000
rect 16090 19200 16202 20000
rect 17378 19200 17490 20000
rect 19310 19200 19422 20000
rect 20598 19200 20710 20000
rect 22530 19200 22642 20000
rect 23818 19200 23930 20000
rect 25750 19200 25862 20000
rect 27682 19200 27794 20000
rect 28970 19200 29082 20000
rect 30902 19200 31014 20000
rect 32190 19200 32302 20000
rect 34122 19200 34234 20000
rect 35410 19200 35522 20000
rect 37342 19200 37454 20000
rect 38630 19200 38742 20000
rect 40562 19200 40674 20000
rect 41850 19200 41962 20000
rect 43782 19200 43894 20000
rect 45070 19200 45182 20000
rect 32 16590 60 19200
rect 1030 18456 1086 18465
rect 1030 18391 1086 18400
rect 940 17264 992 17270
rect 940 17206 992 17212
rect 952 17105 980 17206
rect 938 17096 994 17105
rect 938 17031 994 17040
rect 20 16584 72 16590
rect 20 16526 72 16532
rect 1044 16114 1072 18391
rect 1320 17202 1348 19200
rect 3252 17270 3280 19200
rect 3240 17264 3292 17270
rect 3240 17206 3292 17212
rect 4540 17202 4568 19200
rect 6472 17202 6500 19200
rect 7760 17202 7788 19200
rect 9692 17202 9720 19200
rect 10980 19122 11008 19200
rect 10980 19094 11100 19122
rect 11072 17270 11100 19094
rect 11896 17436 12204 17445
rect 11896 17434 11902 17436
rect 11958 17434 11982 17436
rect 12038 17434 12062 17436
rect 12118 17434 12142 17436
rect 12198 17434 12204 17436
rect 11958 17382 11960 17434
rect 12140 17382 12142 17434
rect 11896 17380 11902 17382
rect 11958 17380 11982 17382
rect 12038 17380 12062 17382
rect 12118 17380 12142 17382
rect 12198 17380 12204 17382
rect 11896 17371 12204 17380
rect 11060 17264 11112 17270
rect 11060 17206 11112 17212
rect 12912 17202 12940 19200
rect 14200 17202 14228 19200
rect 16132 19106 16160 19200
rect 16120 19100 16172 19106
rect 16120 19042 16172 19048
rect 16856 19100 16908 19106
rect 16856 19042 16908 19048
rect 16868 17202 16896 19042
rect 17420 17354 17448 19200
rect 17236 17326 17448 17354
rect 1308 17196 1360 17202
rect 1308 17138 1360 17144
rect 4528 17196 4580 17202
rect 4528 17138 4580 17144
rect 6460 17196 6512 17202
rect 6460 17138 6512 17144
rect 7748 17196 7800 17202
rect 7748 17138 7800 17144
rect 9680 17196 9732 17202
rect 9680 17138 9732 17144
rect 12900 17196 12952 17202
rect 12900 17138 12952 17144
rect 14188 17196 14240 17202
rect 14188 17138 14240 17144
rect 16856 17196 16908 17202
rect 16856 17138 16908 17144
rect 10876 17128 10928 17134
rect 10876 17070 10928 17076
rect 3608 17060 3660 17066
rect 3608 17002 3660 17008
rect 1768 16992 1820 16998
rect 1768 16934 1820 16940
rect 2504 16992 2556 16998
rect 2504 16934 2556 16940
rect 1032 16108 1084 16114
rect 1032 16050 1084 16056
rect 1030 15056 1086 15065
rect 1030 14991 1086 15000
rect 1044 13938 1072 14991
rect 1032 13932 1084 13938
rect 1032 13874 1084 13880
rect 940 13864 992 13870
rect 940 13806 992 13812
rect 952 13705 980 13806
rect 938 13696 994 13705
rect 938 13631 994 13640
rect 940 10464 992 10470
rect 940 10406 992 10412
rect 952 10305 980 10406
rect 938 10296 994 10305
rect 938 10231 994 10240
rect 1780 9489 1808 16934
rect 2134 12200 2190 12209
rect 2134 12135 2190 12144
rect 2148 11762 2176 12135
rect 2136 11756 2188 11762
rect 2136 11698 2188 11704
rect 2516 9654 2544 16934
rect 3056 13932 3108 13938
rect 3056 13874 3108 13880
rect 3068 12986 3096 13874
rect 3056 12980 3108 12986
rect 3056 12922 3108 12928
rect 3424 12844 3476 12850
rect 3424 12786 3476 12792
rect 3332 11756 3384 11762
rect 3332 11698 3384 11704
rect 2780 11688 2832 11694
rect 2780 11630 2832 11636
rect 2792 10470 2820 11630
rect 3344 11150 3372 11698
rect 3436 11354 3464 12786
rect 3424 11348 3476 11354
rect 3424 11290 3476 11296
rect 3436 11150 3464 11290
rect 3332 11144 3384 11150
rect 3332 11086 3384 11092
rect 3424 11144 3476 11150
rect 3424 11086 3476 11092
rect 2872 11076 2924 11082
rect 2872 11018 2924 11024
rect 2780 10464 2832 10470
rect 2780 10406 2832 10412
rect 2884 10266 2912 11018
rect 3344 10674 3372 11086
rect 3240 10668 3292 10674
rect 3240 10610 3292 10616
rect 3332 10668 3384 10674
rect 3332 10610 3384 10616
rect 3252 10266 3280 10610
rect 2872 10260 2924 10266
rect 2872 10202 2924 10208
rect 3240 10260 3292 10266
rect 3240 10202 3292 10208
rect 2504 9648 2556 9654
rect 2504 9590 2556 9596
rect 3148 9580 3200 9586
rect 3148 9522 3200 9528
rect 1766 9480 1822 9489
rect 1766 9415 1822 9424
rect 2780 9376 2832 9382
rect 2780 9318 2832 9324
rect 2792 8634 2820 9318
rect 2780 8628 2832 8634
rect 2780 8570 2832 8576
rect 938 8256 994 8265
rect 938 8191 994 8200
rect 952 7886 980 8191
rect 3160 7954 3188 9522
rect 3620 8537 3648 17002
rect 10232 16992 10284 16998
rect 10232 16934 10284 16940
rect 6423 16892 6731 16901
rect 6423 16890 6429 16892
rect 6485 16890 6509 16892
rect 6565 16890 6589 16892
rect 6645 16890 6669 16892
rect 6725 16890 6731 16892
rect 6485 16838 6487 16890
rect 6667 16838 6669 16890
rect 6423 16836 6429 16838
rect 6485 16836 6509 16838
rect 6565 16836 6589 16838
rect 6645 16836 6669 16838
rect 6725 16836 6731 16838
rect 6423 16827 6731 16836
rect 5172 16652 5224 16658
rect 5172 16594 5224 16600
rect 4712 14408 4764 14414
rect 4712 14350 4764 14356
rect 4344 14340 4396 14346
rect 4344 14282 4396 14288
rect 4160 14272 4212 14278
rect 4160 14214 4212 14220
rect 4172 13530 4200 14214
rect 4160 13524 4212 13530
rect 4160 13466 4212 13472
rect 4068 13320 4120 13326
rect 4068 13262 4120 13268
rect 4080 12306 4108 13262
rect 4356 13190 4384 14282
rect 4724 14074 4752 14350
rect 4712 14068 4764 14074
rect 4712 14010 4764 14016
rect 4988 13932 5040 13938
rect 4988 13874 5040 13880
rect 5000 13530 5028 13874
rect 4988 13524 5040 13530
rect 4988 13466 5040 13472
rect 4344 13184 4396 13190
rect 4344 13126 4396 13132
rect 4356 12850 4384 13126
rect 4528 12980 4580 12986
rect 4528 12922 4580 12928
rect 4344 12844 4396 12850
rect 4344 12786 4396 12792
rect 4436 12776 4488 12782
rect 4436 12718 4488 12724
rect 4068 12300 4120 12306
rect 4068 12242 4120 12248
rect 3884 12096 3936 12102
rect 3884 12038 3936 12044
rect 3896 11762 3924 12038
rect 4080 11898 4108 12242
rect 4344 12232 4396 12238
rect 4344 12174 4396 12180
rect 4068 11892 4120 11898
rect 4068 11834 4120 11840
rect 4356 11762 4384 12174
rect 3884 11756 3936 11762
rect 3884 11698 3936 11704
rect 4344 11756 4396 11762
rect 4344 11698 4396 11704
rect 4066 11656 4122 11665
rect 4122 11614 4200 11642
rect 4066 11591 4122 11600
rect 3884 11076 3936 11082
rect 3884 11018 3936 11024
rect 3896 9450 3924 11018
rect 3976 11008 4028 11014
rect 3976 10950 4028 10956
rect 3988 10062 4016 10950
rect 3976 10056 4028 10062
rect 3976 9998 4028 10004
rect 3884 9444 3936 9450
rect 3884 9386 3936 9392
rect 4172 8974 4200 11614
rect 4448 11354 4476 12718
rect 4540 12374 4568 12922
rect 4896 12912 4948 12918
rect 4896 12854 4948 12860
rect 4528 12368 4580 12374
rect 4528 12310 4580 12316
rect 4908 12238 4936 12854
rect 4896 12232 4948 12238
rect 4896 12174 4948 12180
rect 4988 12232 5040 12238
rect 4988 12174 5040 12180
rect 5000 11898 5028 12174
rect 4988 11892 5040 11898
rect 4988 11834 5040 11840
rect 4436 11348 4488 11354
rect 4436 11290 4488 11296
rect 4620 11212 4672 11218
rect 4620 11154 4672 11160
rect 4344 10532 4396 10538
rect 4344 10474 4396 10480
rect 4356 10062 4384 10474
rect 4632 10130 4660 11154
rect 5184 11150 5212 16594
rect 7012 16584 7064 16590
rect 7012 16526 7064 16532
rect 6423 15804 6731 15813
rect 6423 15802 6429 15804
rect 6485 15802 6509 15804
rect 6565 15802 6589 15804
rect 6645 15802 6669 15804
rect 6725 15802 6731 15804
rect 6485 15750 6487 15802
rect 6667 15750 6669 15802
rect 6423 15748 6429 15750
rect 6485 15748 6509 15750
rect 6565 15748 6589 15750
rect 6645 15748 6669 15750
rect 6725 15748 6731 15750
rect 6423 15739 6731 15748
rect 5632 15020 5684 15026
rect 5632 14962 5684 14968
rect 5644 14618 5672 14962
rect 6828 14816 6880 14822
rect 6828 14758 6880 14764
rect 6423 14716 6731 14725
rect 6423 14714 6429 14716
rect 6485 14714 6509 14716
rect 6565 14714 6589 14716
rect 6645 14714 6669 14716
rect 6725 14714 6731 14716
rect 6485 14662 6487 14714
rect 6667 14662 6669 14714
rect 6423 14660 6429 14662
rect 6485 14660 6509 14662
rect 6565 14660 6589 14662
rect 6645 14660 6669 14662
rect 6725 14660 6731 14662
rect 6423 14651 6731 14660
rect 5632 14612 5684 14618
rect 5632 14554 5684 14560
rect 5816 14612 5868 14618
rect 5816 14554 5868 14560
rect 5632 14408 5684 14414
rect 5632 14350 5684 14356
rect 5724 14408 5776 14414
rect 5724 14350 5776 14356
rect 5644 14074 5672 14350
rect 5632 14068 5684 14074
rect 5632 14010 5684 14016
rect 5540 14000 5592 14006
rect 5540 13942 5592 13948
rect 5264 13864 5316 13870
rect 5264 13806 5316 13812
rect 5276 12918 5304 13806
rect 5264 12912 5316 12918
rect 5264 12854 5316 12860
rect 5552 12238 5580 13942
rect 5736 13802 5764 14350
rect 5828 13938 5856 14554
rect 6552 14408 6604 14414
rect 6552 14350 6604 14356
rect 6564 13938 6592 14350
rect 6840 14006 6868 14758
rect 6828 14000 6880 14006
rect 6828 13942 6880 13948
rect 5816 13932 5868 13938
rect 5816 13874 5868 13880
rect 6552 13932 6604 13938
rect 6552 13874 6604 13880
rect 5724 13796 5776 13802
rect 5724 13738 5776 13744
rect 5828 13258 5856 13874
rect 6000 13728 6052 13734
rect 6000 13670 6052 13676
rect 6012 13258 6040 13670
rect 6423 13628 6731 13637
rect 6423 13626 6429 13628
rect 6485 13626 6509 13628
rect 6565 13626 6589 13628
rect 6645 13626 6669 13628
rect 6725 13626 6731 13628
rect 6485 13574 6487 13626
rect 6667 13574 6669 13626
rect 6423 13572 6429 13574
rect 6485 13572 6509 13574
rect 6565 13572 6589 13574
rect 6645 13572 6669 13574
rect 6725 13572 6731 13574
rect 6423 13563 6731 13572
rect 6828 13524 6880 13530
rect 6828 13466 6880 13472
rect 5816 13252 5868 13258
rect 5816 13194 5868 13200
rect 6000 13252 6052 13258
rect 6000 13194 6052 13200
rect 6552 13184 6604 13190
rect 6552 13126 6604 13132
rect 5724 12980 5776 12986
rect 5724 12922 5776 12928
rect 5736 12730 5764 12922
rect 6564 12850 6592 13126
rect 6840 12850 6868 13466
rect 6552 12844 6604 12850
rect 6552 12786 6604 12792
rect 6828 12844 6880 12850
rect 6828 12786 6880 12792
rect 5736 12702 5856 12730
rect 5828 12646 5856 12702
rect 5724 12640 5776 12646
rect 5724 12582 5776 12588
rect 5816 12640 5868 12646
rect 5816 12582 5868 12588
rect 6920 12640 6972 12646
rect 6920 12582 6972 12588
rect 5540 12232 5592 12238
rect 5540 12174 5592 12180
rect 5356 11348 5408 11354
rect 5356 11290 5408 11296
rect 5172 11144 5224 11150
rect 5172 11086 5224 11092
rect 5184 10742 5212 11086
rect 5172 10736 5224 10742
rect 5368 10713 5396 11290
rect 5552 11150 5580 12174
rect 5736 12170 5764 12582
rect 5724 12164 5776 12170
rect 5724 12106 5776 12112
rect 5828 11762 5856 12582
rect 6423 12540 6731 12549
rect 6423 12538 6429 12540
rect 6485 12538 6509 12540
rect 6565 12538 6589 12540
rect 6645 12538 6669 12540
rect 6725 12538 6731 12540
rect 6485 12486 6487 12538
rect 6667 12486 6669 12538
rect 6423 12484 6429 12486
rect 6485 12484 6509 12486
rect 6565 12484 6589 12486
rect 6645 12484 6669 12486
rect 6725 12484 6731 12486
rect 6423 12475 6731 12484
rect 6932 12442 6960 12582
rect 6920 12436 6972 12442
rect 6920 12378 6972 12384
rect 6932 12238 6960 12378
rect 6920 12232 6972 12238
rect 6920 12174 6972 12180
rect 5908 12164 5960 12170
rect 5908 12106 5960 12112
rect 5920 11830 5948 12106
rect 5908 11824 5960 11830
rect 5908 11766 5960 11772
rect 6918 11792 6974 11801
rect 5816 11756 5868 11762
rect 6918 11727 6920 11736
rect 5816 11698 5868 11704
rect 6972 11727 6974 11736
rect 6920 11698 6972 11704
rect 6423 11452 6731 11461
rect 6423 11450 6429 11452
rect 6485 11450 6509 11452
rect 6565 11450 6589 11452
rect 6645 11450 6669 11452
rect 6725 11450 6731 11452
rect 6485 11398 6487 11450
rect 6667 11398 6669 11450
rect 6423 11396 6429 11398
rect 6485 11396 6509 11398
rect 6565 11396 6589 11398
rect 6645 11396 6669 11398
rect 6725 11396 6731 11398
rect 6423 11387 6731 11396
rect 6932 11354 6960 11698
rect 6920 11348 6972 11354
rect 6920 11290 6972 11296
rect 5540 11144 5592 11150
rect 5540 11086 5592 11092
rect 5172 10678 5224 10684
rect 5354 10704 5410 10713
rect 4988 10668 5040 10674
rect 5354 10639 5356 10648
rect 4988 10610 5040 10616
rect 5408 10639 5410 10648
rect 5356 10610 5408 10616
rect 4620 10124 4672 10130
rect 4620 10066 4672 10072
rect 4344 10056 4396 10062
rect 4344 9998 4396 10004
rect 4436 9920 4488 9926
rect 4436 9862 4488 9868
rect 4160 8968 4212 8974
rect 4160 8910 4212 8916
rect 3792 8628 3844 8634
rect 3844 8588 4016 8616
rect 3792 8570 3844 8576
rect 3606 8528 3662 8537
rect 3988 8498 4016 8588
rect 4448 8566 4476 9862
rect 4436 8560 4488 8566
rect 4436 8502 4488 8508
rect 3606 8463 3662 8472
rect 3976 8492 4028 8498
rect 3976 8434 4028 8440
rect 3148 7948 3200 7954
rect 3148 7890 3200 7896
rect 940 7880 992 7886
rect 940 7822 992 7828
rect 2964 7744 3016 7750
rect 2964 7686 3016 7692
rect 938 6896 994 6905
rect 938 6831 994 6840
rect 952 5914 980 6831
rect 940 5908 992 5914
rect 940 5850 992 5856
rect 2976 5710 3004 7686
rect 3160 7002 3188 7890
rect 3988 7546 4016 8434
rect 3976 7540 4028 7546
rect 3976 7482 4028 7488
rect 3148 6996 3200 7002
rect 3148 6938 3200 6944
rect 3988 6914 4016 7482
rect 5000 7206 5028 10610
rect 5552 10470 5580 11086
rect 7024 10810 7052 16526
rect 10244 15502 10272 16934
rect 10888 16574 10916 17070
rect 15660 17060 15712 17066
rect 15660 17002 15712 17008
rect 10704 16546 10916 16574
rect 10140 15496 10192 15502
rect 10140 15438 10192 15444
rect 10232 15496 10284 15502
rect 10232 15438 10284 15444
rect 7380 15020 7432 15026
rect 7380 14962 7432 14968
rect 7196 14816 7248 14822
rect 7196 14758 7248 14764
rect 7208 14414 7236 14758
rect 7196 14408 7248 14414
rect 7196 14350 7248 14356
rect 7104 13932 7156 13938
rect 7104 13874 7156 13880
rect 7116 13258 7144 13874
rect 7392 13462 7420 14962
rect 7840 14612 7892 14618
rect 7840 14554 7892 14560
rect 7852 14074 7880 14554
rect 10152 14482 10180 15438
rect 10140 14476 10192 14482
rect 10140 14418 10192 14424
rect 8208 14272 8260 14278
rect 8208 14214 8260 14220
rect 8484 14272 8536 14278
rect 8484 14214 8536 14220
rect 7840 14068 7892 14074
rect 7840 14010 7892 14016
rect 8220 14006 8248 14214
rect 8208 14000 8260 14006
rect 8208 13942 8260 13948
rect 7380 13456 7432 13462
rect 7380 13398 7432 13404
rect 8220 13326 8248 13942
rect 8496 13938 8524 14214
rect 9772 14068 9824 14074
rect 9772 14010 9824 14016
rect 8484 13932 8536 13938
rect 8484 13874 8536 13880
rect 9404 13932 9456 13938
rect 9404 13874 9456 13880
rect 8208 13320 8260 13326
rect 8208 13262 8260 13268
rect 8496 13258 8524 13874
rect 8760 13728 8812 13734
rect 8760 13670 8812 13676
rect 8772 13530 8800 13670
rect 8760 13524 8812 13530
rect 8760 13466 8812 13472
rect 7104 13252 7156 13258
rect 7104 13194 7156 13200
rect 8484 13252 8536 13258
rect 8484 13194 8536 13200
rect 9416 12850 9444 13874
rect 9404 12844 9456 12850
rect 9404 12786 9456 12792
rect 9784 12238 9812 14010
rect 9864 12300 9916 12306
rect 9864 12242 9916 12248
rect 9772 12232 9824 12238
rect 9772 12174 9824 12180
rect 7748 12096 7800 12102
rect 7748 12038 7800 12044
rect 7760 11762 7788 12038
rect 7656 11756 7708 11762
rect 7656 11698 7708 11704
rect 7748 11756 7800 11762
rect 7748 11698 7800 11704
rect 7104 11688 7156 11694
rect 7104 11630 7156 11636
rect 7012 10804 7064 10810
rect 7012 10746 7064 10752
rect 5540 10464 5592 10470
rect 5540 10406 5592 10412
rect 6423 10364 6731 10373
rect 6423 10362 6429 10364
rect 6485 10362 6509 10364
rect 6565 10362 6589 10364
rect 6645 10362 6669 10364
rect 6725 10362 6731 10364
rect 6485 10310 6487 10362
rect 6667 10310 6669 10362
rect 6423 10308 6429 10310
rect 6485 10308 6509 10310
rect 6565 10308 6589 10310
rect 6645 10308 6669 10310
rect 6725 10308 6731 10310
rect 6423 10299 6731 10308
rect 5816 10124 5868 10130
rect 5816 10066 5868 10072
rect 5632 9580 5684 9586
rect 5632 9522 5684 9528
rect 5644 8974 5672 9522
rect 5828 9518 5856 10066
rect 6276 10056 6328 10062
rect 6276 9998 6328 10004
rect 6288 9518 6316 9998
rect 5816 9512 5868 9518
rect 5816 9454 5868 9460
rect 6276 9512 6328 9518
rect 6276 9454 6328 9460
rect 5828 9178 5856 9454
rect 6184 9376 6236 9382
rect 6184 9318 6236 9324
rect 5816 9172 5868 9178
rect 5816 9114 5868 9120
rect 5632 8968 5684 8974
rect 5632 8910 5684 8916
rect 5540 8832 5592 8838
rect 5540 8774 5592 8780
rect 5356 8288 5408 8294
rect 5356 8230 5408 8236
rect 5264 7744 5316 7750
rect 5264 7686 5316 7692
rect 5172 7404 5224 7410
rect 5172 7346 5224 7352
rect 5080 7336 5132 7342
rect 5080 7278 5132 7284
rect 4252 7200 4304 7206
rect 4252 7142 4304 7148
rect 4988 7200 5040 7206
rect 4988 7142 5040 7148
rect 3896 6886 4016 6914
rect 3896 6798 3924 6886
rect 3884 6792 3936 6798
rect 3884 6734 3936 6740
rect 4264 6390 4292 7142
rect 4436 6724 4488 6730
rect 4436 6666 4488 6672
rect 4344 6452 4396 6458
rect 4344 6394 4396 6400
rect 4252 6384 4304 6390
rect 4252 6326 4304 6332
rect 3976 6248 4028 6254
rect 3976 6190 4028 6196
rect 3988 5710 4016 6190
rect 2964 5704 3016 5710
rect 2964 5646 3016 5652
rect 3976 5704 4028 5710
rect 3976 5646 4028 5652
rect 4356 5370 4384 6394
rect 4448 5370 4476 6666
rect 4528 6316 4580 6322
rect 4528 6258 4580 6264
rect 4344 5364 4396 5370
rect 4344 5306 4396 5312
rect 4436 5364 4488 5370
rect 4436 5306 4488 5312
rect 940 5160 992 5166
rect 940 5102 992 5108
rect 1860 5160 1912 5166
rect 1860 5102 1912 5108
rect 952 4865 980 5102
rect 938 4856 994 4865
rect 938 4791 994 4800
rect 1872 4758 1900 5102
rect 1860 4752 1912 4758
rect 1860 4694 1912 4700
rect 4356 4690 4384 5306
rect 4540 5098 4568 6258
rect 4712 5704 4764 5710
rect 4712 5646 4764 5652
rect 4724 5234 4752 5646
rect 4712 5228 4764 5234
rect 4712 5170 4764 5176
rect 4528 5092 4580 5098
rect 4528 5034 4580 5040
rect 4344 4684 4396 4690
rect 4344 4626 4396 4632
rect 4724 4622 4752 5170
rect 5092 5166 5120 7278
rect 5184 6458 5212 7346
rect 5172 6452 5224 6458
rect 5172 6394 5224 6400
rect 5276 5914 5304 7686
rect 5368 7546 5396 8230
rect 5552 7886 5580 8774
rect 5828 7886 5856 9114
rect 5540 7880 5592 7886
rect 5540 7822 5592 7828
rect 5816 7880 5868 7886
rect 5816 7822 5868 7828
rect 5448 7812 5500 7818
rect 5448 7754 5500 7760
rect 5356 7540 5408 7546
rect 5356 7482 5408 7488
rect 5368 6798 5396 7482
rect 5460 7342 5488 7754
rect 5552 7478 5580 7822
rect 5540 7472 5592 7478
rect 5540 7414 5592 7420
rect 5448 7336 5500 7342
rect 5448 7278 5500 7284
rect 5448 7200 5500 7206
rect 5448 7142 5500 7148
rect 5356 6792 5408 6798
rect 5356 6734 5408 6740
rect 5264 5908 5316 5914
rect 5264 5850 5316 5856
rect 5276 5234 5304 5850
rect 5460 5710 5488 7142
rect 6196 6798 6224 9318
rect 6288 8906 6316 9454
rect 6423 9276 6731 9285
rect 6423 9274 6429 9276
rect 6485 9274 6509 9276
rect 6565 9274 6589 9276
rect 6645 9274 6669 9276
rect 6725 9274 6731 9276
rect 6485 9222 6487 9274
rect 6667 9222 6669 9274
rect 6423 9220 6429 9222
rect 6485 9220 6509 9222
rect 6565 9220 6589 9222
rect 6645 9220 6669 9222
rect 6725 9220 6731 9222
rect 6423 9211 6731 9220
rect 7116 9178 7144 11630
rect 7668 9450 7696 11698
rect 7932 11552 7984 11558
rect 7932 11494 7984 11500
rect 7944 11150 7972 11494
rect 9876 11354 9904 12242
rect 9864 11348 9916 11354
rect 9864 11290 9916 11296
rect 7932 11144 7984 11150
rect 7932 11086 7984 11092
rect 9956 11144 10008 11150
rect 9956 11086 10008 11092
rect 9968 10810 9996 11086
rect 9956 10804 10008 10810
rect 9956 10746 10008 10752
rect 10152 10470 10180 14418
rect 10704 11642 10732 16546
rect 11896 16348 12204 16357
rect 11896 16346 11902 16348
rect 11958 16346 11982 16348
rect 12038 16346 12062 16348
rect 12118 16346 12142 16348
rect 12198 16346 12204 16348
rect 11958 16294 11960 16346
rect 12140 16294 12142 16346
rect 11896 16292 11902 16294
rect 11958 16292 11982 16294
rect 12038 16292 12062 16294
rect 12118 16292 12142 16294
rect 12198 16292 12204 16294
rect 11896 16283 12204 16292
rect 12624 15360 12676 15366
rect 12624 15302 12676 15308
rect 11896 15260 12204 15269
rect 11896 15258 11902 15260
rect 11958 15258 11982 15260
rect 12038 15258 12062 15260
rect 12118 15258 12142 15260
rect 12198 15258 12204 15260
rect 11958 15206 11960 15258
rect 12140 15206 12142 15258
rect 11896 15204 11902 15206
rect 11958 15204 11982 15206
rect 12038 15204 12062 15206
rect 12118 15204 12142 15206
rect 12198 15204 12204 15206
rect 11896 15195 12204 15204
rect 12636 15026 12664 15302
rect 12624 15020 12676 15026
rect 12624 14962 12676 14968
rect 13820 15020 13872 15026
rect 13820 14962 13872 14968
rect 15200 15020 15252 15026
rect 15200 14962 15252 14968
rect 12256 14408 12308 14414
rect 12256 14350 12308 14356
rect 11336 14272 11388 14278
rect 11336 14214 11388 14220
rect 11244 14000 11296 14006
rect 11244 13942 11296 13948
rect 11152 13932 11204 13938
rect 11152 13874 11204 13880
rect 11060 13524 11112 13530
rect 11060 13466 11112 13472
rect 11072 12986 11100 13466
rect 11164 13394 11192 13874
rect 11256 13462 11284 13942
rect 11348 13870 11376 14214
rect 11896 14172 12204 14181
rect 11896 14170 11902 14172
rect 11958 14170 11982 14172
rect 12038 14170 12062 14172
rect 12118 14170 12142 14172
rect 12198 14170 12204 14172
rect 11958 14118 11960 14170
rect 12140 14118 12142 14170
rect 11896 14116 11902 14118
rect 11958 14116 11982 14118
rect 12038 14116 12062 14118
rect 12118 14116 12142 14118
rect 12198 14116 12204 14118
rect 11896 14107 12204 14116
rect 12268 14074 12296 14350
rect 12348 14272 12400 14278
rect 12348 14214 12400 14220
rect 13544 14272 13596 14278
rect 13544 14214 13596 14220
rect 12256 14068 12308 14074
rect 12256 14010 12308 14016
rect 11336 13864 11388 13870
rect 11336 13806 11388 13812
rect 11244 13456 11296 13462
rect 11244 13398 11296 13404
rect 11152 13388 11204 13394
rect 11152 13330 11204 13336
rect 11348 13326 11376 13806
rect 12360 13462 12388 14214
rect 12624 13864 12676 13870
rect 12624 13806 12676 13812
rect 12636 13530 12664 13806
rect 12716 13728 12768 13734
rect 12716 13670 12768 13676
rect 12624 13524 12676 13530
rect 12624 13466 12676 13472
rect 12348 13456 12400 13462
rect 12348 13398 12400 13404
rect 11520 13388 11572 13394
rect 11520 13330 11572 13336
rect 11336 13320 11388 13326
rect 11336 13262 11388 13268
rect 11060 12980 11112 12986
rect 11060 12922 11112 12928
rect 11336 12912 11388 12918
rect 11336 12854 11388 12860
rect 11060 12844 11112 12850
rect 11060 12786 11112 12792
rect 11152 12844 11204 12850
rect 11152 12786 11204 12792
rect 11244 12844 11296 12850
rect 11244 12786 11296 12792
rect 10784 12708 10836 12714
rect 10784 12650 10836 12656
rect 10796 12306 10824 12650
rect 10784 12300 10836 12306
rect 10784 12242 10836 12248
rect 10968 12300 11020 12306
rect 10968 12242 11020 12248
rect 10980 12186 11008 12242
rect 10888 12158 11008 12186
rect 10888 11762 10916 12158
rect 11072 12102 11100 12786
rect 11164 12170 11192 12786
rect 11152 12164 11204 12170
rect 11152 12106 11204 12112
rect 11060 12096 11112 12102
rect 11060 12038 11112 12044
rect 11256 11898 11284 12786
rect 11348 12238 11376 12854
rect 11532 12442 11560 13330
rect 12532 13252 12584 13258
rect 12532 13194 12584 13200
rect 11896 13084 12204 13093
rect 11896 13082 11902 13084
rect 11958 13082 11982 13084
rect 12038 13082 12062 13084
rect 12118 13082 12142 13084
rect 12198 13082 12204 13084
rect 11958 13030 11960 13082
rect 12140 13030 12142 13082
rect 11896 13028 11902 13030
rect 11958 13028 11982 13030
rect 12038 13028 12062 13030
rect 12118 13028 12142 13030
rect 12198 13028 12204 13030
rect 11896 13019 12204 13028
rect 12440 12912 12492 12918
rect 12440 12854 12492 12860
rect 12348 12844 12400 12850
rect 12348 12786 12400 12792
rect 11520 12436 11572 12442
rect 11520 12378 11572 12384
rect 11336 12232 11388 12238
rect 11336 12174 11388 12180
rect 11428 12232 11480 12238
rect 11428 12174 11480 12180
rect 11244 11892 11296 11898
rect 11244 11834 11296 11840
rect 10876 11756 10928 11762
rect 10876 11698 10928 11704
rect 10704 11614 10916 11642
rect 10692 11008 10744 11014
rect 10692 10950 10744 10956
rect 10140 10464 10192 10470
rect 10140 10406 10192 10412
rect 10324 10464 10376 10470
rect 10324 10406 10376 10412
rect 10336 10130 10364 10406
rect 10704 10130 10732 10950
rect 10888 10606 10916 11614
rect 11244 11552 11296 11558
rect 11244 11494 11296 11500
rect 11256 11218 11284 11494
rect 11244 11212 11296 11218
rect 11244 11154 11296 11160
rect 11152 11008 11204 11014
rect 11152 10950 11204 10956
rect 11164 10674 11192 10950
rect 11256 10810 11284 11154
rect 11348 10810 11376 12174
rect 11440 11762 11468 12174
rect 11520 12164 11572 12170
rect 11520 12106 11572 12112
rect 12256 12164 12308 12170
rect 12256 12106 12308 12112
rect 11428 11756 11480 11762
rect 11428 11698 11480 11704
rect 11244 10804 11296 10810
rect 11244 10746 11296 10752
rect 11336 10804 11388 10810
rect 11336 10746 11388 10752
rect 11152 10668 11204 10674
rect 11152 10610 11204 10616
rect 10876 10600 10928 10606
rect 10876 10542 10928 10548
rect 10968 10600 11020 10606
rect 10968 10542 11020 10548
rect 10888 10470 10916 10542
rect 10876 10464 10928 10470
rect 10876 10406 10928 10412
rect 10324 10124 10376 10130
rect 10324 10066 10376 10072
rect 10692 10124 10744 10130
rect 10692 10066 10744 10072
rect 7932 9920 7984 9926
rect 7932 9862 7984 9868
rect 7944 9654 7972 9862
rect 7932 9648 7984 9654
rect 7932 9590 7984 9596
rect 10692 9580 10744 9586
rect 10692 9522 10744 9528
rect 7656 9444 7708 9450
rect 7656 9386 7708 9392
rect 7104 9172 7156 9178
rect 7104 9114 7156 9120
rect 7564 9104 7616 9110
rect 7564 9046 7616 9052
rect 6276 8900 6328 8906
rect 6276 8842 6328 8848
rect 6288 8430 6316 8842
rect 7012 8560 7064 8566
rect 6840 8508 7012 8514
rect 6840 8502 7064 8508
rect 6840 8486 7052 8502
rect 6276 8424 6328 8430
rect 6276 8366 6328 8372
rect 6288 8090 6316 8366
rect 6423 8188 6731 8197
rect 6423 8186 6429 8188
rect 6485 8186 6509 8188
rect 6565 8186 6589 8188
rect 6645 8186 6669 8188
rect 6725 8186 6731 8188
rect 6485 8134 6487 8186
rect 6667 8134 6669 8186
rect 6423 8132 6429 8134
rect 6485 8132 6509 8134
rect 6565 8132 6589 8134
rect 6645 8132 6669 8134
rect 6725 8132 6731 8134
rect 6423 8123 6731 8132
rect 6276 8084 6328 8090
rect 6276 8026 6328 8032
rect 6423 7100 6731 7109
rect 6423 7098 6429 7100
rect 6485 7098 6509 7100
rect 6565 7098 6589 7100
rect 6645 7098 6669 7100
rect 6725 7098 6731 7100
rect 6485 7046 6487 7098
rect 6667 7046 6669 7098
rect 6423 7044 6429 7046
rect 6485 7044 6509 7046
rect 6565 7044 6589 7046
rect 6645 7044 6669 7046
rect 6725 7044 6731 7046
rect 6423 7035 6731 7044
rect 6184 6792 6236 6798
rect 6184 6734 6236 6740
rect 6840 6662 6868 8486
rect 7288 7744 7340 7750
rect 7288 7686 7340 7692
rect 6920 7472 6972 7478
rect 6920 7414 6972 7420
rect 6932 6866 6960 7414
rect 7300 7410 7328 7686
rect 7288 7404 7340 7410
rect 7288 7346 7340 7352
rect 6920 6860 6972 6866
rect 6920 6802 6972 6808
rect 6828 6656 6880 6662
rect 6828 6598 6880 6604
rect 6000 6452 6052 6458
rect 6000 6394 6052 6400
rect 6012 5710 6040 6394
rect 6423 6012 6731 6021
rect 6423 6010 6429 6012
rect 6485 6010 6509 6012
rect 6565 6010 6589 6012
rect 6645 6010 6669 6012
rect 6725 6010 6731 6012
rect 6485 5958 6487 6010
rect 6667 5958 6669 6010
rect 6423 5956 6429 5958
rect 6485 5956 6509 5958
rect 6565 5956 6589 5958
rect 6645 5956 6669 5958
rect 6725 5956 6731 5958
rect 6423 5947 6731 5956
rect 5448 5704 5500 5710
rect 5448 5646 5500 5652
rect 6000 5704 6052 5710
rect 6000 5646 6052 5652
rect 6932 5642 6960 6802
rect 7576 6798 7604 9046
rect 7668 8634 7696 9386
rect 10704 9042 10732 9522
rect 10980 9518 11008 10542
rect 11256 10266 11284 10746
rect 11244 10260 11296 10266
rect 11244 10202 11296 10208
rect 11532 10198 11560 12106
rect 11796 12096 11848 12102
rect 11796 12038 11848 12044
rect 11808 11762 11836 12038
rect 11896 11996 12204 12005
rect 11896 11994 11902 11996
rect 11958 11994 11982 11996
rect 12038 11994 12062 11996
rect 12118 11994 12142 11996
rect 12198 11994 12204 11996
rect 11958 11942 11960 11994
rect 12140 11942 12142 11994
rect 11896 11940 11902 11942
rect 11958 11940 11982 11942
rect 12038 11940 12062 11942
rect 12118 11940 12142 11942
rect 12198 11940 12204 11942
rect 11896 11931 12204 11940
rect 11796 11756 11848 11762
rect 11796 11698 11848 11704
rect 12072 11756 12124 11762
rect 12072 11698 12124 11704
rect 12084 11354 12112 11698
rect 12268 11642 12296 12106
rect 12360 11762 12388 12786
rect 12452 11762 12480 12854
rect 12544 12442 12572 13194
rect 12532 12436 12584 12442
rect 12532 12378 12584 12384
rect 12636 12238 12664 13466
rect 12728 13326 12756 13670
rect 12716 13320 12768 13326
rect 12716 13262 12768 13268
rect 12808 13320 12860 13326
rect 12808 13262 12860 13268
rect 12820 12986 12848 13262
rect 13084 13252 13136 13258
rect 13084 13194 13136 13200
rect 12992 13184 13044 13190
rect 12992 13126 13044 13132
rect 12808 12980 12860 12986
rect 12808 12922 12860 12928
rect 13004 12442 13032 13126
rect 13096 12850 13124 13194
rect 13084 12844 13136 12850
rect 13084 12786 13136 12792
rect 12992 12436 13044 12442
rect 12992 12378 13044 12384
rect 13360 12436 13412 12442
rect 13556 12434 13584 14214
rect 13636 13932 13688 13938
rect 13832 13920 13860 14962
rect 14280 14408 14332 14414
rect 14280 14350 14332 14356
rect 14464 14408 14516 14414
rect 14464 14350 14516 14356
rect 14292 14074 14320 14350
rect 14280 14068 14332 14074
rect 14280 14010 14332 14016
rect 13688 13892 13860 13920
rect 13636 13874 13688 13880
rect 13728 12912 13780 12918
rect 13832 12866 13860 13892
rect 14292 13326 14320 14010
rect 14476 13326 14504 14350
rect 15108 13932 15160 13938
rect 15108 13874 15160 13880
rect 14280 13320 14332 13326
rect 14280 13262 14332 13268
rect 14464 13320 14516 13326
rect 14464 13262 14516 13268
rect 13780 12860 13860 12866
rect 13728 12854 13860 12860
rect 13740 12838 13860 12854
rect 14292 12850 14320 13262
rect 14476 12986 14504 13262
rect 15120 13258 15148 13874
rect 15108 13252 15160 13258
rect 15108 13194 15160 13200
rect 14464 12980 14516 12986
rect 14464 12922 14516 12928
rect 13556 12406 13676 12434
rect 13360 12378 13412 12384
rect 12624 12232 12676 12238
rect 12624 12174 12676 12180
rect 12716 12232 12768 12238
rect 12716 12174 12768 12180
rect 12728 11898 12756 12174
rect 13372 12102 13400 12378
rect 13452 12300 13504 12306
rect 13452 12242 13504 12248
rect 13360 12096 13412 12102
rect 13360 12038 13412 12044
rect 12716 11892 12768 11898
rect 12716 11834 12768 11840
rect 12348 11756 12400 11762
rect 12348 11698 12400 11704
rect 12440 11756 12492 11762
rect 12440 11698 12492 11704
rect 12268 11614 12388 11642
rect 12072 11348 12124 11354
rect 12072 11290 12124 11296
rect 12256 11008 12308 11014
rect 12256 10950 12308 10956
rect 11896 10908 12204 10917
rect 11896 10906 11902 10908
rect 11958 10906 11982 10908
rect 12038 10906 12062 10908
rect 12118 10906 12142 10908
rect 12198 10906 12204 10908
rect 11958 10854 11960 10906
rect 12140 10854 12142 10906
rect 11896 10852 11902 10854
rect 11958 10852 11982 10854
rect 12038 10852 12062 10854
rect 12118 10852 12142 10854
rect 12198 10852 12204 10854
rect 11896 10843 12204 10852
rect 12268 10810 12296 10950
rect 12256 10804 12308 10810
rect 12256 10746 12308 10752
rect 11520 10192 11572 10198
rect 11520 10134 11572 10140
rect 11896 9820 12204 9829
rect 11896 9818 11902 9820
rect 11958 9818 11982 9820
rect 12038 9818 12062 9820
rect 12118 9818 12142 9820
rect 12198 9818 12204 9820
rect 11958 9766 11960 9818
rect 12140 9766 12142 9818
rect 11896 9764 11902 9766
rect 11958 9764 11982 9766
rect 12038 9764 12062 9766
rect 12118 9764 12142 9766
rect 12198 9764 12204 9766
rect 11896 9755 12204 9764
rect 12268 9654 12296 10746
rect 12360 9926 12388 11614
rect 13464 11354 13492 12242
rect 13648 12238 13676 12406
rect 13636 12232 13688 12238
rect 13636 12174 13688 12180
rect 13452 11348 13504 11354
rect 13452 11290 13504 11296
rect 12440 11212 12492 11218
rect 12440 11154 12492 11160
rect 12452 10606 12480 11154
rect 13648 11150 13676 12174
rect 13728 11688 13780 11694
rect 13728 11630 13780 11636
rect 13740 11286 13768 11630
rect 13728 11280 13780 11286
rect 13728 11222 13780 11228
rect 13636 11144 13688 11150
rect 13636 11086 13688 11092
rect 13176 11076 13228 11082
rect 13176 11018 13228 11024
rect 12900 10668 12952 10674
rect 12900 10610 12952 10616
rect 12440 10600 12492 10606
rect 12440 10542 12492 10548
rect 12452 10062 12480 10542
rect 12440 10056 12492 10062
rect 12440 9998 12492 10004
rect 12348 9920 12400 9926
rect 12348 9862 12400 9868
rect 12256 9648 12308 9654
rect 12256 9590 12308 9596
rect 10876 9512 10928 9518
rect 10876 9454 10928 9460
rect 10968 9512 11020 9518
rect 10968 9454 11020 9460
rect 10888 9178 10916 9454
rect 10876 9172 10928 9178
rect 10876 9114 10928 9120
rect 10980 9058 11008 9454
rect 11152 9376 11204 9382
rect 11152 9318 11204 9324
rect 10692 9036 10744 9042
rect 10692 8978 10744 8984
rect 10888 9030 11008 9058
rect 9956 8968 10008 8974
rect 9956 8910 10008 8916
rect 8024 8832 8076 8838
rect 8024 8774 8076 8780
rect 9772 8832 9824 8838
rect 9772 8774 9824 8780
rect 8036 8634 8064 8774
rect 7656 8628 7708 8634
rect 7656 8570 7708 8576
rect 8024 8628 8076 8634
rect 8024 8570 8076 8576
rect 8208 8492 8260 8498
rect 8208 8434 8260 8440
rect 7932 8356 7984 8362
rect 7932 8298 7984 8304
rect 7748 8288 7800 8294
rect 7748 8230 7800 8236
rect 7760 7410 7788 8230
rect 7944 7954 7972 8298
rect 8220 8022 8248 8434
rect 8208 8016 8260 8022
rect 8208 7958 8260 7964
rect 7932 7948 7984 7954
rect 7932 7890 7984 7896
rect 9784 7818 9812 8774
rect 9864 7880 9916 7886
rect 9864 7822 9916 7828
rect 9128 7812 9180 7818
rect 9128 7754 9180 7760
rect 9772 7812 9824 7818
rect 9772 7754 9824 7760
rect 9140 7546 9168 7754
rect 9128 7540 9180 7546
rect 9128 7482 9180 7488
rect 7748 7404 7800 7410
rect 7748 7346 7800 7352
rect 9140 6914 9168 7482
rect 9876 7410 9904 7822
rect 9864 7404 9916 7410
rect 9864 7346 9916 7352
rect 9048 6886 9168 6914
rect 7564 6792 7616 6798
rect 7564 6734 7616 6740
rect 9048 6322 9076 6886
rect 9404 6860 9456 6866
rect 9404 6802 9456 6808
rect 8484 6316 8536 6322
rect 8484 6258 8536 6264
rect 9036 6316 9088 6322
rect 9036 6258 9088 6264
rect 8300 6112 8352 6118
rect 8300 6054 8352 6060
rect 6920 5636 6972 5642
rect 6920 5578 6972 5584
rect 6184 5568 6236 5574
rect 6184 5510 6236 5516
rect 7196 5568 7248 5574
rect 7196 5510 7248 5516
rect 6196 5273 6224 5510
rect 7208 5302 7236 5510
rect 7196 5296 7248 5302
rect 6182 5264 6238 5273
rect 5264 5228 5316 5234
rect 7196 5238 7248 5244
rect 8312 5234 8340 6054
rect 8390 5808 8446 5817
rect 8390 5743 8446 5752
rect 8404 5710 8432 5743
rect 8392 5704 8444 5710
rect 8392 5646 8444 5652
rect 6182 5199 6238 5208
rect 8300 5228 8352 5234
rect 5264 5170 5316 5176
rect 8300 5170 8352 5176
rect 5080 5160 5132 5166
rect 5080 5102 5132 5108
rect 7196 5024 7248 5030
rect 7196 4966 7248 4972
rect 6423 4924 6731 4933
rect 6423 4922 6429 4924
rect 6485 4922 6509 4924
rect 6565 4922 6589 4924
rect 6645 4922 6669 4924
rect 6725 4922 6731 4924
rect 6485 4870 6487 4922
rect 6667 4870 6669 4922
rect 6423 4868 6429 4870
rect 6485 4868 6509 4870
rect 6565 4868 6589 4870
rect 6645 4868 6669 4870
rect 6725 4868 6731 4870
rect 6423 4859 6731 4868
rect 4712 4616 4764 4622
rect 4712 4558 4764 4564
rect 5632 4480 5684 4486
rect 5632 4422 5684 4428
rect 5644 3534 5672 4422
rect 6423 3836 6731 3845
rect 6423 3834 6429 3836
rect 6485 3834 6509 3836
rect 6565 3834 6589 3836
rect 6645 3834 6669 3836
rect 6725 3834 6731 3836
rect 6485 3782 6487 3834
rect 6667 3782 6669 3834
rect 6423 3780 6429 3782
rect 6485 3780 6509 3782
rect 6565 3780 6589 3782
rect 6645 3780 6669 3782
rect 6725 3780 6731 3782
rect 6423 3771 6731 3780
rect 6276 3596 6328 3602
rect 6276 3538 6328 3544
rect 940 3528 992 3534
rect 938 3496 940 3505
rect 5632 3528 5684 3534
rect 992 3496 994 3505
rect 5632 3470 5684 3476
rect 938 3431 994 3440
rect 940 2848 992 2854
rect 940 2790 992 2796
rect 20 2508 72 2514
rect 20 2450 72 2456
rect 32 800 60 2450
rect 952 1465 980 2790
rect 1308 2440 1360 2446
rect 1308 2382 1360 2388
rect 4160 2440 4212 2446
rect 4160 2382 4212 2388
rect 4528 2440 4580 2446
rect 4528 2382 4580 2388
rect 938 1456 994 1465
rect 938 1391 994 1400
rect 1320 800 1348 2382
rect 4172 950 4200 2382
rect 3240 944 3292 950
rect 3240 886 3292 892
rect 4160 944 4212 950
rect 4160 886 4212 892
rect 3252 800 3280 886
rect 4540 800 4568 2382
rect 6288 1714 6316 3538
rect 7208 3058 7236 4966
rect 8496 4010 8524 6258
rect 8944 6248 8996 6254
rect 8944 6190 8996 6196
rect 8956 5846 8984 6190
rect 9312 6112 9364 6118
rect 9312 6054 9364 6060
rect 8944 5840 8996 5846
rect 8944 5782 8996 5788
rect 8484 4004 8536 4010
rect 8484 3946 8536 3952
rect 9324 3194 9352 6054
rect 9416 5302 9444 6802
rect 9404 5296 9456 5302
rect 9404 5238 9456 5244
rect 9876 4622 9904 7346
rect 9968 6458 9996 8910
rect 10232 8900 10284 8906
rect 10232 8842 10284 8848
rect 10600 8900 10652 8906
rect 10600 8842 10652 8848
rect 10244 8566 10272 8842
rect 10324 8832 10376 8838
rect 10324 8774 10376 8780
rect 10336 8634 10364 8774
rect 10324 8628 10376 8634
rect 10324 8570 10376 8576
rect 10232 8560 10284 8566
rect 10232 8502 10284 8508
rect 10508 8492 10560 8498
rect 10508 8434 10560 8440
rect 10520 8090 10548 8434
rect 10612 8430 10640 8842
rect 10600 8424 10652 8430
rect 10600 8366 10652 8372
rect 10508 8084 10560 8090
rect 10508 8026 10560 8032
rect 10612 7886 10640 8366
rect 10888 8090 10916 9030
rect 10968 8900 11020 8906
rect 10968 8842 11020 8848
rect 10980 8634 11008 8842
rect 10968 8628 11020 8634
rect 10968 8570 11020 8576
rect 11164 8498 11192 9318
rect 12268 9178 12296 9590
rect 12256 9172 12308 9178
rect 12256 9114 12308 9120
rect 11896 8732 12204 8741
rect 11896 8730 11902 8732
rect 11958 8730 11982 8732
rect 12038 8730 12062 8732
rect 12118 8730 12142 8732
rect 12198 8730 12204 8732
rect 11958 8678 11960 8730
rect 12140 8678 12142 8730
rect 11896 8676 11902 8678
rect 11958 8676 11982 8678
rect 12038 8676 12062 8678
rect 12118 8676 12142 8678
rect 12198 8676 12204 8678
rect 11896 8667 12204 8676
rect 12912 8634 12940 10610
rect 13188 10062 13216 11018
rect 13832 10810 13860 12838
rect 14280 12844 14332 12850
rect 14280 12786 14332 12792
rect 14832 12640 14884 12646
rect 14832 12582 14884 12588
rect 14844 12374 14872 12582
rect 15120 12442 15148 13194
rect 15108 12436 15160 12442
rect 15108 12378 15160 12384
rect 14832 12368 14884 12374
rect 14832 12310 14884 12316
rect 14464 12096 14516 12102
rect 14464 12038 14516 12044
rect 14476 11898 14504 12038
rect 14464 11892 14516 11898
rect 14464 11834 14516 11840
rect 14476 11218 14504 11834
rect 14464 11212 14516 11218
rect 14464 11154 14516 11160
rect 13820 10804 13872 10810
rect 13820 10746 13872 10752
rect 13268 10668 13320 10674
rect 13268 10610 13320 10616
rect 13176 10056 13228 10062
rect 13176 9998 13228 10004
rect 13280 9654 13308 10610
rect 15212 10470 15240 14962
rect 15672 14414 15700 17002
rect 16580 16992 16632 16998
rect 16580 16934 16632 16940
rect 15660 14408 15712 14414
rect 15660 14350 15712 14356
rect 15292 14340 15344 14346
rect 15292 14282 15344 14288
rect 15476 14340 15528 14346
rect 15476 14282 15528 14288
rect 15304 13258 15332 14282
rect 15292 13252 15344 13258
rect 15292 13194 15344 13200
rect 15384 11144 15436 11150
rect 15384 11086 15436 11092
rect 15200 10464 15252 10470
rect 15200 10406 15252 10412
rect 14280 10260 14332 10266
rect 14280 10202 14332 10208
rect 14292 10062 14320 10202
rect 14832 10192 14884 10198
rect 14832 10134 14884 10140
rect 13452 10056 13504 10062
rect 13452 9998 13504 10004
rect 14280 10056 14332 10062
rect 14280 9998 14332 10004
rect 13464 9722 13492 9998
rect 14844 9926 14872 10134
rect 14832 9920 14884 9926
rect 14832 9862 14884 9868
rect 13452 9716 13504 9722
rect 13452 9658 13504 9664
rect 13544 9716 13596 9722
rect 13544 9658 13596 9664
rect 13268 9648 13320 9654
rect 13268 9590 13320 9596
rect 13084 9580 13136 9586
rect 13084 9522 13136 9528
rect 12992 9444 13044 9450
rect 12992 9386 13044 9392
rect 13004 9178 13032 9386
rect 13096 9178 13124 9522
rect 12992 9172 13044 9178
rect 12992 9114 13044 9120
rect 13084 9172 13136 9178
rect 13084 9114 13136 9120
rect 11612 8628 11664 8634
rect 11612 8570 11664 8576
rect 12900 8628 12952 8634
rect 12900 8570 12952 8576
rect 11520 8560 11572 8566
rect 11520 8502 11572 8508
rect 11152 8492 11204 8498
rect 11152 8434 11204 8440
rect 11532 8294 11560 8502
rect 11520 8288 11572 8294
rect 11520 8230 11572 8236
rect 10876 8084 10928 8090
rect 10876 8026 10928 8032
rect 10600 7880 10652 7886
rect 10600 7822 10652 7828
rect 10612 7002 10640 7822
rect 10968 7200 11020 7206
rect 10968 7142 11020 7148
rect 11060 7200 11112 7206
rect 11060 7142 11112 7148
rect 10140 6996 10192 7002
rect 10140 6938 10192 6944
rect 10600 6996 10652 7002
rect 10600 6938 10652 6944
rect 9956 6452 10008 6458
rect 9956 6394 10008 6400
rect 10152 6186 10180 6938
rect 10612 6866 10640 6938
rect 10600 6860 10652 6866
rect 10600 6802 10652 6808
rect 10692 6724 10744 6730
rect 10692 6666 10744 6672
rect 10704 6458 10732 6666
rect 10876 6656 10928 6662
rect 10876 6598 10928 6604
rect 10692 6452 10744 6458
rect 10692 6394 10744 6400
rect 10888 6390 10916 6598
rect 10876 6384 10928 6390
rect 10876 6326 10928 6332
rect 10980 6322 11008 7142
rect 11072 6798 11100 7142
rect 11060 6792 11112 6798
rect 11060 6734 11112 6740
rect 11624 6662 11652 8570
rect 11888 8560 11940 8566
rect 11888 8502 11940 8508
rect 11900 7834 11928 8502
rect 12912 7886 12940 8570
rect 11808 7806 11928 7834
rect 12900 7880 12952 7886
rect 12900 7822 12952 7828
rect 11808 7546 11836 7806
rect 12256 7744 12308 7750
rect 12256 7686 12308 7692
rect 12900 7744 12952 7750
rect 12900 7686 12952 7692
rect 11896 7644 12204 7653
rect 11896 7642 11902 7644
rect 11958 7642 11982 7644
rect 12038 7642 12062 7644
rect 12118 7642 12142 7644
rect 12198 7642 12204 7644
rect 11958 7590 11960 7642
rect 12140 7590 12142 7642
rect 11896 7588 11902 7590
rect 11958 7588 11982 7590
rect 12038 7588 12062 7590
rect 12118 7588 12142 7590
rect 12198 7588 12204 7590
rect 11896 7579 12204 7588
rect 11796 7540 11848 7546
rect 11796 7482 11848 7488
rect 12268 7410 12296 7686
rect 12256 7404 12308 7410
rect 12256 7346 12308 7352
rect 12624 7404 12676 7410
rect 12624 7346 12676 7352
rect 11796 6996 11848 7002
rect 11796 6938 11848 6944
rect 11612 6656 11664 6662
rect 11612 6598 11664 6604
rect 10968 6316 11020 6322
rect 10968 6258 11020 6264
rect 10140 6180 10192 6186
rect 10140 6122 10192 6128
rect 10876 6180 10928 6186
rect 10876 6122 10928 6128
rect 10888 5370 10916 6122
rect 11808 5914 11836 6938
rect 11896 6556 12204 6565
rect 11896 6554 11902 6556
rect 11958 6554 11982 6556
rect 12038 6554 12062 6556
rect 12118 6554 12142 6556
rect 12198 6554 12204 6556
rect 11958 6502 11960 6554
rect 12140 6502 12142 6554
rect 11896 6500 11902 6502
rect 11958 6500 11982 6502
rect 12038 6500 12062 6502
rect 12118 6500 12142 6502
rect 12198 6500 12204 6502
rect 11896 6491 12204 6500
rect 12532 6384 12584 6390
rect 12532 6326 12584 6332
rect 11796 5908 11848 5914
rect 11796 5850 11848 5856
rect 10876 5364 10928 5370
rect 10876 5306 10928 5312
rect 10416 5296 10468 5302
rect 10416 5238 10468 5244
rect 10428 4826 10456 5238
rect 10416 4820 10468 4826
rect 10416 4762 10468 4768
rect 11808 4690 11836 5850
rect 12544 5710 12572 6326
rect 12636 5710 12664 7346
rect 12912 7206 12940 7686
rect 12900 7200 12952 7206
rect 12900 7142 12952 7148
rect 12532 5704 12584 5710
rect 12532 5646 12584 5652
rect 12624 5704 12676 5710
rect 12624 5646 12676 5652
rect 12716 5568 12768 5574
rect 12716 5510 12768 5516
rect 12808 5568 12860 5574
rect 12808 5510 12860 5516
rect 11896 5468 12204 5477
rect 11896 5466 11902 5468
rect 11958 5466 11982 5468
rect 12038 5466 12062 5468
rect 12118 5466 12142 5468
rect 12198 5466 12204 5468
rect 11958 5414 11960 5466
rect 12140 5414 12142 5466
rect 11896 5412 11902 5414
rect 11958 5412 11982 5414
rect 12038 5412 12062 5414
rect 12118 5412 12142 5414
rect 12198 5412 12204 5414
rect 11896 5403 12204 5412
rect 12728 5234 12756 5510
rect 12820 5302 12848 5510
rect 12808 5296 12860 5302
rect 12808 5238 12860 5244
rect 12716 5228 12768 5234
rect 12716 5170 12768 5176
rect 12912 5114 12940 7142
rect 13280 6390 13308 9590
rect 13360 9580 13412 9586
rect 13360 9522 13412 9528
rect 13372 9450 13400 9522
rect 13360 9444 13412 9450
rect 13360 9386 13412 9392
rect 13372 7562 13400 9386
rect 13464 8974 13492 9658
rect 13556 9042 13584 9658
rect 14096 9580 14148 9586
rect 14096 9522 14148 9528
rect 14004 9444 14056 9450
rect 14004 9386 14056 9392
rect 13820 9376 13872 9382
rect 14016 9330 14044 9386
rect 13872 9324 14044 9330
rect 13820 9318 14044 9324
rect 13832 9302 14044 9318
rect 14108 9110 14136 9522
rect 14924 9512 14976 9518
rect 14924 9454 14976 9460
rect 14096 9104 14148 9110
rect 14096 9046 14148 9052
rect 13544 9036 13596 9042
rect 13544 8978 13596 8984
rect 13452 8968 13504 8974
rect 13452 8910 13504 8916
rect 13556 7954 13584 8978
rect 14936 8974 14964 9454
rect 14464 8968 14516 8974
rect 14464 8910 14516 8916
rect 14924 8968 14976 8974
rect 14924 8910 14976 8916
rect 13544 7948 13596 7954
rect 13544 7890 13596 7896
rect 13372 7534 13492 7562
rect 14476 7546 14504 8910
rect 14936 7886 14964 8910
rect 15396 8430 15424 11086
rect 15384 8424 15436 8430
rect 15384 8366 15436 8372
rect 15488 7886 15516 14282
rect 15672 14278 15700 14350
rect 15660 14272 15712 14278
rect 15660 14214 15712 14220
rect 16592 13977 16620 16934
rect 17236 16522 17264 17326
rect 19352 17202 19380 19200
rect 19340 17196 19392 17202
rect 19340 17138 19392 17144
rect 17370 16892 17678 16901
rect 17370 16890 17376 16892
rect 17432 16890 17456 16892
rect 17512 16890 17536 16892
rect 17592 16890 17616 16892
rect 17672 16890 17678 16892
rect 17432 16838 17434 16890
rect 17614 16838 17616 16890
rect 17370 16836 17376 16838
rect 17432 16836 17456 16838
rect 17512 16836 17536 16838
rect 17592 16836 17616 16838
rect 17672 16836 17678 16838
rect 17370 16827 17678 16836
rect 20640 16590 20668 19200
rect 22572 17202 22600 19200
rect 22843 17436 23151 17445
rect 22843 17434 22849 17436
rect 22905 17434 22929 17436
rect 22985 17434 23009 17436
rect 23065 17434 23089 17436
rect 23145 17434 23151 17436
rect 22905 17382 22907 17434
rect 23087 17382 23089 17434
rect 22843 17380 22849 17382
rect 22905 17380 22929 17382
rect 22985 17380 23009 17382
rect 23065 17380 23089 17382
rect 23145 17380 23151 17382
rect 22843 17371 23151 17380
rect 23860 17202 23888 19200
rect 25792 17202 25820 19200
rect 27724 17202 27752 19200
rect 29012 17202 29040 19200
rect 30944 17202 30972 19200
rect 32232 17202 32260 19200
rect 34164 19106 34192 19200
rect 34152 19100 34204 19106
rect 34152 19042 34204 19048
rect 35072 19100 35124 19106
rect 35072 19042 35124 19048
rect 33790 17436 34098 17445
rect 33790 17434 33796 17436
rect 33852 17434 33876 17436
rect 33932 17434 33956 17436
rect 34012 17434 34036 17436
rect 34092 17434 34098 17436
rect 33852 17382 33854 17434
rect 34034 17382 34036 17434
rect 33790 17380 33796 17382
rect 33852 17380 33876 17382
rect 33932 17380 33956 17382
rect 34012 17380 34036 17382
rect 34092 17380 34098 17382
rect 33790 17371 34098 17380
rect 35084 17202 35112 19042
rect 35452 17202 35480 19200
rect 37384 17202 37412 19200
rect 38672 17270 38700 19200
rect 38660 17264 38712 17270
rect 38660 17206 38712 17212
rect 22560 17196 22612 17202
rect 22560 17138 22612 17144
rect 23848 17196 23900 17202
rect 23848 17138 23900 17144
rect 25780 17196 25832 17202
rect 25780 17138 25832 17144
rect 27712 17196 27764 17202
rect 27712 17138 27764 17144
rect 29000 17196 29052 17202
rect 29000 17138 29052 17144
rect 30932 17196 30984 17202
rect 30932 17138 30984 17144
rect 32220 17196 32272 17202
rect 32220 17138 32272 17144
rect 35072 17196 35124 17202
rect 35072 17138 35124 17144
rect 35440 17196 35492 17202
rect 35440 17138 35492 17144
rect 37372 17196 37424 17202
rect 37372 17138 37424 17144
rect 32588 17128 32640 17134
rect 32588 17070 32640 17076
rect 23756 16992 23808 16998
rect 23756 16934 23808 16940
rect 31300 16992 31352 16998
rect 31300 16934 31352 16940
rect 19524 16584 19576 16590
rect 19524 16526 19576 16532
rect 20628 16584 20680 16590
rect 20628 16526 20680 16532
rect 17224 16516 17276 16522
rect 17224 16458 17276 16464
rect 17370 15804 17678 15813
rect 17370 15802 17376 15804
rect 17432 15802 17456 15804
rect 17512 15802 17536 15804
rect 17592 15802 17616 15804
rect 17672 15802 17678 15804
rect 17432 15750 17434 15802
rect 17614 15750 17616 15802
rect 17370 15748 17376 15750
rect 17432 15748 17456 15750
rect 17512 15748 17536 15750
rect 17592 15748 17616 15750
rect 17672 15748 17678 15750
rect 17370 15739 17678 15748
rect 19536 15706 19564 16526
rect 22843 16348 23151 16357
rect 22843 16346 22849 16348
rect 22905 16346 22929 16348
rect 22985 16346 23009 16348
rect 23065 16346 23089 16348
rect 23145 16346 23151 16348
rect 22905 16294 22907 16346
rect 23087 16294 23089 16346
rect 22843 16292 22849 16294
rect 22905 16292 22929 16294
rect 22985 16292 23009 16294
rect 23065 16292 23089 16294
rect 23145 16292 23151 16294
rect 22843 16283 23151 16292
rect 19524 15700 19576 15706
rect 19524 15642 19576 15648
rect 17132 15496 17184 15502
rect 17132 15438 17184 15444
rect 17776 15496 17828 15502
rect 17776 15438 17828 15444
rect 16578 13968 16634 13977
rect 15568 13932 15620 13938
rect 16578 13903 16634 13912
rect 15568 13874 15620 13880
rect 15580 13530 15608 13874
rect 15568 13524 15620 13530
rect 15568 13466 15620 13472
rect 16304 11076 16356 11082
rect 16304 11018 16356 11024
rect 16028 11008 16080 11014
rect 16028 10950 16080 10956
rect 16040 10674 16068 10950
rect 16028 10668 16080 10674
rect 16028 10610 16080 10616
rect 15660 10464 15712 10470
rect 15660 10406 15712 10412
rect 15568 8900 15620 8906
rect 15568 8842 15620 8848
rect 14924 7880 14976 7886
rect 14924 7822 14976 7828
rect 15476 7880 15528 7886
rect 15476 7822 15528 7828
rect 13360 7404 13412 7410
rect 13360 7346 13412 7352
rect 13372 7002 13400 7346
rect 13360 6996 13412 7002
rect 13360 6938 13412 6944
rect 13464 6866 13492 7534
rect 14464 7540 14516 7546
rect 14464 7482 14516 7488
rect 14936 7478 14964 7822
rect 14924 7472 14976 7478
rect 14924 7414 14976 7420
rect 14936 6866 14964 7414
rect 15476 7404 15528 7410
rect 15476 7346 15528 7352
rect 15016 7200 15068 7206
rect 15016 7142 15068 7148
rect 15108 7200 15160 7206
rect 15108 7142 15160 7148
rect 13452 6860 13504 6866
rect 13452 6802 13504 6808
rect 14924 6860 14976 6866
rect 14924 6802 14976 6808
rect 13268 6384 13320 6390
rect 13268 6326 13320 6332
rect 13360 5704 13412 5710
rect 13360 5646 13412 5652
rect 13372 5545 13400 5646
rect 13358 5536 13414 5545
rect 13280 5494 13358 5522
rect 13280 5370 13308 5494
rect 13358 5471 13414 5480
rect 13268 5364 13320 5370
rect 13464 5352 13492 6802
rect 14188 6724 14240 6730
rect 14188 6666 14240 6672
rect 13544 5704 13596 5710
rect 13544 5646 13596 5652
rect 13820 5704 13872 5710
rect 13820 5646 13872 5652
rect 13268 5306 13320 5312
rect 13372 5324 13492 5352
rect 12820 5086 12940 5114
rect 12164 5024 12216 5030
rect 12164 4966 12216 4972
rect 11796 4684 11848 4690
rect 11796 4626 11848 4632
rect 9864 4616 9916 4622
rect 9864 4558 9916 4564
rect 9876 4146 9904 4558
rect 12176 4554 12204 4966
rect 12716 4684 12768 4690
rect 12716 4626 12768 4632
rect 12164 4548 12216 4554
rect 12164 4490 12216 4496
rect 11896 4380 12204 4389
rect 11896 4378 11902 4380
rect 11958 4378 11982 4380
rect 12038 4378 12062 4380
rect 12118 4378 12142 4380
rect 12198 4378 12204 4380
rect 11958 4326 11960 4378
rect 12140 4326 12142 4378
rect 11896 4324 11902 4326
rect 11958 4324 11982 4326
rect 12038 4324 12062 4326
rect 12118 4324 12142 4326
rect 12198 4324 12204 4326
rect 11896 4315 12204 4324
rect 12728 4282 12756 4626
rect 12716 4276 12768 4282
rect 12716 4218 12768 4224
rect 9864 4140 9916 4146
rect 9864 4082 9916 4088
rect 11896 3292 12204 3301
rect 11896 3290 11902 3292
rect 11958 3290 11982 3292
rect 12038 3290 12062 3292
rect 12118 3290 12142 3292
rect 12198 3290 12204 3292
rect 11958 3238 11960 3290
rect 12140 3238 12142 3290
rect 11896 3236 11902 3238
rect 11958 3236 11982 3238
rect 12038 3236 12062 3238
rect 12118 3236 12142 3238
rect 12198 3236 12204 3238
rect 11896 3227 12204 3236
rect 9312 3188 9364 3194
rect 9312 3130 9364 3136
rect 7196 3052 7248 3058
rect 7196 2994 7248 3000
rect 9680 2984 9732 2990
rect 9680 2926 9732 2932
rect 6423 2748 6731 2757
rect 6423 2746 6429 2748
rect 6485 2746 6509 2748
rect 6565 2746 6589 2748
rect 6645 2746 6669 2748
rect 6725 2746 6731 2748
rect 6485 2694 6487 2746
rect 6667 2694 6669 2746
rect 6423 2692 6429 2694
rect 6485 2692 6509 2694
rect 6565 2692 6589 2694
rect 6645 2692 6669 2694
rect 6725 2692 6731 2694
rect 6423 2683 6731 2692
rect 7748 2440 7800 2446
rect 7748 2382 7800 2388
rect 6288 1686 6500 1714
rect 6472 800 6500 1686
rect 7760 800 7788 2382
rect 9692 800 9720 2926
rect 12820 2650 12848 5086
rect 12900 5024 12952 5030
rect 12900 4966 12952 4972
rect 12912 4146 12940 4966
rect 13280 4758 13308 5306
rect 13372 4826 13400 5324
rect 13556 5250 13584 5646
rect 13832 5556 13860 5646
rect 13740 5528 13860 5556
rect 13740 5302 13768 5528
rect 13464 5234 13584 5250
rect 13728 5296 13780 5302
rect 13728 5238 13780 5244
rect 13452 5228 13584 5234
rect 13504 5222 13584 5228
rect 13452 5170 13504 5176
rect 13360 4820 13412 4826
rect 13360 4762 13412 4768
rect 13268 4752 13320 4758
rect 13268 4694 13320 4700
rect 13556 4554 13584 5222
rect 13544 4548 13596 4554
rect 13544 4490 13596 4496
rect 12900 4140 12952 4146
rect 12900 4082 12952 4088
rect 13740 3534 13768 5238
rect 13820 5160 13872 5166
rect 13820 5102 13872 5108
rect 13832 4282 13860 5102
rect 13820 4276 13872 4282
rect 13820 4218 13872 4224
rect 13728 3528 13780 3534
rect 13728 3470 13780 3476
rect 13636 3392 13688 3398
rect 13636 3334 13688 3340
rect 13648 3058 13676 3334
rect 13636 3052 13688 3058
rect 13636 2994 13688 3000
rect 12808 2644 12860 2650
rect 12808 2586 12860 2592
rect 11060 2440 11112 2446
rect 11060 2382 11112 2388
rect 12900 2440 12952 2446
rect 12900 2382 12952 2388
rect 11072 898 11100 2382
rect 11896 2204 12204 2213
rect 11896 2202 11902 2204
rect 11958 2202 11982 2204
rect 12038 2202 12062 2204
rect 12118 2202 12142 2204
rect 12198 2202 12204 2204
rect 11958 2150 11960 2202
rect 12140 2150 12142 2202
rect 11896 2148 11902 2150
rect 11958 2148 11982 2150
rect 12038 2148 12062 2150
rect 12118 2148 12142 2150
rect 12198 2148 12204 2150
rect 11896 2139 12204 2148
rect 10980 870 11100 898
rect 10980 800 11008 870
rect 12912 800 12940 2382
rect 14200 800 14228 6666
rect 14556 6656 14608 6662
rect 14556 6598 14608 6604
rect 14462 5672 14518 5681
rect 14568 5642 14596 6598
rect 14936 6390 14964 6802
rect 15028 6730 15056 7142
rect 15120 6798 15148 7142
rect 15108 6792 15160 6798
rect 15108 6734 15160 6740
rect 15016 6724 15068 6730
rect 15016 6666 15068 6672
rect 15028 6390 15056 6666
rect 14924 6384 14976 6390
rect 14924 6326 14976 6332
rect 15016 6384 15068 6390
rect 15016 6326 15068 6332
rect 14936 5710 14964 6326
rect 15488 6254 15516 7346
rect 15580 7342 15608 8842
rect 15672 8566 15700 10406
rect 16040 10266 16068 10610
rect 16028 10260 16080 10266
rect 16028 10202 16080 10208
rect 16316 9450 16344 11018
rect 16488 10600 16540 10606
rect 16488 10542 16540 10548
rect 16500 10266 16528 10542
rect 16488 10260 16540 10266
rect 16488 10202 16540 10208
rect 16592 10130 16620 13903
rect 16948 12232 17000 12238
rect 16948 12174 17000 12180
rect 16960 11830 16988 12174
rect 16948 11824 17000 11830
rect 16948 11766 17000 11772
rect 17144 11218 17172 15438
rect 17788 15162 17816 15438
rect 19892 15428 19944 15434
rect 19892 15370 19944 15376
rect 19800 15360 19852 15366
rect 19800 15302 19852 15308
rect 17776 15156 17828 15162
rect 17776 15098 17828 15104
rect 19708 15088 19760 15094
rect 19708 15030 19760 15036
rect 17224 15020 17276 15026
rect 17224 14962 17276 14968
rect 17868 15020 17920 15026
rect 17868 14962 17920 14968
rect 17236 14618 17264 14962
rect 17370 14716 17678 14725
rect 17370 14714 17376 14716
rect 17432 14714 17456 14716
rect 17512 14714 17536 14716
rect 17592 14714 17616 14716
rect 17672 14714 17678 14716
rect 17432 14662 17434 14714
rect 17614 14662 17616 14714
rect 17370 14660 17376 14662
rect 17432 14660 17456 14662
rect 17512 14660 17536 14662
rect 17592 14660 17616 14662
rect 17672 14660 17678 14662
rect 17370 14651 17678 14660
rect 17224 14612 17276 14618
rect 17224 14554 17276 14560
rect 17880 13870 17908 14962
rect 19720 14414 19748 15030
rect 19812 15026 19840 15302
rect 19800 15020 19852 15026
rect 19800 14962 19852 14968
rect 19904 14550 19932 15370
rect 19984 15360 20036 15366
rect 19984 15302 20036 15308
rect 19996 15162 20024 15302
rect 22843 15260 23151 15269
rect 22843 15258 22849 15260
rect 22905 15258 22929 15260
rect 22985 15258 23009 15260
rect 23065 15258 23089 15260
rect 23145 15258 23151 15260
rect 22905 15206 22907 15258
rect 23087 15206 23089 15258
rect 22843 15204 22849 15206
rect 22905 15204 22929 15206
rect 22985 15204 23009 15206
rect 23065 15204 23089 15206
rect 23145 15204 23151 15206
rect 22843 15195 23151 15204
rect 19984 15156 20036 15162
rect 19984 15098 20036 15104
rect 22100 15020 22152 15026
rect 22100 14962 22152 14968
rect 19892 14544 19944 14550
rect 19892 14486 19944 14492
rect 19984 14476 20036 14482
rect 19984 14418 20036 14424
rect 20996 14476 21048 14482
rect 20996 14418 21048 14424
rect 19708 14408 19760 14414
rect 19708 14350 19760 14356
rect 18512 14272 18564 14278
rect 18512 14214 18564 14220
rect 19892 14272 19944 14278
rect 19892 14214 19944 14220
rect 17868 13864 17920 13870
rect 17868 13806 17920 13812
rect 17370 13628 17678 13637
rect 17370 13626 17376 13628
rect 17432 13626 17456 13628
rect 17512 13626 17536 13628
rect 17592 13626 17616 13628
rect 17672 13626 17678 13628
rect 17432 13574 17434 13626
rect 17614 13574 17616 13626
rect 17370 13572 17376 13574
rect 17432 13572 17456 13574
rect 17512 13572 17536 13574
rect 17592 13572 17616 13574
rect 17672 13572 17678 13574
rect 17370 13563 17678 13572
rect 17880 13258 17908 13806
rect 18524 13530 18552 14214
rect 19904 14074 19932 14214
rect 19892 14068 19944 14074
rect 19892 14010 19944 14016
rect 19340 13932 19392 13938
rect 19340 13874 19392 13880
rect 19352 13530 19380 13874
rect 18512 13524 18564 13530
rect 18512 13466 18564 13472
rect 19340 13524 19392 13530
rect 19340 13466 19392 13472
rect 19996 13394 20024 14418
rect 20628 14340 20680 14346
rect 20628 14282 20680 14288
rect 20352 13728 20404 13734
rect 20352 13670 20404 13676
rect 19984 13388 20036 13394
rect 19984 13330 20036 13336
rect 20364 13326 20392 13670
rect 20352 13320 20404 13326
rect 20352 13262 20404 13268
rect 17776 13252 17828 13258
rect 17776 13194 17828 13200
rect 17868 13252 17920 13258
rect 17868 13194 17920 13200
rect 17370 12540 17678 12549
rect 17370 12538 17376 12540
rect 17432 12538 17456 12540
rect 17512 12538 17536 12540
rect 17592 12538 17616 12540
rect 17672 12538 17678 12540
rect 17432 12486 17434 12538
rect 17614 12486 17616 12538
rect 17370 12484 17376 12486
rect 17432 12484 17456 12486
rect 17512 12484 17536 12486
rect 17592 12484 17616 12486
rect 17672 12484 17678 12486
rect 17370 12475 17678 12484
rect 17788 12442 17816 13194
rect 17880 12918 17908 13194
rect 18880 13184 18932 13190
rect 18880 13126 18932 13132
rect 18892 12986 18920 13126
rect 18880 12980 18932 12986
rect 18880 12922 18932 12928
rect 17868 12912 17920 12918
rect 17868 12854 17920 12860
rect 18052 12844 18104 12850
rect 18052 12786 18104 12792
rect 19432 12844 19484 12850
rect 19432 12786 19484 12792
rect 17776 12436 17828 12442
rect 17776 12378 17828 12384
rect 17776 12232 17828 12238
rect 17776 12174 17828 12180
rect 17224 11756 17276 11762
rect 17224 11698 17276 11704
rect 17132 11212 17184 11218
rect 17132 11154 17184 11160
rect 17236 10810 17264 11698
rect 17370 11452 17678 11461
rect 17370 11450 17376 11452
rect 17432 11450 17456 11452
rect 17512 11450 17536 11452
rect 17592 11450 17616 11452
rect 17672 11450 17678 11452
rect 17432 11398 17434 11450
rect 17614 11398 17616 11450
rect 17370 11396 17376 11398
rect 17432 11396 17456 11398
rect 17512 11396 17536 11398
rect 17592 11396 17616 11398
rect 17672 11396 17678 11398
rect 17370 11387 17678 11396
rect 17788 11354 17816 12174
rect 18064 11898 18092 12786
rect 19444 11898 19472 12786
rect 20640 12442 20668 14282
rect 21008 13870 21036 14418
rect 21916 14272 21968 14278
rect 21916 14214 21968 14220
rect 21928 14006 21956 14214
rect 21916 14000 21968 14006
rect 21916 13942 21968 13948
rect 22112 13938 22140 14962
rect 22376 14816 22428 14822
rect 22376 14758 22428 14764
rect 22192 14408 22244 14414
rect 22192 14350 22244 14356
rect 22100 13932 22152 13938
rect 22100 13874 22152 13880
rect 20996 13864 21048 13870
rect 20996 13806 21048 13812
rect 22204 13530 22232 14350
rect 22192 13524 22244 13530
rect 22192 13466 22244 13472
rect 22008 13184 22060 13190
rect 22008 13126 22060 13132
rect 20720 12912 20772 12918
rect 20720 12854 20772 12860
rect 20628 12436 20680 12442
rect 20628 12378 20680 12384
rect 19524 12096 19576 12102
rect 19524 12038 19576 12044
rect 19536 11898 19564 12038
rect 18052 11892 18104 11898
rect 18052 11834 18104 11840
rect 19432 11892 19484 11898
rect 19432 11834 19484 11840
rect 19524 11892 19576 11898
rect 19524 11834 19576 11840
rect 18236 11756 18288 11762
rect 18236 11698 18288 11704
rect 18880 11756 18932 11762
rect 18880 11698 18932 11704
rect 17776 11348 17828 11354
rect 17776 11290 17828 11296
rect 18248 11286 18276 11698
rect 18236 11280 18288 11286
rect 18236 11222 18288 11228
rect 18328 11212 18380 11218
rect 18328 11154 18380 11160
rect 18236 11144 18288 11150
rect 18236 11086 18288 11092
rect 17224 10804 17276 10810
rect 17224 10746 17276 10752
rect 16580 10124 16632 10130
rect 16580 10066 16632 10072
rect 17236 10062 17264 10746
rect 17958 10568 18014 10577
rect 17958 10503 18014 10512
rect 17370 10364 17678 10373
rect 17370 10362 17376 10364
rect 17432 10362 17456 10364
rect 17512 10362 17536 10364
rect 17592 10362 17616 10364
rect 17672 10362 17678 10364
rect 17432 10310 17434 10362
rect 17614 10310 17616 10362
rect 17370 10308 17376 10310
rect 17432 10308 17456 10310
rect 17512 10308 17536 10310
rect 17592 10308 17616 10310
rect 17672 10308 17678 10310
rect 17370 10299 17678 10308
rect 17776 10124 17828 10130
rect 17776 10066 17828 10072
rect 17224 10056 17276 10062
rect 17224 9998 17276 10004
rect 17788 9722 17816 10066
rect 17972 10062 18000 10503
rect 17960 10056 18012 10062
rect 17960 9998 18012 10004
rect 17776 9716 17828 9722
rect 17776 9658 17828 9664
rect 17132 9580 17184 9586
rect 17184 9540 17264 9568
rect 17132 9522 17184 9528
rect 16856 9512 16908 9518
rect 16856 9454 16908 9460
rect 16304 9444 16356 9450
rect 16304 9386 16356 9392
rect 16868 8974 16896 9454
rect 17236 9178 17264 9540
rect 17370 9276 17678 9285
rect 17370 9274 17376 9276
rect 17432 9274 17456 9276
rect 17512 9274 17536 9276
rect 17592 9274 17616 9276
rect 17672 9274 17678 9276
rect 17432 9222 17434 9274
rect 17614 9222 17616 9274
rect 17370 9220 17376 9222
rect 17432 9220 17456 9222
rect 17512 9220 17536 9222
rect 17592 9220 17616 9222
rect 17672 9220 17678 9222
rect 17370 9211 17678 9220
rect 17224 9172 17276 9178
rect 17224 9114 17276 9120
rect 16856 8968 16908 8974
rect 16856 8910 16908 8916
rect 16868 8566 16896 8910
rect 15660 8560 15712 8566
rect 15660 8502 15712 8508
rect 16856 8560 16908 8566
rect 16856 8502 16908 8508
rect 16212 8492 16264 8498
rect 16212 8434 16264 8440
rect 15660 8424 15712 8430
rect 15660 8366 15712 8372
rect 15672 7886 15700 8366
rect 16224 8090 16252 8434
rect 16856 8356 16908 8362
rect 16856 8298 16908 8304
rect 16212 8084 16264 8090
rect 16212 8026 16264 8032
rect 15660 7880 15712 7886
rect 15660 7822 15712 7828
rect 15672 7342 15700 7822
rect 16224 7410 16252 8026
rect 16868 7886 16896 8298
rect 16856 7880 16908 7886
rect 16856 7822 16908 7828
rect 16212 7404 16264 7410
rect 16212 7346 16264 7352
rect 15568 7336 15620 7342
rect 15568 7278 15620 7284
rect 15660 7336 15712 7342
rect 15660 7278 15712 7284
rect 15672 7002 15700 7278
rect 15660 6996 15712 7002
rect 15660 6938 15712 6944
rect 15568 6724 15620 6730
rect 15568 6666 15620 6672
rect 15580 6458 15608 6666
rect 17236 6662 17264 9114
rect 17370 8188 17678 8197
rect 17370 8186 17376 8188
rect 17432 8186 17456 8188
rect 17512 8186 17536 8188
rect 17592 8186 17616 8188
rect 17672 8186 17678 8188
rect 17432 8134 17434 8186
rect 17614 8134 17616 8186
rect 17370 8132 17376 8134
rect 17432 8132 17456 8134
rect 17512 8132 17536 8134
rect 17592 8132 17616 8134
rect 17672 8132 17678 8134
rect 17370 8123 17678 8132
rect 17972 7818 18000 9998
rect 18248 9382 18276 11086
rect 18340 10062 18368 11154
rect 18604 10464 18656 10470
rect 18604 10406 18656 10412
rect 18616 10198 18644 10406
rect 18892 10266 18920 11698
rect 20076 11552 20128 11558
rect 20076 11494 20128 11500
rect 20088 11354 20116 11494
rect 20076 11348 20128 11354
rect 20076 11290 20128 11296
rect 20260 11280 20312 11286
rect 20260 11222 20312 11228
rect 19984 11212 20036 11218
rect 19984 11154 20036 11160
rect 19248 10804 19300 10810
rect 19248 10746 19300 10752
rect 18880 10260 18932 10266
rect 18880 10202 18932 10208
rect 18604 10192 18656 10198
rect 18604 10134 18656 10140
rect 18328 10056 18380 10062
rect 18328 9998 18380 10004
rect 18512 10056 18564 10062
rect 18512 9998 18564 10004
rect 18236 9376 18288 9382
rect 18236 9318 18288 9324
rect 18524 9178 18552 9998
rect 19260 9926 19288 10746
rect 19708 10532 19760 10538
rect 19708 10474 19760 10480
rect 19720 10062 19748 10474
rect 19708 10056 19760 10062
rect 19706 10024 19708 10033
rect 19760 10024 19762 10033
rect 19706 9959 19762 9968
rect 19248 9920 19300 9926
rect 19248 9862 19300 9868
rect 19340 9376 19392 9382
rect 19340 9318 19392 9324
rect 18512 9172 18564 9178
rect 18512 9114 18564 9120
rect 19352 9110 19380 9318
rect 19340 9104 19392 9110
rect 19340 9046 19392 9052
rect 19892 9036 19944 9042
rect 19892 8978 19944 8984
rect 18236 8968 18288 8974
rect 18236 8910 18288 8916
rect 18052 8832 18104 8838
rect 18052 8774 18104 8780
rect 18064 8498 18092 8774
rect 18052 8492 18104 8498
rect 18052 8434 18104 8440
rect 18248 8090 18276 8910
rect 19524 8832 19576 8838
rect 19524 8774 19576 8780
rect 18604 8288 18656 8294
rect 18604 8230 18656 8236
rect 18236 8084 18288 8090
rect 18236 8026 18288 8032
rect 18616 7886 18644 8230
rect 19536 7886 19564 8774
rect 19708 8492 19760 8498
rect 19904 8480 19932 8978
rect 19760 8452 19932 8480
rect 19708 8434 19760 8440
rect 19904 7954 19932 8452
rect 19996 8430 20024 11154
rect 20272 10674 20300 11222
rect 20640 11218 20668 12378
rect 20732 11218 20760 12854
rect 22020 12714 22048 13126
rect 22008 12708 22060 12714
rect 22008 12650 22060 12656
rect 21364 12232 21416 12238
rect 21364 12174 21416 12180
rect 21456 12232 21508 12238
rect 21456 12174 21508 12180
rect 20996 12096 21048 12102
rect 20996 12038 21048 12044
rect 20904 11892 20956 11898
rect 20904 11834 20956 11840
rect 20916 11694 20944 11834
rect 20904 11688 20956 11694
rect 20904 11630 20956 11636
rect 20812 11552 20864 11558
rect 20812 11494 20864 11500
rect 20904 11552 20956 11558
rect 20904 11494 20956 11500
rect 20628 11212 20680 11218
rect 20628 11154 20680 11160
rect 20720 11212 20772 11218
rect 20720 11154 20772 11160
rect 20720 11076 20772 11082
rect 20720 11018 20772 11024
rect 20260 10668 20312 10674
rect 20260 10610 20312 10616
rect 20732 9382 20760 11018
rect 20824 10062 20852 11494
rect 20916 11014 20944 11494
rect 21008 11218 21036 12038
rect 21376 11898 21404 12174
rect 21088 11892 21140 11898
rect 21088 11834 21140 11840
rect 21364 11892 21416 11898
rect 21364 11834 21416 11840
rect 20996 11212 21048 11218
rect 20996 11154 21048 11160
rect 20904 11008 20956 11014
rect 20904 10950 20956 10956
rect 20996 11008 21048 11014
rect 20996 10950 21048 10956
rect 21008 10810 21036 10950
rect 20996 10804 21048 10810
rect 20996 10746 21048 10752
rect 20904 10260 20956 10266
rect 20904 10202 20956 10208
rect 20812 10056 20864 10062
rect 20812 9998 20864 10004
rect 20812 9648 20864 9654
rect 20812 9590 20864 9596
rect 20352 9376 20404 9382
rect 20352 9318 20404 9324
rect 20720 9376 20772 9382
rect 20720 9318 20772 9324
rect 20364 8974 20392 9318
rect 20168 8968 20220 8974
rect 20168 8910 20220 8916
rect 20352 8968 20404 8974
rect 20352 8910 20404 8916
rect 20180 8634 20208 8910
rect 20824 8906 20852 9590
rect 20916 9518 20944 10202
rect 20996 9920 21048 9926
rect 20996 9862 21048 9868
rect 21100 9908 21128 11834
rect 21180 11688 21232 11694
rect 21180 11630 21232 11636
rect 21192 10810 21220 11630
rect 21468 11558 21496 12174
rect 22100 12096 22152 12102
rect 22100 12038 22152 12044
rect 22008 11756 22060 11762
rect 22008 11698 22060 11704
rect 21456 11552 21508 11558
rect 21456 11494 21508 11500
rect 22020 11286 22048 11698
rect 22008 11280 22060 11286
rect 22008 11222 22060 11228
rect 22112 11150 22140 12038
rect 22284 11552 22336 11558
rect 22284 11494 22336 11500
rect 22100 11144 22152 11150
rect 22100 11086 22152 11092
rect 21180 10804 21232 10810
rect 21180 10746 21232 10752
rect 22192 10600 22244 10606
rect 22192 10542 22244 10548
rect 21272 10532 21324 10538
rect 21272 10474 21324 10480
rect 21284 9994 21312 10474
rect 21732 10192 21784 10198
rect 21732 10134 21784 10140
rect 21272 9988 21324 9994
rect 21272 9930 21324 9936
rect 21180 9920 21232 9926
rect 21100 9880 21180 9908
rect 21008 9518 21036 9862
rect 21100 9586 21128 9880
rect 21180 9862 21232 9868
rect 21088 9580 21140 9586
rect 21088 9522 21140 9528
rect 21180 9580 21232 9586
rect 21180 9522 21232 9528
rect 20904 9512 20956 9518
rect 20904 9454 20956 9460
rect 20996 9512 21048 9518
rect 20996 9454 21048 9460
rect 20812 8900 20864 8906
rect 20812 8842 20864 8848
rect 21192 8634 21220 9522
rect 21744 9518 21772 10134
rect 22204 10130 22232 10542
rect 22192 10124 22244 10130
rect 22192 10066 22244 10072
rect 22006 9752 22062 9761
rect 22006 9687 22008 9696
rect 22060 9687 22062 9696
rect 22008 9658 22060 9664
rect 22100 9580 22152 9586
rect 22100 9522 22152 9528
rect 21732 9512 21784 9518
rect 21732 9454 21784 9460
rect 22112 9382 22140 9522
rect 22100 9376 22152 9382
rect 22100 9318 22152 9324
rect 20168 8628 20220 8634
rect 20168 8570 20220 8576
rect 21180 8628 21232 8634
rect 21180 8570 21232 8576
rect 20904 8492 20956 8498
rect 20904 8434 20956 8440
rect 21272 8492 21324 8498
rect 21272 8434 21324 8440
rect 19984 8424 20036 8430
rect 19984 8366 20036 8372
rect 20076 8424 20128 8430
rect 20076 8366 20128 8372
rect 20088 8090 20116 8366
rect 20076 8084 20128 8090
rect 20076 8026 20128 8032
rect 19892 7948 19944 7954
rect 19892 7890 19944 7896
rect 18604 7880 18656 7886
rect 18604 7822 18656 7828
rect 19524 7880 19576 7886
rect 19524 7822 19576 7828
rect 17960 7812 18012 7818
rect 17960 7754 18012 7760
rect 17960 7200 18012 7206
rect 17960 7142 18012 7148
rect 17370 7100 17678 7109
rect 17370 7098 17376 7100
rect 17432 7098 17456 7100
rect 17512 7098 17536 7100
rect 17592 7098 17616 7100
rect 17672 7098 17678 7100
rect 17432 7046 17434 7098
rect 17614 7046 17616 7098
rect 17370 7044 17376 7046
rect 17432 7044 17456 7046
rect 17512 7044 17536 7046
rect 17592 7044 17616 7046
rect 17672 7044 17678 7046
rect 17370 7035 17678 7044
rect 17776 6724 17828 6730
rect 17776 6666 17828 6672
rect 17132 6656 17184 6662
rect 17132 6598 17184 6604
rect 17224 6656 17276 6662
rect 17224 6598 17276 6604
rect 15568 6452 15620 6458
rect 15568 6394 15620 6400
rect 17144 6322 17172 6598
rect 17132 6316 17184 6322
rect 17132 6258 17184 6264
rect 15476 6248 15528 6254
rect 15476 6190 15528 6196
rect 15488 5914 15516 6190
rect 17370 6012 17678 6021
rect 17370 6010 17376 6012
rect 17432 6010 17456 6012
rect 17512 6010 17536 6012
rect 17592 6010 17616 6012
rect 17672 6010 17678 6012
rect 17432 5958 17434 6010
rect 17614 5958 17616 6010
rect 17370 5956 17376 5958
rect 17432 5956 17456 5958
rect 17512 5956 17536 5958
rect 17592 5956 17616 5958
rect 17672 5956 17678 5958
rect 17370 5947 17678 5956
rect 15476 5908 15528 5914
rect 15476 5850 15528 5856
rect 16120 5840 16172 5846
rect 16120 5782 16172 5788
rect 15752 5772 15804 5778
rect 15752 5714 15804 5720
rect 14924 5704 14976 5710
rect 14924 5646 14976 5652
rect 14462 5607 14518 5616
rect 14556 5636 14608 5642
rect 14476 5574 14504 5607
rect 14556 5578 14608 5584
rect 14464 5568 14516 5574
rect 14464 5510 14516 5516
rect 14476 4622 14504 5510
rect 15764 5234 15792 5714
rect 15844 5568 15896 5574
rect 15844 5510 15896 5516
rect 15856 5302 15884 5510
rect 15844 5296 15896 5302
rect 15844 5238 15896 5244
rect 15752 5228 15804 5234
rect 15752 5170 15804 5176
rect 16132 5166 16160 5782
rect 17788 5710 17816 6666
rect 17868 6656 17920 6662
rect 17868 6598 17920 6604
rect 16304 5704 16356 5710
rect 16304 5646 16356 5652
rect 17684 5704 17736 5710
rect 17684 5646 17736 5652
rect 17776 5704 17828 5710
rect 17776 5646 17828 5652
rect 15844 5160 15896 5166
rect 15842 5128 15844 5137
rect 15936 5160 15988 5166
rect 15896 5128 15898 5137
rect 15936 5102 15988 5108
rect 16120 5160 16172 5166
rect 16120 5102 16172 5108
rect 15842 5063 15898 5072
rect 15948 4690 15976 5102
rect 16316 4826 16344 5646
rect 16580 5636 16632 5642
rect 16580 5578 16632 5584
rect 16304 4820 16356 4826
rect 16304 4762 16356 4768
rect 16592 4690 16620 5578
rect 16948 5296 17000 5302
rect 16948 5238 17000 5244
rect 16960 5166 16988 5238
rect 17696 5234 17724 5646
rect 17684 5228 17736 5234
rect 17684 5170 17736 5176
rect 16948 5160 17000 5166
rect 16948 5102 17000 5108
rect 15936 4684 15988 4690
rect 15936 4626 15988 4632
rect 16580 4684 16632 4690
rect 16580 4626 16632 4632
rect 14464 4616 14516 4622
rect 14464 4558 14516 4564
rect 15108 4480 15160 4486
rect 15108 4422 15160 4428
rect 15120 4146 15148 4422
rect 16960 4282 16988 5102
rect 17776 5024 17828 5030
rect 17776 4966 17828 4972
rect 17370 4924 17678 4933
rect 17370 4922 17376 4924
rect 17432 4922 17456 4924
rect 17512 4922 17536 4924
rect 17592 4922 17616 4924
rect 17672 4922 17678 4924
rect 17432 4870 17434 4922
rect 17614 4870 17616 4922
rect 17370 4868 17376 4870
rect 17432 4868 17456 4870
rect 17512 4868 17536 4870
rect 17592 4868 17616 4870
rect 17672 4868 17678 4870
rect 17370 4859 17678 4868
rect 17408 4548 17460 4554
rect 17408 4490 17460 4496
rect 17420 4282 17448 4490
rect 16948 4276 17000 4282
rect 16948 4218 17000 4224
rect 17408 4276 17460 4282
rect 17408 4218 17460 4224
rect 17788 4146 17816 4966
rect 15108 4140 15160 4146
rect 15108 4082 15160 4088
rect 16856 4140 16908 4146
rect 16856 4082 16908 4088
rect 17776 4140 17828 4146
rect 17776 4082 17828 4088
rect 16580 3936 16632 3942
rect 16580 3878 16632 3884
rect 14832 3528 14884 3534
rect 14832 3470 14884 3476
rect 15384 3528 15436 3534
rect 15384 3470 15436 3476
rect 16120 3528 16172 3534
rect 16120 3470 16172 3476
rect 16212 3528 16264 3534
rect 16212 3470 16264 3476
rect 14844 3058 14872 3470
rect 15200 3392 15252 3398
rect 15200 3334 15252 3340
rect 15212 3126 15240 3334
rect 15200 3120 15252 3126
rect 15200 3062 15252 3068
rect 14832 3052 14884 3058
rect 14832 2994 14884 3000
rect 15396 2650 15424 3470
rect 16132 3194 16160 3470
rect 16120 3188 16172 3194
rect 16120 3130 16172 3136
rect 16224 3058 16252 3470
rect 16592 3466 16620 3878
rect 16580 3460 16632 3466
rect 16580 3402 16632 3408
rect 16212 3052 16264 3058
rect 16212 2994 16264 3000
rect 15384 2644 15436 2650
rect 15384 2586 15436 2592
rect 16120 2576 16172 2582
rect 16120 2518 16172 2524
rect 16132 800 16160 2518
rect 16868 2446 16896 4082
rect 17370 3836 17678 3845
rect 17370 3834 17376 3836
rect 17432 3834 17456 3836
rect 17512 3834 17536 3836
rect 17592 3834 17616 3836
rect 17672 3834 17678 3836
rect 17432 3782 17434 3834
rect 17614 3782 17616 3834
rect 17370 3780 17376 3782
rect 17432 3780 17456 3782
rect 17512 3780 17536 3782
rect 17592 3780 17616 3782
rect 17672 3780 17678 3782
rect 17370 3771 17678 3780
rect 17776 3392 17828 3398
rect 17776 3334 17828 3340
rect 17788 3058 17816 3334
rect 17776 3052 17828 3058
rect 17776 2994 17828 3000
rect 17132 2984 17184 2990
rect 17132 2926 17184 2932
rect 17144 2650 17172 2926
rect 17370 2748 17678 2757
rect 17370 2746 17376 2748
rect 17432 2746 17456 2748
rect 17512 2746 17536 2748
rect 17592 2746 17616 2748
rect 17672 2746 17678 2748
rect 17432 2694 17434 2746
rect 17614 2694 17616 2746
rect 17370 2692 17376 2694
rect 17432 2692 17456 2694
rect 17512 2692 17536 2694
rect 17592 2692 17616 2694
rect 17672 2692 17678 2694
rect 17370 2683 17678 2692
rect 17880 2650 17908 6598
rect 17972 6458 18000 7142
rect 18616 6866 18644 7822
rect 19904 7410 19932 7890
rect 19892 7404 19944 7410
rect 19892 7346 19944 7352
rect 20916 7274 20944 8434
rect 21284 7750 21312 8434
rect 22204 8430 22232 10066
rect 22296 9761 22324 11494
rect 22388 10690 22416 14758
rect 23768 14482 23796 16934
rect 28317 16892 28625 16901
rect 28317 16890 28323 16892
rect 28379 16890 28403 16892
rect 28459 16890 28483 16892
rect 28539 16890 28563 16892
rect 28619 16890 28625 16892
rect 28379 16838 28381 16890
rect 28561 16838 28563 16890
rect 28317 16836 28323 16838
rect 28379 16836 28403 16838
rect 28459 16836 28483 16838
rect 28539 16836 28563 16838
rect 28619 16836 28625 16838
rect 28317 16827 28625 16836
rect 28317 15804 28625 15813
rect 28317 15802 28323 15804
rect 28379 15802 28403 15804
rect 28459 15802 28483 15804
rect 28539 15802 28563 15804
rect 28619 15802 28625 15804
rect 28379 15750 28381 15802
rect 28561 15750 28563 15802
rect 28317 15748 28323 15750
rect 28379 15748 28403 15750
rect 28459 15748 28483 15750
rect 28539 15748 28563 15750
rect 28619 15748 28625 15750
rect 28317 15739 28625 15748
rect 25228 15496 25280 15502
rect 25228 15438 25280 15444
rect 25136 15360 25188 15366
rect 25136 15302 25188 15308
rect 25148 15026 25176 15302
rect 24860 15020 24912 15026
rect 24860 14962 24912 14968
rect 25136 15020 25188 15026
rect 25136 14962 25188 14968
rect 24400 14816 24452 14822
rect 24400 14758 24452 14764
rect 23756 14476 23808 14482
rect 23756 14418 23808 14424
rect 23848 14476 23900 14482
rect 23848 14418 23900 14424
rect 23662 14376 23718 14385
rect 23662 14311 23664 14320
rect 23716 14311 23718 14320
rect 23664 14282 23716 14288
rect 23572 14272 23624 14278
rect 23572 14214 23624 14220
rect 22843 14172 23151 14181
rect 22843 14170 22849 14172
rect 22905 14170 22929 14172
rect 22985 14170 23009 14172
rect 23065 14170 23089 14172
rect 23145 14170 23151 14172
rect 22905 14118 22907 14170
rect 23087 14118 23089 14170
rect 22843 14116 22849 14118
rect 22905 14116 22929 14118
rect 22985 14116 23009 14118
rect 23065 14116 23089 14118
rect 23145 14116 23151 14118
rect 22843 14107 23151 14116
rect 23020 13864 23072 13870
rect 23020 13806 23072 13812
rect 23032 13326 23060 13806
rect 23584 13326 23612 14214
rect 23020 13320 23072 13326
rect 23020 13262 23072 13268
rect 23572 13320 23624 13326
rect 23572 13262 23624 13268
rect 22652 13184 22704 13190
rect 22652 13126 22704 13132
rect 22468 12436 22520 12442
rect 22468 12378 22520 12384
rect 22480 11898 22508 12378
rect 22468 11892 22520 11898
rect 22468 11834 22520 11840
rect 22388 10674 22600 10690
rect 22388 10668 22612 10674
rect 22388 10662 22560 10668
rect 22560 10610 22612 10616
rect 22282 9752 22338 9761
rect 22282 9687 22338 9696
rect 22572 9110 22600 10610
rect 22560 9104 22612 9110
rect 22560 9046 22612 9052
rect 22468 8492 22520 8498
rect 22468 8434 22520 8440
rect 22192 8424 22244 8430
rect 22192 8366 22244 8372
rect 21916 8356 21968 8362
rect 21916 8298 21968 8304
rect 21928 7886 21956 8298
rect 21916 7880 21968 7886
rect 21916 7822 21968 7828
rect 21272 7744 21324 7750
rect 21272 7686 21324 7692
rect 21732 7744 21784 7750
rect 21732 7686 21784 7692
rect 20904 7268 20956 7274
rect 20904 7210 20956 7216
rect 20916 6934 20944 7210
rect 20996 6996 21048 7002
rect 20996 6938 21048 6944
rect 20444 6928 20496 6934
rect 20444 6870 20496 6876
rect 20904 6928 20956 6934
rect 20904 6870 20956 6876
rect 18604 6860 18656 6866
rect 18604 6802 18656 6808
rect 20456 6798 20484 6870
rect 18512 6792 18564 6798
rect 18512 6734 18564 6740
rect 20444 6792 20496 6798
rect 20444 6734 20496 6740
rect 18144 6724 18196 6730
rect 18144 6666 18196 6672
rect 17960 6452 18012 6458
rect 17960 6394 18012 6400
rect 17972 5846 18000 6394
rect 18156 5914 18184 6666
rect 18236 6316 18288 6322
rect 18236 6258 18288 6264
rect 18144 5908 18196 5914
rect 18144 5850 18196 5856
rect 17960 5840 18012 5846
rect 17960 5782 18012 5788
rect 18248 5778 18276 6258
rect 18328 6112 18380 6118
rect 18328 6054 18380 6060
rect 18236 5772 18288 5778
rect 18236 5714 18288 5720
rect 17960 5364 18012 5370
rect 17960 5306 18012 5312
rect 17972 5166 18000 5306
rect 18248 5234 18276 5714
rect 18340 5642 18368 6054
rect 18328 5636 18380 5642
rect 18328 5578 18380 5584
rect 18524 5545 18552 6734
rect 20720 6656 20772 6662
rect 20720 6598 20772 6604
rect 19248 6452 19300 6458
rect 19248 6394 19300 6400
rect 18604 6384 18656 6390
rect 18604 6326 18656 6332
rect 18616 5710 18644 6326
rect 19260 6322 19288 6394
rect 19156 6316 19208 6322
rect 19156 6258 19208 6264
rect 19248 6316 19300 6322
rect 19248 6258 19300 6264
rect 19340 6316 19392 6322
rect 19340 6258 19392 6264
rect 20352 6316 20404 6322
rect 20352 6258 20404 6264
rect 19168 5846 19196 6258
rect 19156 5840 19208 5846
rect 19156 5782 19208 5788
rect 18604 5704 18656 5710
rect 18604 5646 18656 5652
rect 19260 5658 19288 6258
rect 19352 5914 19380 6258
rect 19432 6248 19484 6254
rect 19432 6190 19484 6196
rect 20168 6248 20220 6254
rect 20168 6190 20220 6196
rect 19340 5908 19392 5914
rect 19340 5850 19392 5856
rect 19444 5794 19472 6190
rect 20180 5914 20208 6190
rect 20364 5914 20392 6258
rect 20628 6112 20680 6118
rect 20628 6054 20680 6060
rect 20168 5908 20220 5914
rect 20168 5850 20220 5856
rect 20352 5908 20404 5914
rect 20352 5850 20404 5856
rect 19444 5778 19564 5794
rect 19444 5772 19576 5778
rect 19444 5766 19524 5772
rect 19524 5714 19576 5720
rect 20640 5710 20668 6054
rect 20732 5710 20760 6598
rect 20812 6248 20864 6254
rect 20812 6190 20864 6196
rect 20628 5704 20680 5710
rect 19260 5642 19656 5658
rect 20628 5646 20680 5652
rect 20720 5704 20772 5710
rect 20720 5646 20772 5652
rect 19260 5636 19668 5642
rect 19260 5630 19616 5636
rect 19616 5578 19668 5584
rect 20824 5574 20852 6190
rect 20812 5568 20864 5574
rect 18510 5536 18566 5545
rect 20812 5510 20864 5516
rect 20904 5568 20956 5574
rect 20904 5510 20956 5516
rect 18510 5471 18566 5480
rect 18524 5302 18552 5471
rect 20916 5386 20944 5510
rect 20548 5370 20944 5386
rect 20536 5364 20944 5370
rect 20588 5358 20944 5364
rect 20536 5306 20588 5312
rect 18512 5296 18564 5302
rect 18512 5238 18564 5244
rect 19708 5296 19760 5302
rect 20444 5296 20496 5302
rect 19760 5256 19840 5284
rect 19708 5238 19760 5244
rect 18236 5228 18288 5234
rect 18236 5170 18288 5176
rect 17960 5160 18012 5166
rect 17958 5128 17960 5137
rect 18420 5160 18472 5166
rect 18012 5128 18014 5137
rect 18420 5102 18472 5108
rect 17958 5063 18014 5072
rect 18432 4826 18460 5102
rect 18524 5030 18552 5238
rect 18880 5228 18932 5234
rect 18880 5170 18932 5176
rect 18604 5092 18656 5098
rect 18604 5034 18656 5040
rect 18512 5024 18564 5030
rect 18512 4966 18564 4972
rect 18420 4820 18472 4826
rect 18420 4762 18472 4768
rect 18144 4684 18196 4690
rect 18144 4626 18196 4632
rect 18156 3534 18184 4626
rect 18616 4282 18644 5034
rect 18892 4826 18920 5170
rect 19812 5098 19840 5256
rect 20904 5296 20956 5302
rect 20640 5256 20904 5284
rect 20640 5250 20668 5256
rect 20496 5244 20668 5250
rect 20444 5238 20668 5244
rect 20904 5238 20956 5244
rect 20456 5222 20668 5238
rect 21008 5234 21036 6938
rect 21284 6934 21312 7686
rect 21744 7478 21772 7686
rect 21732 7472 21784 7478
rect 21732 7414 21784 7420
rect 22204 7342 22232 8366
rect 22480 8090 22508 8434
rect 22468 8084 22520 8090
rect 22468 8026 22520 8032
rect 22192 7336 22244 7342
rect 22192 7278 22244 7284
rect 21824 7268 21876 7274
rect 21824 7210 21876 7216
rect 21456 6996 21508 7002
rect 21456 6938 21508 6944
rect 21272 6928 21324 6934
rect 21272 6870 21324 6876
rect 21468 6798 21496 6938
rect 21640 6928 21692 6934
rect 21640 6870 21692 6876
rect 21652 6798 21680 6870
rect 21836 6798 21864 7210
rect 21456 6792 21508 6798
rect 21456 6734 21508 6740
rect 21640 6792 21692 6798
rect 21640 6734 21692 6740
rect 21824 6792 21876 6798
rect 21824 6734 21876 6740
rect 21732 6724 21784 6730
rect 21732 6666 21784 6672
rect 21744 6458 21772 6666
rect 22008 6656 22060 6662
rect 22008 6598 22060 6604
rect 21732 6452 21784 6458
rect 21732 6394 21784 6400
rect 22020 5778 22048 6598
rect 22560 6180 22612 6186
rect 22560 6122 22612 6128
rect 22468 6112 22520 6118
rect 22468 6054 22520 6060
rect 22008 5772 22060 5778
rect 22008 5714 22060 5720
rect 21180 5704 21232 5710
rect 21180 5646 21232 5652
rect 20996 5228 21048 5234
rect 20996 5170 21048 5176
rect 21192 5166 21220 5646
rect 22480 5574 22508 6054
rect 22468 5568 22520 5574
rect 22468 5510 22520 5516
rect 22480 5370 22508 5510
rect 22468 5364 22520 5370
rect 22468 5306 22520 5312
rect 21180 5160 21232 5166
rect 21180 5102 21232 5108
rect 19800 5092 19852 5098
rect 19800 5034 19852 5040
rect 19064 5024 19116 5030
rect 19064 4966 19116 4972
rect 20168 5024 20220 5030
rect 20168 4966 20220 4972
rect 18880 4820 18932 4826
rect 18880 4762 18932 4768
rect 18604 4276 18656 4282
rect 18604 4218 18656 4224
rect 19076 4146 19104 4966
rect 19432 4548 19484 4554
rect 19432 4490 19484 4496
rect 19064 4140 19116 4146
rect 19064 4082 19116 4088
rect 19444 3738 19472 4490
rect 20180 4282 20208 4966
rect 21192 4826 21220 5102
rect 22572 5098 22600 6122
rect 22560 5092 22612 5098
rect 22560 5034 22612 5040
rect 21364 5024 21416 5030
rect 21364 4966 21416 4972
rect 21180 4820 21232 4826
rect 21180 4762 21232 4768
rect 20720 4548 20772 4554
rect 20720 4490 20772 4496
rect 20168 4276 20220 4282
rect 20168 4218 20220 4224
rect 19800 4140 19852 4146
rect 19800 4082 19852 4088
rect 19616 3936 19668 3942
rect 19616 3878 19668 3884
rect 19432 3732 19484 3738
rect 19432 3674 19484 3680
rect 19628 3534 19656 3878
rect 18144 3528 18196 3534
rect 18144 3470 18196 3476
rect 19616 3528 19668 3534
rect 19616 3470 19668 3476
rect 18052 3460 18104 3466
rect 18052 3402 18104 3408
rect 18064 3058 18092 3402
rect 18052 3052 18104 3058
rect 18052 2994 18104 3000
rect 17132 2644 17184 2650
rect 17132 2586 17184 2592
rect 17868 2644 17920 2650
rect 17868 2586 17920 2592
rect 18156 2514 18184 3470
rect 19812 3126 19840 4082
rect 20628 3936 20680 3942
rect 20628 3878 20680 3884
rect 20640 3534 20668 3878
rect 20732 3738 20760 4490
rect 21376 4078 21404 4966
rect 21824 4616 21876 4622
rect 21824 4558 21876 4564
rect 21364 4072 21416 4078
rect 21364 4014 21416 4020
rect 21836 4010 21864 4558
rect 21824 4004 21876 4010
rect 21824 3946 21876 3952
rect 20720 3732 20772 3738
rect 20720 3674 20772 3680
rect 20628 3528 20680 3534
rect 20628 3470 20680 3476
rect 19800 3120 19852 3126
rect 19800 3062 19852 3068
rect 22664 3058 22692 13126
rect 22843 13084 23151 13093
rect 22843 13082 22849 13084
rect 22905 13082 22929 13084
rect 22985 13082 23009 13084
rect 23065 13082 23089 13084
rect 23145 13082 23151 13084
rect 22905 13030 22907 13082
rect 23087 13030 23089 13082
rect 22843 13028 22849 13030
rect 22905 13028 22929 13030
rect 22985 13028 23009 13030
rect 23065 13028 23089 13030
rect 23145 13028 23151 13030
rect 22843 13019 23151 13028
rect 22744 12844 22796 12850
rect 22744 12786 22796 12792
rect 22756 12442 22784 12786
rect 22744 12436 22796 12442
rect 22744 12378 22796 12384
rect 22843 11996 23151 12005
rect 22843 11994 22849 11996
rect 22905 11994 22929 11996
rect 22985 11994 23009 11996
rect 23065 11994 23089 11996
rect 23145 11994 23151 11996
rect 22905 11942 22907 11994
rect 23087 11942 23089 11994
rect 22843 11940 22849 11942
rect 22905 11940 22929 11942
rect 22985 11940 23009 11942
rect 23065 11940 23089 11942
rect 23145 11940 23151 11942
rect 22843 11931 23151 11940
rect 22744 11688 22796 11694
rect 22744 11630 22796 11636
rect 22756 10198 22784 11630
rect 23388 11552 23440 11558
rect 23388 11494 23440 11500
rect 23400 11150 23428 11494
rect 23388 11144 23440 11150
rect 23388 11086 23440 11092
rect 22843 10908 23151 10917
rect 22843 10906 22849 10908
rect 22905 10906 22929 10908
rect 22985 10906 23009 10908
rect 23065 10906 23089 10908
rect 23145 10906 23151 10908
rect 22905 10854 22907 10906
rect 23087 10854 23089 10906
rect 22843 10852 22849 10854
rect 22905 10852 22929 10854
rect 22985 10852 23009 10854
rect 23065 10852 23089 10854
rect 23145 10852 23151 10854
rect 22843 10843 23151 10852
rect 23204 10736 23256 10742
rect 23204 10678 23256 10684
rect 22744 10192 22796 10198
rect 22744 10134 22796 10140
rect 23216 10062 23244 10678
rect 23676 10577 23704 14282
rect 23860 13938 23888 14418
rect 24412 14414 24440 14758
rect 24400 14408 24452 14414
rect 24400 14350 24452 14356
rect 23848 13932 23900 13938
rect 23848 13874 23900 13880
rect 23860 12434 23888 13874
rect 24872 13870 24900 14962
rect 25240 14618 25268 15438
rect 27712 15020 27764 15026
rect 27712 14962 27764 14968
rect 30196 15020 30248 15026
rect 30196 14962 30248 14968
rect 26608 14816 26660 14822
rect 26608 14758 26660 14764
rect 25228 14612 25280 14618
rect 25228 14554 25280 14560
rect 25504 14476 25556 14482
rect 25504 14418 25556 14424
rect 25516 14006 25544 14418
rect 26620 14414 26648 14758
rect 26792 14476 26844 14482
rect 26792 14418 26844 14424
rect 26608 14408 26660 14414
rect 26608 14350 26660 14356
rect 26620 14074 26648 14350
rect 26804 14278 26832 14418
rect 26792 14272 26844 14278
rect 26792 14214 26844 14220
rect 26608 14068 26660 14074
rect 26608 14010 26660 14016
rect 25504 14000 25556 14006
rect 25504 13942 25556 13948
rect 24860 13864 24912 13870
rect 24860 13806 24912 13812
rect 24676 13388 24728 13394
rect 24676 13330 24728 13336
rect 24584 12844 24636 12850
rect 24584 12786 24636 12792
rect 24596 12442 24624 12786
rect 24584 12436 24636 12442
rect 23860 12406 23980 12434
rect 23848 12300 23900 12306
rect 23848 12242 23900 12248
rect 23860 11830 23888 12242
rect 23848 11824 23900 11830
rect 23848 11766 23900 11772
rect 23662 10568 23718 10577
rect 23662 10503 23718 10512
rect 23664 10464 23716 10470
rect 23664 10406 23716 10412
rect 23204 10056 23256 10062
rect 23204 9998 23256 10004
rect 22843 9820 23151 9829
rect 22843 9818 22849 9820
rect 22905 9818 22929 9820
rect 22985 9818 23009 9820
rect 23065 9818 23089 9820
rect 23145 9818 23151 9820
rect 22905 9766 22907 9818
rect 23087 9766 23089 9818
rect 22843 9764 22849 9766
rect 22905 9764 22929 9766
rect 22985 9764 23009 9766
rect 23065 9764 23089 9766
rect 23145 9764 23151 9766
rect 22843 9755 23151 9764
rect 23216 8838 23244 9998
rect 23480 9920 23532 9926
rect 23480 9862 23532 9868
rect 23296 9580 23348 9586
rect 23296 9522 23348 9528
rect 23204 8832 23256 8838
rect 23204 8774 23256 8780
rect 22843 8732 23151 8741
rect 22843 8730 22849 8732
rect 22905 8730 22929 8732
rect 22985 8730 23009 8732
rect 23065 8730 23089 8732
rect 23145 8730 23151 8732
rect 22905 8678 22907 8730
rect 23087 8678 23089 8730
rect 22843 8676 22849 8678
rect 22905 8676 22929 8678
rect 22985 8676 23009 8678
rect 23065 8676 23089 8678
rect 23145 8676 23151 8678
rect 22843 8667 23151 8676
rect 22843 7644 23151 7653
rect 22843 7642 22849 7644
rect 22905 7642 22929 7644
rect 22985 7642 23009 7644
rect 23065 7642 23089 7644
rect 23145 7642 23151 7644
rect 22905 7590 22907 7642
rect 23087 7590 23089 7642
rect 22843 7588 22849 7590
rect 22905 7588 22929 7590
rect 22985 7588 23009 7590
rect 23065 7588 23089 7590
rect 23145 7588 23151 7590
rect 22843 7579 23151 7588
rect 22843 6556 23151 6565
rect 22843 6554 22849 6556
rect 22905 6554 22929 6556
rect 22985 6554 23009 6556
rect 23065 6554 23089 6556
rect 23145 6554 23151 6556
rect 22905 6502 22907 6554
rect 23087 6502 23089 6554
rect 22843 6500 22849 6502
rect 22905 6500 22929 6502
rect 22985 6500 23009 6502
rect 23065 6500 23089 6502
rect 23145 6500 23151 6502
rect 22843 6491 23151 6500
rect 22744 6316 22796 6322
rect 22744 6258 22796 6264
rect 23112 6316 23164 6322
rect 23112 6258 23164 6264
rect 22756 5370 22784 6258
rect 23020 6180 23072 6186
rect 23020 6122 23072 6128
rect 23032 5914 23060 6122
rect 23124 5914 23152 6258
rect 23020 5908 23072 5914
rect 23020 5850 23072 5856
rect 23112 5908 23164 5914
rect 23112 5850 23164 5856
rect 22843 5468 23151 5477
rect 22843 5466 22849 5468
rect 22905 5466 22929 5468
rect 22985 5466 23009 5468
rect 23065 5466 23089 5468
rect 23145 5466 23151 5468
rect 22905 5414 22907 5466
rect 23087 5414 23089 5466
rect 22843 5412 22849 5414
rect 22905 5412 22929 5414
rect 22985 5412 23009 5414
rect 23065 5412 23089 5414
rect 23145 5412 23151 5414
rect 22843 5403 23151 5412
rect 22744 5364 22796 5370
rect 22744 5306 22796 5312
rect 22843 4380 23151 4389
rect 22843 4378 22849 4380
rect 22905 4378 22929 4380
rect 22985 4378 23009 4380
rect 23065 4378 23089 4380
rect 23145 4378 23151 4380
rect 22905 4326 22907 4378
rect 23087 4326 23089 4378
rect 22843 4324 22849 4326
rect 22905 4324 22929 4326
rect 22985 4324 23009 4326
rect 23065 4324 23089 4326
rect 23145 4324 23151 4326
rect 22843 4315 23151 4324
rect 23308 3466 23336 9522
rect 23492 9178 23520 9862
rect 23480 9172 23532 9178
rect 23480 9114 23532 9120
rect 23676 9042 23704 10406
rect 23848 9648 23900 9654
rect 23846 9616 23848 9625
rect 23900 9616 23902 9625
rect 23846 9551 23902 9560
rect 23756 9172 23808 9178
rect 23756 9114 23808 9120
rect 23664 9036 23716 9042
rect 23664 8978 23716 8984
rect 23480 8832 23532 8838
rect 23480 8774 23532 8780
rect 23388 7880 23440 7886
rect 23492 7868 23520 8774
rect 23440 7840 23520 7868
rect 23572 7880 23624 7886
rect 23388 7822 23440 7828
rect 23572 7822 23624 7828
rect 23388 7744 23440 7750
rect 23388 7686 23440 7692
rect 23400 7478 23428 7686
rect 23388 7472 23440 7478
rect 23388 7414 23440 7420
rect 23388 7200 23440 7206
rect 23440 7148 23520 7154
rect 23388 7142 23520 7148
rect 23400 7126 23520 7142
rect 23492 6254 23520 7126
rect 23584 6662 23612 7822
rect 23768 6866 23796 9114
rect 23848 8356 23900 8362
rect 23848 8298 23900 8304
rect 23860 6866 23888 8298
rect 23756 6860 23808 6866
rect 23756 6802 23808 6808
rect 23848 6860 23900 6866
rect 23848 6802 23900 6808
rect 23572 6656 23624 6662
rect 23572 6598 23624 6604
rect 23756 6384 23808 6390
rect 23756 6326 23808 6332
rect 23480 6248 23532 6254
rect 23480 6190 23532 6196
rect 23388 5840 23440 5846
rect 23388 5782 23440 5788
rect 23400 5302 23428 5782
rect 23388 5296 23440 5302
rect 23388 5238 23440 5244
rect 23768 4826 23796 6326
rect 23952 5817 23980 12406
rect 24584 12378 24636 12384
rect 24688 10418 24716 13330
rect 24872 13326 24900 13806
rect 25516 13530 25544 13942
rect 26148 13864 26200 13870
rect 26148 13806 26200 13812
rect 25504 13524 25556 13530
rect 25504 13466 25556 13472
rect 24860 13320 24912 13326
rect 24860 13262 24912 13268
rect 24872 12986 24900 13262
rect 24860 12980 24912 12986
rect 24860 12922 24912 12928
rect 24872 11218 24900 12922
rect 24952 12640 25004 12646
rect 24952 12582 25004 12588
rect 24964 12102 24992 12582
rect 26160 12306 26188 13806
rect 26804 13802 26832 14214
rect 26792 13796 26844 13802
rect 26792 13738 26844 13744
rect 27160 12844 27212 12850
rect 27160 12786 27212 12792
rect 26884 12640 26936 12646
rect 26884 12582 26936 12588
rect 26148 12300 26200 12306
rect 26148 12242 26200 12248
rect 25228 12232 25280 12238
rect 25228 12174 25280 12180
rect 24952 12096 25004 12102
rect 24952 12038 25004 12044
rect 24964 11830 24992 12038
rect 24952 11824 25004 11830
rect 24952 11766 25004 11772
rect 24860 11212 24912 11218
rect 24860 11154 24912 11160
rect 25240 10674 25268 12174
rect 26896 12170 26924 12582
rect 26424 12164 26476 12170
rect 26424 12106 26476 12112
rect 26884 12164 26936 12170
rect 26884 12106 26936 12112
rect 26436 11898 26464 12106
rect 26424 11892 26476 11898
rect 26424 11834 26476 11840
rect 25596 11620 25648 11626
rect 25596 11562 25648 11568
rect 25608 11354 25636 11562
rect 27172 11558 27200 12786
rect 27436 12300 27488 12306
rect 27436 12242 27488 12248
rect 27448 11762 27476 12242
rect 27436 11756 27488 11762
rect 27436 11698 27488 11704
rect 27620 11756 27672 11762
rect 27620 11698 27672 11704
rect 27632 11626 27660 11698
rect 27620 11620 27672 11626
rect 27620 11562 27672 11568
rect 27160 11552 27212 11558
rect 27160 11494 27212 11500
rect 25596 11348 25648 11354
rect 25596 11290 25648 11296
rect 25608 10810 25636 11290
rect 27172 11286 27200 11494
rect 27160 11280 27212 11286
rect 27160 11222 27212 11228
rect 26792 11212 26844 11218
rect 26792 11154 26844 11160
rect 26884 11212 26936 11218
rect 26884 11154 26936 11160
rect 26424 11076 26476 11082
rect 26424 11018 26476 11024
rect 25596 10804 25648 10810
rect 25596 10746 25648 10752
rect 25228 10668 25280 10674
rect 25228 10610 25280 10616
rect 26056 10668 26108 10674
rect 26056 10610 26108 10616
rect 24688 10390 24900 10418
rect 24766 10024 24822 10033
rect 24872 10010 24900 10390
rect 24822 9982 24900 10010
rect 24766 9959 24822 9968
rect 24492 8968 24544 8974
rect 24492 8910 24544 8916
rect 24400 7200 24452 7206
rect 24400 7142 24452 7148
rect 24412 6798 24440 7142
rect 24400 6792 24452 6798
rect 24400 6734 24452 6740
rect 24504 6254 24532 8910
rect 24872 8906 24900 9982
rect 25228 9580 25280 9586
rect 25228 9522 25280 9528
rect 24860 8900 24912 8906
rect 24860 8842 24912 8848
rect 25136 8832 25188 8838
rect 25136 8774 25188 8780
rect 25148 8634 25176 8774
rect 25240 8634 25268 9522
rect 25320 9376 25372 9382
rect 25320 9318 25372 9324
rect 25332 8906 25360 9318
rect 25320 8900 25372 8906
rect 25320 8842 25372 8848
rect 25136 8628 25188 8634
rect 25136 8570 25188 8576
rect 25228 8628 25280 8634
rect 25228 8570 25280 8576
rect 26068 8566 26096 10610
rect 26332 10464 26384 10470
rect 26332 10406 26384 10412
rect 26344 10062 26372 10406
rect 26436 10266 26464 11018
rect 26700 11008 26752 11014
rect 26700 10950 26752 10956
rect 26712 10810 26740 10950
rect 26700 10804 26752 10810
rect 26700 10746 26752 10752
rect 26804 10266 26832 11154
rect 26896 10742 26924 11154
rect 27632 11150 27660 11562
rect 27620 11144 27672 11150
rect 27620 11086 27672 11092
rect 27436 11076 27488 11082
rect 27436 11018 27488 11024
rect 26884 10736 26936 10742
rect 27448 10690 27476 11018
rect 27620 11008 27672 11014
rect 27620 10950 27672 10956
rect 26884 10678 26936 10684
rect 27356 10662 27476 10690
rect 27160 10600 27212 10606
rect 27160 10542 27212 10548
rect 26424 10260 26476 10266
rect 26424 10202 26476 10208
rect 26792 10260 26844 10266
rect 26792 10202 26844 10208
rect 26332 10056 26384 10062
rect 26332 9998 26384 10004
rect 26332 9580 26384 9586
rect 26332 9522 26384 9528
rect 26344 9178 26372 9522
rect 27068 9376 27120 9382
rect 27068 9318 27120 9324
rect 26332 9172 26384 9178
rect 26332 9114 26384 9120
rect 27080 8974 27108 9318
rect 27068 8968 27120 8974
rect 27068 8910 27120 8916
rect 26240 8832 26292 8838
rect 26240 8774 26292 8780
rect 26056 8560 26108 8566
rect 26056 8502 26108 8508
rect 25964 8492 26016 8498
rect 25964 8434 26016 8440
rect 25976 7410 26004 8434
rect 26252 7970 26280 8774
rect 26160 7954 26280 7970
rect 26148 7948 26280 7954
rect 26200 7942 26280 7948
rect 26148 7890 26200 7896
rect 25964 7404 26016 7410
rect 25964 7346 26016 7352
rect 25044 6792 25096 6798
rect 25044 6734 25096 6740
rect 24584 6384 24636 6390
rect 24584 6326 24636 6332
rect 24492 6248 24544 6254
rect 24492 6190 24544 6196
rect 24124 6112 24176 6118
rect 24124 6054 24176 6060
rect 23938 5808 23994 5817
rect 23938 5743 23994 5752
rect 24136 5710 24164 6054
rect 24124 5704 24176 5710
rect 24124 5646 24176 5652
rect 24308 5568 24360 5574
rect 24308 5510 24360 5516
rect 24032 5364 24084 5370
rect 24032 5306 24084 5312
rect 23940 5228 23992 5234
rect 23940 5170 23992 5176
rect 23952 5030 23980 5170
rect 23940 5024 23992 5030
rect 23940 4966 23992 4972
rect 23756 4820 23808 4826
rect 23756 4762 23808 4768
rect 23664 4684 23716 4690
rect 23664 4626 23716 4632
rect 23676 4146 23704 4626
rect 23768 4282 23796 4762
rect 23952 4758 23980 4966
rect 23940 4752 23992 4758
rect 23940 4694 23992 4700
rect 24044 4622 24072 5306
rect 24320 5234 24348 5510
rect 24308 5228 24360 5234
rect 24308 5170 24360 5176
rect 24504 4690 24532 6190
rect 24596 5914 24624 6326
rect 24860 6112 24912 6118
rect 24860 6054 24912 6060
rect 24584 5908 24636 5914
rect 24584 5850 24636 5856
rect 24872 5710 24900 6054
rect 25056 5710 25084 6734
rect 25872 6656 25924 6662
rect 25872 6598 25924 6604
rect 25884 6390 25912 6598
rect 25872 6384 25924 6390
rect 25872 6326 25924 6332
rect 24860 5704 24912 5710
rect 24860 5646 24912 5652
rect 25044 5704 25096 5710
rect 25872 5704 25924 5710
rect 25044 5646 25096 5652
rect 25870 5672 25872 5681
rect 25924 5672 25926 5681
rect 25870 5607 25926 5616
rect 25228 5568 25280 5574
rect 25228 5510 25280 5516
rect 25240 5234 25268 5510
rect 25228 5228 25280 5234
rect 25228 5170 25280 5176
rect 25320 5228 25372 5234
rect 25320 5170 25372 5176
rect 25332 4826 25360 5170
rect 25872 5024 25924 5030
rect 25872 4966 25924 4972
rect 24584 4820 24636 4826
rect 24584 4762 24636 4768
rect 25320 4820 25372 4826
rect 25320 4762 25372 4768
rect 24492 4684 24544 4690
rect 24492 4626 24544 4632
rect 24596 4622 24624 4762
rect 24032 4616 24084 4622
rect 24584 4616 24636 4622
rect 24084 4576 24164 4604
rect 24032 4558 24084 4564
rect 24136 4486 24164 4576
rect 24584 4558 24636 4564
rect 25884 4554 25912 4966
rect 25872 4548 25924 4554
rect 25872 4490 25924 4496
rect 24032 4480 24084 4486
rect 24032 4422 24084 4428
rect 24124 4480 24176 4486
rect 24124 4422 24176 4428
rect 25412 4480 25464 4486
rect 25412 4422 25464 4428
rect 23756 4276 23808 4282
rect 23756 4218 23808 4224
rect 23664 4140 23716 4146
rect 23664 4082 23716 4088
rect 23940 4072 23992 4078
rect 23940 4014 23992 4020
rect 23952 3738 23980 4014
rect 23940 3732 23992 3738
rect 23940 3674 23992 3680
rect 24044 3534 24072 4422
rect 25424 4282 25452 4422
rect 25412 4276 25464 4282
rect 25412 4218 25464 4224
rect 25976 4078 26004 7346
rect 26240 7336 26292 7342
rect 26240 7278 26292 7284
rect 26056 6792 26108 6798
rect 26056 6734 26108 6740
rect 26068 5914 26096 6734
rect 26056 5908 26108 5914
rect 26056 5850 26108 5856
rect 26252 5710 26280 7278
rect 27080 6322 27108 8910
rect 27172 8362 27200 10542
rect 27356 9586 27384 10662
rect 27436 10600 27488 10606
rect 27436 10542 27488 10548
rect 27448 9722 27476 10542
rect 27632 10130 27660 10950
rect 27620 10124 27672 10130
rect 27620 10066 27672 10072
rect 27436 9716 27488 9722
rect 27436 9658 27488 9664
rect 27344 9580 27396 9586
rect 27344 9522 27396 9528
rect 27724 9450 27752 14962
rect 29552 14952 29604 14958
rect 29552 14894 29604 14900
rect 28908 14816 28960 14822
rect 28908 14758 28960 14764
rect 28317 14716 28625 14725
rect 28317 14714 28323 14716
rect 28379 14714 28403 14716
rect 28459 14714 28483 14716
rect 28539 14714 28563 14716
rect 28619 14714 28625 14716
rect 28379 14662 28381 14714
rect 28561 14662 28563 14714
rect 28317 14660 28323 14662
rect 28379 14660 28403 14662
rect 28459 14660 28483 14662
rect 28539 14660 28563 14662
rect 28619 14660 28625 14662
rect 28317 14651 28625 14660
rect 28920 14414 28948 14758
rect 27804 14408 27856 14414
rect 27804 14350 27856 14356
rect 28908 14408 28960 14414
rect 28908 14350 28960 14356
rect 27816 13870 27844 14350
rect 27804 13864 27856 13870
rect 27804 13806 27856 13812
rect 28317 13628 28625 13637
rect 28317 13626 28323 13628
rect 28379 13626 28403 13628
rect 28459 13626 28483 13628
rect 28539 13626 28563 13628
rect 28619 13626 28625 13628
rect 28379 13574 28381 13626
rect 28561 13574 28563 13626
rect 28317 13572 28323 13574
rect 28379 13572 28403 13574
rect 28459 13572 28483 13574
rect 28539 13572 28563 13574
rect 28619 13572 28625 13574
rect 28317 13563 28625 13572
rect 28920 13326 28948 14350
rect 29564 13938 29592 14894
rect 29644 14884 29696 14890
rect 29644 14826 29696 14832
rect 29656 14618 29684 14826
rect 30012 14816 30064 14822
rect 30012 14758 30064 14764
rect 29644 14612 29696 14618
rect 29644 14554 29696 14560
rect 29736 14408 29788 14414
rect 29736 14350 29788 14356
rect 29552 13932 29604 13938
rect 29552 13874 29604 13880
rect 29748 13870 29776 14350
rect 30024 13938 30052 14758
rect 30208 14074 30236 14962
rect 31116 14816 31168 14822
rect 31116 14758 31168 14764
rect 31208 14816 31260 14822
rect 31208 14758 31260 14764
rect 31128 14414 31156 14758
rect 30932 14408 30984 14414
rect 30932 14350 30984 14356
rect 31116 14408 31168 14414
rect 31116 14350 31168 14356
rect 30196 14068 30248 14074
rect 30196 14010 30248 14016
rect 30012 13932 30064 13938
rect 30012 13874 30064 13880
rect 30288 13932 30340 13938
rect 30288 13874 30340 13880
rect 29000 13864 29052 13870
rect 29000 13806 29052 13812
rect 29736 13864 29788 13870
rect 29736 13806 29788 13812
rect 27896 13320 27948 13326
rect 27896 13262 27948 13268
rect 28172 13320 28224 13326
rect 28172 13262 28224 13268
rect 28908 13320 28960 13326
rect 28908 13262 28960 13268
rect 27908 12442 27936 13262
rect 28080 13184 28132 13190
rect 28080 13126 28132 13132
rect 28092 12646 28120 13126
rect 28080 12640 28132 12646
rect 28080 12582 28132 12588
rect 28092 12442 28120 12582
rect 27896 12436 27948 12442
rect 27896 12378 27948 12384
rect 28080 12436 28132 12442
rect 28080 12378 28132 12384
rect 28184 11694 28212 13262
rect 28264 13184 28316 13190
rect 28264 13126 28316 13132
rect 28276 12918 28304 13126
rect 28920 12986 28948 13262
rect 28908 12980 28960 12986
rect 28908 12922 28960 12928
rect 28264 12912 28316 12918
rect 28264 12854 28316 12860
rect 28317 12540 28625 12549
rect 28317 12538 28323 12540
rect 28379 12538 28403 12540
rect 28459 12538 28483 12540
rect 28539 12538 28563 12540
rect 28619 12538 28625 12540
rect 28379 12486 28381 12538
rect 28561 12486 28563 12538
rect 28317 12484 28323 12486
rect 28379 12484 28403 12486
rect 28459 12484 28483 12486
rect 28539 12484 28563 12486
rect 28619 12484 28625 12486
rect 28317 12475 28625 12484
rect 28264 12436 28316 12442
rect 28264 12378 28316 12384
rect 28724 12436 28776 12442
rect 29012 12434 29040 13806
rect 30300 12442 30328 13874
rect 30840 13320 30892 13326
rect 30944 13308 30972 14350
rect 31116 14272 31168 14278
rect 31116 14214 31168 14220
rect 30892 13280 30972 13308
rect 30840 13262 30892 13268
rect 30380 12844 30432 12850
rect 30380 12786 30432 12792
rect 30288 12436 30340 12442
rect 29012 12406 29132 12434
rect 28724 12378 28776 12384
rect 28276 12220 28304 12378
rect 28356 12368 28408 12374
rect 28540 12368 28592 12374
rect 28408 12316 28540 12322
rect 28356 12310 28592 12316
rect 28368 12294 28580 12310
rect 28540 12232 28592 12238
rect 28276 12192 28540 12220
rect 28540 12174 28592 12180
rect 28632 12232 28684 12238
rect 28632 12174 28684 12180
rect 28644 12102 28672 12174
rect 28632 12096 28684 12102
rect 28632 12038 28684 12044
rect 28172 11688 28224 11694
rect 28172 11630 28224 11636
rect 28317 11452 28625 11461
rect 28317 11450 28323 11452
rect 28379 11450 28403 11452
rect 28459 11450 28483 11452
rect 28539 11450 28563 11452
rect 28619 11450 28625 11452
rect 28379 11398 28381 11450
rect 28561 11398 28563 11450
rect 28317 11396 28323 11398
rect 28379 11396 28403 11398
rect 28459 11396 28483 11398
rect 28539 11396 28563 11398
rect 28619 11396 28625 11398
rect 28317 11387 28625 11396
rect 28736 11286 28764 12378
rect 28908 12164 28960 12170
rect 28908 12106 28960 12112
rect 28920 11694 28948 12106
rect 29000 11756 29052 11762
rect 29000 11698 29052 11704
rect 28908 11688 28960 11694
rect 28908 11630 28960 11636
rect 27896 11280 27948 11286
rect 28724 11280 28776 11286
rect 27896 11222 27948 11228
rect 28552 11228 28724 11234
rect 28552 11222 28776 11228
rect 27908 11121 27936 11222
rect 28552 11218 28764 11222
rect 28540 11212 28764 11218
rect 28592 11206 28764 11212
rect 28540 11154 28592 11160
rect 28920 11150 28948 11630
rect 28908 11144 28960 11150
rect 27894 11112 27950 11121
rect 28908 11086 28960 11092
rect 27894 11047 27950 11056
rect 27908 10130 27936 11047
rect 28172 10736 28224 10742
rect 28078 10704 28134 10713
rect 28172 10678 28224 10684
rect 28078 10639 28134 10648
rect 27896 10124 27948 10130
rect 27896 10066 27948 10072
rect 27894 9616 27950 9625
rect 28092 9586 28120 10639
rect 28184 10266 28212 10678
rect 29012 10470 29040 11698
rect 29104 10713 29132 12406
rect 30288 12378 30340 12384
rect 30392 11830 30420 12786
rect 30564 12300 30616 12306
rect 30564 12242 30616 12248
rect 30472 12232 30524 12238
rect 30472 12174 30524 12180
rect 30380 11824 30432 11830
rect 30380 11766 30432 11772
rect 30484 11626 30512 12174
rect 30472 11620 30524 11626
rect 30472 11562 30524 11568
rect 30576 11354 30604 12242
rect 30944 12238 30972 13280
rect 31024 12640 31076 12646
rect 31024 12582 31076 12588
rect 30932 12232 30984 12238
rect 31036 12209 31064 12582
rect 30932 12174 30984 12180
rect 31022 12200 31078 12209
rect 30656 11756 30708 11762
rect 30656 11698 30708 11704
rect 30840 11756 30892 11762
rect 30840 11698 30892 11704
rect 30380 11348 30432 11354
rect 30380 11290 30432 11296
rect 30564 11348 30616 11354
rect 30564 11290 30616 11296
rect 30288 11008 30340 11014
rect 30288 10950 30340 10956
rect 29090 10704 29146 10713
rect 29090 10639 29146 10648
rect 29644 10668 29696 10674
rect 29644 10610 29696 10616
rect 29092 10600 29144 10606
rect 29092 10542 29144 10548
rect 29000 10464 29052 10470
rect 29000 10406 29052 10412
rect 28317 10364 28625 10373
rect 28317 10362 28323 10364
rect 28379 10362 28403 10364
rect 28459 10362 28483 10364
rect 28539 10362 28563 10364
rect 28619 10362 28625 10364
rect 28379 10310 28381 10362
rect 28561 10310 28563 10362
rect 28317 10308 28323 10310
rect 28379 10308 28403 10310
rect 28459 10308 28483 10310
rect 28539 10308 28563 10310
rect 28619 10308 28625 10310
rect 28317 10299 28625 10308
rect 28172 10260 28224 10266
rect 28172 10202 28224 10208
rect 28172 10124 28224 10130
rect 28172 10066 28224 10072
rect 27894 9551 27950 9560
rect 27988 9580 28040 9586
rect 27712 9444 27764 9450
rect 27712 9386 27764 9392
rect 27908 9382 27936 9551
rect 27988 9522 28040 9528
rect 28080 9580 28132 9586
rect 28080 9522 28132 9528
rect 27804 9376 27856 9382
rect 27804 9318 27856 9324
rect 27896 9376 27948 9382
rect 27896 9318 27948 9324
rect 27528 8968 27580 8974
rect 27528 8910 27580 8916
rect 27436 8560 27488 8566
rect 27436 8502 27488 8508
rect 27160 8356 27212 8362
rect 27160 8298 27212 8304
rect 27172 7954 27200 8298
rect 27160 7948 27212 7954
rect 27160 7890 27212 7896
rect 27172 7342 27200 7890
rect 27448 7886 27476 8502
rect 27540 8362 27568 8910
rect 27528 8356 27580 8362
rect 27528 8298 27580 8304
rect 27436 7880 27488 7886
rect 27436 7822 27488 7828
rect 27816 7818 27844 9318
rect 27896 8832 27948 8838
rect 27896 8774 27948 8780
rect 27908 7954 27936 8774
rect 28000 8090 28028 9522
rect 28080 9172 28132 9178
rect 28080 9114 28132 9120
rect 28092 8906 28120 9114
rect 28080 8900 28132 8906
rect 28080 8842 28132 8848
rect 28184 8566 28212 10066
rect 29000 10056 29052 10062
rect 29000 9998 29052 10004
rect 29012 9518 29040 9998
rect 29000 9512 29052 9518
rect 29000 9454 29052 9460
rect 28317 9276 28625 9285
rect 28317 9274 28323 9276
rect 28379 9274 28403 9276
rect 28459 9274 28483 9276
rect 28539 9274 28563 9276
rect 28619 9274 28625 9276
rect 28379 9222 28381 9274
rect 28561 9222 28563 9274
rect 28317 9220 28323 9222
rect 28379 9220 28403 9222
rect 28459 9220 28483 9222
rect 28539 9220 28563 9222
rect 28619 9220 28625 9222
rect 28317 9211 28625 9220
rect 29104 8838 29132 10542
rect 29552 9920 29604 9926
rect 29552 9862 29604 9868
rect 29564 9586 29592 9862
rect 29656 9654 29684 10610
rect 30300 9994 30328 10950
rect 30392 10062 30420 11290
rect 30472 11144 30524 11150
rect 30472 11086 30524 11092
rect 30484 10198 30512 11086
rect 30668 11082 30696 11698
rect 30656 11076 30708 11082
rect 30656 11018 30708 11024
rect 30852 10266 30880 11698
rect 30944 11150 30972 12174
rect 31022 12135 31078 12144
rect 31024 11756 31076 11762
rect 31024 11698 31076 11704
rect 31036 11558 31064 11698
rect 31024 11552 31076 11558
rect 31024 11494 31076 11500
rect 30932 11144 30984 11150
rect 30932 11086 30984 11092
rect 30944 10810 30972 11086
rect 30932 10804 30984 10810
rect 30932 10746 30984 10752
rect 30840 10260 30892 10266
rect 30840 10202 30892 10208
rect 30472 10192 30524 10198
rect 30472 10134 30524 10140
rect 30380 10056 30432 10062
rect 30380 9998 30432 10004
rect 31128 9994 31156 14214
rect 31220 14006 31248 14758
rect 31208 14000 31260 14006
rect 31208 13942 31260 13948
rect 31208 12844 31260 12850
rect 31208 12786 31260 12792
rect 31220 11762 31248 12786
rect 31208 11756 31260 11762
rect 31208 11698 31260 11704
rect 31312 10690 31340 16934
rect 32600 15162 32628 17070
rect 34520 16992 34572 16998
rect 34520 16934 34572 16940
rect 38844 16992 38896 16998
rect 38844 16934 38896 16940
rect 33790 16348 34098 16357
rect 33790 16346 33796 16348
rect 33852 16346 33876 16348
rect 33932 16346 33956 16348
rect 34012 16346 34036 16348
rect 34092 16346 34098 16348
rect 33852 16294 33854 16346
rect 34034 16294 34036 16346
rect 33790 16292 33796 16294
rect 33852 16292 33876 16294
rect 33932 16292 33956 16294
rect 34012 16292 34036 16294
rect 34092 16292 34098 16294
rect 33790 16283 34098 16292
rect 33790 15260 34098 15269
rect 33790 15258 33796 15260
rect 33852 15258 33876 15260
rect 33932 15258 33956 15260
rect 34012 15258 34036 15260
rect 34092 15258 34098 15260
rect 33852 15206 33854 15258
rect 34034 15206 34036 15258
rect 33790 15204 33796 15206
rect 33852 15204 33876 15206
rect 33932 15204 33956 15206
rect 34012 15204 34036 15206
rect 34092 15204 34098 15206
rect 33790 15195 34098 15204
rect 32588 15156 32640 15162
rect 32588 15098 32640 15104
rect 32036 15088 32088 15094
rect 32036 15030 32088 15036
rect 31392 15020 31444 15026
rect 31392 14962 31444 14968
rect 31404 14618 31432 14962
rect 31392 14612 31444 14618
rect 31392 14554 31444 14560
rect 31392 14068 31444 14074
rect 31392 14010 31444 14016
rect 31404 12170 31432 14010
rect 31484 13184 31536 13190
rect 31484 13126 31536 13132
rect 31496 12986 31524 13126
rect 31484 12980 31536 12986
rect 31484 12922 31536 12928
rect 32048 12918 32076 15030
rect 33600 15020 33652 15026
rect 33600 14962 33652 14968
rect 33612 14618 33640 14962
rect 34532 14958 34560 16934
rect 35716 16040 35768 16046
rect 36176 16040 36228 16046
rect 35716 15982 35768 15988
rect 36096 16000 36176 16028
rect 35728 15706 35756 15982
rect 35716 15700 35768 15706
rect 35716 15642 35768 15648
rect 35900 15564 35952 15570
rect 35900 15506 35952 15512
rect 34520 14952 34572 14958
rect 34520 14894 34572 14900
rect 34612 14952 34664 14958
rect 34612 14894 34664 14900
rect 33600 14612 33652 14618
rect 33600 14554 33652 14560
rect 34624 14414 34652 14894
rect 35912 14482 35940 15506
rect 35900 14476 35952 14482
rect 35900 14418 35952 14424
rect 32404 14408 32456 14414
rect 32404 14350 32456 14356
rect 34612 14408 34664 14414
rect 34612 14350 34664 14356
rect 32416 13870 32444 14350
rect 33790 14172 34098 14181
rect 33790 14170 33796 14172
rect 33852 14170 33876 14172
rect 33932 14170 33956 14172
rect 34012 14170 34036 14172
rect 34092 14170 34098 14172
rect 33852 14118 33854 14170
rect 34034 14118 34036 14170
rect 33790 14116 33796 14118
rect 33852 14116 33876 14118
rect 33932 14116 33956 14118
rect 34012 14116 34036 14118
rect 34092 14116 34098 14118
rect 33790 14107 34098 14116
rect 34624 14006 34652 14350
rect 34612 14000 34664 14006
rect 34612 13942 34664 13948
rect 32404 13864 32456 13870
rect 32404 13806 32456 13812
rect 32772 13320 32824 13326
rect 32772 13262 32824 13268
rect 32036 12912 32088 12918
rect 32036 12854 32088 12860
rect 31484 12776 31536 12782
rect 31484 12718 31536 12724
rect 32312 12776 32364 12782
rect 32312 12718 32364 12724
rect 31496 12646 31524 12718
rect 31484 12640 31536 12646
rect 31484 12582 31536 12588
rect 31392 12164 31444 12170
rect 31392 12106 31444 12112
rect 31496 10742 31524 12582
rect 31852 12300 31904 12306
rect 31852 12242 31904 12248
rect 31576 11348 31628 11354
rect 31576 11290 31628 11296
rect 31484 10736 31536 10742
rect 31312 10662 31432 10690
rect 31484 10678 31536 10684
rect 31300 10056 31352 10062
rect 31300 9998 31352 10004
rect 30288 9988 30340 9994
rect 30288 9930 30340 9936
rect 31116 9988 31168 9994
rect 31116 9930 31168 9936
rect 31312 9722 31340 9998
rect 31300 9716 31352 9722
rect 31300 9658 31352 9664
rect 29644 9648 29696 9654
rect 29644 9590 29696 9596
rect 29184 9580 29236 9586
rect 29184 9522 29236 9528
rect 29552 9580 29604 9586
rect 29552 9522 29604 9528
rect 29196 9178 29224 9522
rect 29276 9512 29328 9518
rect 29276 9454 29328 9460
rect 29184 9172 29236 9178
rect 29184 9114 29236 9120
rect 29092 8832 29144 8838
rect 29092 8774 29144 8780
rect 28172 8560 28224 8566
rect 28172 8502 28224 8508
rect 29288 8362 29316 9454
rect 29656 8498 29684 9590
rect 31116 9580 31168 9586
rect 31116 9522 31168 9528
rect 31300 9580 31352 9586
rect 31300 9522 31352 9528
rect 30564 9376 30616 9382
rect 30564 9318 30616 9324
rect 30748 9376 30800 9382
rect 30748 9318 30800 9324
rect 30576 8974 30604 9318
rect 30564 8968 30616 8974
rect 30102 8936 30158 8945
rect 30564 8910 30616 8916
rect 30102 8871 30104 8880
rect 30156 8871 30158 8880
rect 30104 8842 30156 8848
rect 29644 8492 29696 8498
rect 29644 8434 29696 8440
rect 30472 8492 30524 8498
rect 30472 8434 30524 8440
rect 29276 8356 29328 8362
rect 29276 8298 29328 8304
rect 29184 8288 29236 8294
rect 29184 8230 29236 8236
rect 28317 8188 28625 8197
rect 28317 8186 28323 8188
rect 28379 8186 28403 8188
rect 28459 8186 28483 8188
rect 28539 8186 28563 8188
rect 28619 8186 28625 8188
rect 28379 8134 28381 8186
rect 28561 8134 28563 8186
rect 28317 8132 28323 8134
rect 28379 8132 28403 8134
rect 28459 8132 28483 8134
rect 28539 8132 28563 8134
rect 28619 8132 28625 8134
rect 28317 8123 28625 8132
rect 27988 8084 28040 8090
rect 27988 8026 28040 8032
rect 27896 7948 27948 7954
rect 27896 7890 27948 7896
rect 28908 7948 28960 7954
rect 28908 7890 28960 7896
rect 27804 7812 27856 7818
rect 27804 7754 27856 7760
rect 28920 7478 28948 7890
rect 27896 7472 27948 7478
rect 27896 7414 27948 7420
rect 28908 7472 28960 7478
rect 28908 7414 28960 7420
rect 27160 7336 27212 7342
rect 27160 7278 27212 7284
rect 27068 6316 27120 6322
rect 27068 6258 27120 6264
rect 26240 5704 26292 5710
rect 26240 5646 26292 5652
rect 27172 5166 27200 7278
rect 27620 7200 27672 7206
rect 27620 7142 27672 7148
rect 27632 6866 27660 7142
rect 27620 6860 27672 6866
rect 27620 6802 27672 6808
rect 27252 6792 27304 6798
rect 27252 6734 27304 6740
rect 27264 6458 27292 6734
rect 27908 6662 27936 7414
rect 29196 7410 29224 8230
rect 29644 7880 29696 7886
rect 29644 7822 29696 7828
rect 29736 7880 29788 7886
rect 29736 7822 29788 7828
rect 29656 7410 29684 7822
rect 29184 7404 29236 7410
rect 29184 7346 29236 7352
rect 29644 7404 29696 7410
rect 29644 7346 29696 7352
rect 28724 7336 28776 7342
rect 28724 7278 28776 7284
rect 28317 7100 28625 7109
rect 28317 7098 28323 7100
rect 28379 7098 28403 7100
rect 28459 7098 28483 7100
rect 28539 7098 28563 7100
rect 28619 7098 28625 7100
rect 28379 7046 28381 7098
rect 28561 7046 28563 7098
rect 28317 7044 28323 7046
rect 28379 7044 28403 7046
rect 28459 7044 28483 7046
rect 28539 7044 28563 7046
rect 28619 7044 28625 7046
rect 28317 7035 28625 7044
rect 28736 6730 28764 7278
rect 28724 6724 28776 6730
rect 28724 6666 28776 6672
rect 27896 6656 27948 6662
rect 27896 6598 27948 6604
rect 27252 6452 27304 6458
rect 27252 6394 27304 6400
rect 27620 6316 27672 6322
rect 27620 6258 27672 6264
rect 27526 6216 27582 6225
rect 27526 6151 27582 6160
rect 27540 5817 27568 6151
rect 27632 5914 27660 6258
rect 28317 6012 28625 6021
rect 28317 6010 28323 6012
rect 28379 6010 28403 6012
rect 28459 6010 28483 6012
rect 28539 6010 28563 6012
rect 28619 6010 28625 6012
rect 28379 5958 28381 6010
rect 28561 5958 28563 6010
rect 28317 5956 28323 5958
rect 28379 5956 28403 5958
rect 28459 5956 28483 5958
rect 28539 5956 28563 5958
rect 28619 5956 28625 5958
rect 28317 5947 28625 5956
rect 27620 5908 27672 5914
rect 27620 5850 27672 5856
rect 27526 5808 27582 5817
rect 27526 5743 27582 5752
rect 27344 5228 27396 5234
rect 27344 5170 27396 5176
rect 27160 5160 27212 5166
rect 27160 5102 27212 5108
rect 27356 4826 27384 5170
rect 27344 4820 27396 4826
rect 27344 4762 27396 4768
rect 26884 4548 26936 4554
rect 26884 4490 26936 4496
rect 26056 4140 26108 4146
rect 26056 4082 26108 4088
rect 25964 4072 26016 4078
rect 25964 4014 26016 4020
rect 24952 3936 25004 3942
rect 24952 3878 25004 3884
rect 24964 3534 24992 3878
rect 26068 3738 26096 4082
rect 26896 3738 26924 4490
rect 26976 3936 27028 3942
rect 26976 3878 27028 3884
rect 26056 3732 26108 3738
rect 26056 3674 26108 3680
rect 26884 3732 26936 3738
rect 26884 3674 26936 3680
rect 26988 3534 27016 3878
rect 24032 3528 24084 3534
rect 24032 3470 24084 3476
rect 24952 3528 25004 3534
rect 24952 3470 25004 3476
rect 26976 3528 27028 3534
rect 26976 3470 27028 3476
rect 23296 3460 23348 3466
rect 23296 3402 23348 3408
rect 22843 3292 23151 3301
rect 22843 3290 22849 3292
rect 22905 3290 22929 3292
rect 22985 3290 23009 3292
rect 23065 3290 23089 3292
rect 23145 3290 23151 3292
rect 22905 3238 22907 3290
rect 23087 3238 23089 3290
rect 22843 3236 22849 3238
rect 22905 3236 22929 3238
rect 22985 3236 23009 3238
rect 23065 3236 23089 3238
rect 23145 3236 23151 3238
rect 22843 3227 23151 3236
rect 22652 3052 22704 3058
rect 22652 2994 22704 3000
rect 22560 2984 22612 2990
rect 22560 2926 22612 2932
rect 18880 2848 18932 2854
rect 18880 2790 18932 2796
rect 18892 2582 18920 2790
rect 18880 2576 18932 2582
rect 18880 2518 18932 2524
rect 18144 2508 18196 2514
rect 18144 2450 18196 2456
rect 16856 2440 16908 2446
rect 16856 2382 16908 2388
rect 17408 2440 17460 2446
rect 17408 2382 17460 2388
rect 19340 2440 19392 2446
rect 19340 2382 19392 2388
rect 20720 2440 20772 2446
rect 20720 2382 20772 2388
rect 17420 800 17448 2382
rect 19352 800 19380 2382
rect 20732 898 20760 2382
rect 20640 870 20760 898
rect 20640 800 20668 870
rect 22572 800 22600 2926
rect 27540 2650 27568 5743
rect 28736 5370 28764 6666
rect 29196 6254 29224 7346
rect 29748 6798 29776 7822
rect 29736 6792 29788 6798
rect 29736 6734 29788 6740
rect 29276 6316 29328 6322
rect 29276 6258 29328 6264
rect 29184 6248 29236 6254
rect 29184 6190 29236 6196
rect 29000 6112 29052 6118
rect 29000 6054 29052 6060
rect 29092 6112 29144 6118
rect 29092 6054 29144 6060
rect 28724 5364 28776 5370
rect 28724 5306 28776 5312
rect 29012 5302 29040 6054
rect 29000 5296 29052 5302
rect 29000 5238 29052 5244
rect 29104 5166 29132 6054
rect 29196 5574 29224 6190
rect 29288 5914 29316 6258
rect 29276 5908 29328 5914
rect 29276 5850 29328 5856
rect 29748 5846 29776 6734
rect 30380 6656 30432 6662
rect 30380 6598 30432 6604
rect 30012 6248 30064 6254
rect 30012 6190 30064 6196
rect 29828 6112 29880 6118
rect 29828 6054 29880 6060
rect 29920 6112 29972 6118
rect 29920 6054 29972 6060
rect 29736 5840 29788 5846
rect 29736 5782 29788 5788
rect 29840 5710 29868 6054
rect 29932 5778 29960 6054
rect 29920 5772 29972 5778
rect 29920 5714 29972 5720
rect 29828 5704 29880 5710
rect 29828 5646 29880 5652
rect 29184 5568 29236 5574
rect 29184 5510 29236 5516
rect 29840 5166 29868 5646
rect 29092 5160 29144 5166
rect 29092 5102 29144 5108
rect 29828 5160 29880 5166
rect 29828 5102 29880 5108
rect 29368 5024 29420 5030
rect 29368 4966 29420 4972
rect 28317 4924 28625 4933
rect 28317 4922 28323 4924
rect 28379 4922 28403 4924
rect 28459 4922 28483 4924
rect 28539 4922 28563 4924
rect 28619 4922 28625 4924
rect 28379 4870 28381 4922
rect 28561 4870 28563 4922
rect 28317 4868 28323 4870
rect 28379 4868 28403 4870
rect 28459 4868 28483 4870
rect 28539 4868 28563 4870
rect 28619 4868 28625 4870
rect 28317 4859 28625 4868
rect 29380 4690 29408 4966
rect 30024 4758 30052 6190
rect 30392 5710 30420 6598
rect 30484 5710 30512 8434
rect 30564 7812 30616 7818
rect 30564 7754 30616 7760
rect 30576 6458 30604 7754
rect 30656 7472 30708 7478
rect 30656 7414 30708 7420
rect 30668 7206 30696 7414
rect 30656 7200 30708 7206
rect 30656 7142 30708 7148
rect 30668 6458 30696 7142
rect 30564 6452 30616 6458
rect 30564 6394 30616 6400
rect 30656 6452 30708 6458
rect 30656 6394 30708 6400
rect 30760 6322 30788 9318
rect 31128 7546 31156 9522
rect 31208 8832 31260 8838
rect 31208 8774 31260 8780
rect 31116 7540 31168 7546
rect 31116 7482 31168 7488
rect 31024 6724 31076 6730
rect 31024 6666 31076 6672
rect 31036 6458 31064 6666
rect 31024 6452 31076 6458
rect 31024 6394 31076 6400
rect 30748 6316 30800 6322
rect 30748 6258 30800 6264
rect 30656 5772 30708 5778
rect 30656 5714 30708 5720
rect 30380 5704 30432 5710
rect 30380 5646 30432 5652
rect 30472 5704 30524 5710
rect 30472 5646 30524 5652
rect 30012 4752 30064 4758
rect 30012 4694 30064 4700
rect 29368 4684 29420 4690
rect 29368 4626 29420 4632
rect 29000 4616 29052 4622
rect 29000 4558 29052 4564
rect 29012 4146 29040 4558
rect 29380 4146 29408 4626
rect 29736 4480 29788 4486
rect 29736 4422 29788 4428
rect 29748 4214 29776 4422
rect 29736 4208 29788 4214
rect 29736 4150 29788 4156
rect 29000 4140 29052 4146
rect 29000 4082 29052 4088
rect 29368 4140 29420 4146
rect 29368 4082 29420 4088
rect 28317 3836 28625 3845
rect 28317 3834 28323 3836
rect 28379 3834 28403 3836
rect 28459 3834 28483 3836
rect 28539 3834 28563 3836
rect 28619 3834 28625 3836
rect 28379 3782 28381 3834
rect 28561 3782 28563 3834
rect 28317 3780 28323 3782
rect 28379 3780 28403 3782
rect 28459 3780 28483 3782
rect 28539 3780 28563 3782
rect 28619 3780 28625 3782
rect 28317 3771 28625 3780
rect 30024 3602 30052 4694
rect 30564 4616 30616 4622
rect 30564 4558 30616 4564
rect 30380 4480 30432 4486
rect 30380 4422 30432 4428
rect 30392 4078 30420 4422
rect 30380 4072 30432 4078
rect 30380 4014 30432 4020
rect 30576 3670 30604 4558
rect 30564 3664 30616 3670
rect 30564 3606 30616 3612
rect 30012 3596 30064 3602
rect 30012 3538 30064 3544
rect 28317 2748 28625 2757
rect 28317 2746 28323 2748
rect 28379 2746 28403 2748
rect 28459 2746 28483 2748
rect 28539 2746 28563 2748
rect 28619 2746 28625 2748
rect 28379 2694 28381 2746
rect 28561 2694 28563 2746
rect 28317 2692 28323 2694
rect 28379 2692 28403 2694
rect 28459 2692 28483 2694
rect 28539 2692 28563 2694
rect 28619 2692 28625 2694
rect 28317 2683 28625 2692
rect 27528 2644 27580 2650
rect 27528 2586 27580 2592
rect 23848 2440 23900 2446
rect 23848 2382 23900 2388
rect 25780 2440 25832 2446
rect 25780 2382 25832 2388
rect 29000 2440 29052 2446
rect 29000 2382 29052 2388
rect 30380 2440 30432 2446
rect 30380 2382 30432 2388
rect 22843 2204 23151 2213
rect 22843 2202 22849 2204
rect 22905 2202 22929 2204
rect 22985 2202 23009 2204
rect 23065 2202 23089 2204
rect 23145 2202 23151 2204
rect 22905 2150 22907 2202
rect 23087 2150 23089 2202
rect 22843 2148 22849 2150
rect 22905 2148 22929 2150
rect 22985 2148 23009 2150
rect 23065 2148 23089 2150
rect 23145 2148 23151 2150
rect 22843 2139 23151 2148
rect 23860 800 23888 2382
rect 25792 800 25820 2382
rect 27068 2372 27120 2378
rect 27068 2314 27120 2320
rect 27080 800 27108 2314
rect 29012 800 29040 2382
rect 30392 898 30420 2382
rect 30668 2310 30696 5714
rect 30748 5568 30800 5574
rect 30748 5510 30800 5516
rect 30760 5030 30788 5510
rect 30748 5024 30800 5030
rect 30748 4966 30800 4972
rect 31220 4146 31248 8774
rect 31312 8634 31340 9522
rect 31404 9110 31432 10662
rect 31588 9994 31616 11290
rect 31864 10130 31892 12242
rect 32324 11762 32352 12718
rect 32496 12096 32548 12102
rect 32496 12038 32548 12044
rect 32508 11762 32536 12038
rect 32784 11898 32812 13262
rect 33790 13084 34098 13093
rect 33790 13082 33796 13084
rect 33852 13082 33876 13084
rect 33932 13082 33956 13084
rect 34012 13082 34036 13084
rect 34092 13082 34098 13084
rect 33852 13030 33854 13082
rect 34034 13030 34036 13082
rect 33790 13028 33796 13030
rect 33852 13028 33876 13030
rect 33932 13028 33956 13030
rect 34012 13028 34036 13030
rect 34092 13028 34098 13030
rect 33790 13019 34098 13028
rect 33324 12844 33376 12850
rect 33324 12786 33376 12792
rect 33140 12640 33192 12646
rect 33140 12582 33192 12588
rect 33152 12170 33180 12582
rect 33336 12442 33364 12786
rect 34336 12708 34388 12714
rect 34336 12650 34388 12656
rect 33324 12436 33376 12442
rect 33324 12378 33376 12384
rect 34348 12238 34376 12650
rect 35912 12434 35940 14418
rect 36096 14278 36124 16000
rect 36176 15982 36228 15988
rect 36636 15904 36688 15910
rect 36636 15846 36688 15852
rect 36268 15428 36320 15434
rect 36268 15370 36320 15376
rect 36176 15360 36228 15366
rect 36176 15302 36228 15308
rect 36188 14890 36216 15302
rect 36176 14884 36228 14890
rect 36176 14826 36228 14832
rect 36280 14822 36308 15370
rect 36648 15026 36676 15846
rect 36636 15020 36688 15026
rect 36636 14962 36688 14968
rect 37096 14884 37148 14890
rect 37096 14826 37148 14832
rect 36268 14816 36320 14822
rect 36268 14758 36320 14764
rect 36452 14816 36504 14822
rect 36452 14758 36504 14764
rect 36280 14550 36308 14758
rect 36268 14544 36320 14550
rect 36268 14486 36320 14492
rect 36360 14408 36412 14414
rect 36360 14350 36412 14356
rect 36084 14272 36136 14278
rect 36084 14214 36136 14220
rect 36268 14272 36320 14278
rect 36268 14214 36320 14220
rect 36280 13870 36308 14214
rect 36268 13864 36320 13870
rect 36268 13806 36320 13812
rect 36372 13530 36400 14350
rect 36464 14346 36492 14758
rect 37108 14414 37136 14826
rect 38200 14476 38252 14482
rect 38200 14418 38252 14424
rect 37096 14408 37148 14414
rect 37096 14350 37148 14356
rect 36452 14340 36504 14346
rect 36452 14282 36504 14288
rect 37832 14272 37884 14278
rect 37832 14214 37884 14220
rect 37844 14074 37872 14214
rect 37832 14068 37884 14074
rect 37832 14010 37884 14016
rect 36452 13864 36504 13870
rect 36452 13806 36504 13812
rect 36360 13524 36412 13530
rect 36360 13466 36412 13472
rect 36084 12844 36136 12850
rect 36084 12786 36136 12792
rect 35820 12406 35940 12434
rect 33600 12232 33652 12238
rect 33600 12174 33652 12180
rect 34336 12232 34388 12238
rect 34336 12174 34388 12180
rect 34888 12232 34940 12238
rect 34888 12174 34940 12180
rect 33140 12164 33192 12170
rect 33140 12106 33192 12112
rect 32772 11892 32824 11898
rect 32772 11834 32824 11840
rect 33612 11762 33640 12174
rect 33790 11996 34098 12005
rect 33790 11994 33796 11996
rect 33852 11994 33876 11996
rect 33932 11994 33956 11996
rect 34012 11994 34036 11996
rect 34092 11994 34098 11996
rect 33852 11942 33854 11994
rect 34034 11942 34036 11994
rect 33790 11940 33796 11942
rect 33852 11940 33876 11942
rect 33932 11940 33956 11942
rect 34012 11940 34036 11942
rect 34092 11940 34098 11942
rect 33790 11931 34098 11940
rect 32312 11756 32364 11762
rect 32312 11698 32364 11704
rect 32496 11756 32548 11762
rect 32496 11698 32548 11704
rect 33600 11756 33652 11762
rect 33652 11716 33732 11744
rect 33600 11698 33652 11704
rect 32220 11552 32272 11558
rect 32220 11494 32272 11500
rect 32232 11218 32260 11494
rect 32220 11212 32272 11218
rect 32220 11154 32272 11160
rect 32312 11144 32364 11150
rect 32312 11086 32364 11092
rect 33600 11144 33652 11150
rect 33600 11086 33652 11092
rect 31852 10124 31904 10130
rect 31852 10066 31904 10072
rect 32220 10124 32272 10130
rect 32220 10066 32272 10072
rect 31576 9988 31628 9994
rect 31576 9930 31628 9936
rect 31668 9716 31720 9722
rect 31668 9658 31720 9664
rect 31392 9104 31444 9110
rect 31392 9046 31444 9052
rect 31484 8968 31536 8974
rect 31536 8928 31616 8956
rect 31484 8910 31536 8916
rect 31300 8628 31352 8634
rect 31300 8570 31352 8576
rect 31588 8498 31616 8928
rect 31576 8492 31628 8498
rect 31576 8434 31628 8440
rect 31484 8424 31536 8430
rect 31484 8366 31536 8372
rect 31392 7540 31444 7546
rect 31496 7528 31524 8366
rect 31588 8022 31616 8434
rect 31680 8430 31708 9658
rect 32232 9586 32260 10066
rect 32220 9580 32272 9586
rect 32220 9522 32272 9528
rect 32324 9450 32352 11086
rect 33140 11008 33192 11014
rect 33140 10950 33192 10956
rect 33508 11008 33560 11014
rect 33508 10950 33560 10956
rect 33152 10606 33180 10950
rect 33520 10742 33548 10950
rect 33508 10736 33560 10742
rect 33508 10678 33560 10684
rect 33140 10600 33192 10606
rect 33140 10542 33192 10548
rect 32404 10464 32456 10470
rect 32404 10406 32456 10412
rect 32416 10062 32444 10406
rect 33612 10266 33640 11086
rect 33600 10260 33652 10266
rect 33600 10202 33652 10208
rect 33704 10062 33732 11716
rect 34796 11076 34848 11082
rect 34796 11018 34848 11024
rect 34520 11008 34572 11014
rect 34520 10950 34572 10956
rect 33790 10908 34098 10917
rect 33790 10906 33796 10908
rect 33852 10906 33876 10908
rect 33932 10906 33956 10908
rect 34012 10906 34036 10908
rect 34092 10906 34098 10908
rect 33852 10854 33854 10906
rect 34034 10854 34036 10906
rect 33790 10852 33796 10854
rect 33852 10852 33876 10854
rect 33932 10852 33956 10854
rect 34012 10852 34036 10854
rect 34092 10852 34098 10854
rect 33790 10843 34098 10852
rect 34532 10062 34560 10950
rect 32404 10056 32456 10062
rect 32404 9998 32456 10004
rect 33692 10056 33744 10062
rect 33692 9998 33744 10004
rect 34520 10056 34572 10062
rect 34520 9998 34572 10004
rect 34808 9994 34836 11018
rect 34900 10538 34928 12174
rect 35820 11286 35848 12406
rect 35900 11756 35952 11762
rect 35900 11698 35952 11704
rect 35808 11280 35860 11286
rect 35808 11222 35860 11228
rect 35072 11144 35124 11150
rect 35070 11112 35072 11121
rect 35124 11112 35126 11121
rect 35820 11082 35848 11222
rect 35070 11047 35126 11056
rect 35808 11076 35860 11082
rect 35808 11018 35860 11024
rect 34888 10532 34940 10538
rect 34888 10474 34940 10480
rect 34900 10130 34928 10474
rect 35164 10464 35216 10470
rect 35164 10406 35216 10412
rect 35176 10130 35204 10406
rect 35912 10130 35940 11698
rect 35992 11688 36044 11694
rect 35992 11630 36044 11636
rect 36004 11150 36032 11630
rect 36096 11218 36124 12786
rect 36360 11756 36412 11762
rect 36360 11698 36412 11704
rect 36084 11212 36136 11218
rect 36084 11154 36136 11160
rect 35992 11144 36044 11150
rect 35992 11086 36044 11092
rect 36176 11144 36228 11150
rect 36176 11086 36228 11092
rect 34888 10124 34940 10130
rect 34888 10066 34940 10072
rect 35164 10124 35216 10130
rect 35164 10066 35216 10072
rect 35900 10124 35952 10130
rect 35900 10066 35952 10072
rect 34796 9988 34848 9994
rect 34796 9930 34848 9936
rect 32956 9920 33008 9926
rect 32956 9862 33008 9868
rect 32864 9648 32916 9654
rect 32864 9590 32916 9596
rect 32876 9489 32904 9590
rect 32968 9586 32996 9862
rect 33790 9820 34098 9829
rect 33790 9818 33796 9820
rect 33852 9818 33876 9820
rect 33932 9818 33956 9820
rect 34012 9818 34036 9820
rect 34092 9818 34098 9820
rect 33852 9766 33854 9818
rect 34034 9766 34036 9818
rect 33790 9764 33796 9766
rect 33852 9764 33876 9766
rect 33932 9764 33956 9766
rect 34012 9764 34036 9766
rect 34092 9764 34098 9766
rect 33790 9755 34098 9764
rect 35912 9722 35940 10066
rect 36004 9926 36032 11086
rect 35992 9920 36044 9926
rect 35992 9862 36044 9868
rect 35900 9716 35952 9722
rect 35900 9658 35952 9664
rect 35164 9648 35216 9654
rect 35164 9590 35216 9596
rect 32956 9580 33008 9586
rect 32956 9522 33008 9528
rect 33416 9580 33468 9586
rect 33416 9522 33468 9528
rect 32862 9480 32918 9489
rect 32220 9444 32272 9450
rect 32220 9386 32272 9392
rect 32312 9444 32364 9450
rect 32862 9415 32918 9424
rect 32312 9386 32364 9392
rect 32232 9042 32260 9386
rect 32220 9036 32272 9042
rect 32220 8978 32272 8984
rect 32494 8936 32550 8945
rect 32494 8871 32550 8880
rect 31852 8560 31904 8566
rect 31852 8502 31904 8508
rect 31668 8424 31720 8430
rect 31668 8366 31720 8372
rect 31760 8356 31812 8362
rect 31760 8298 31812 8304
rect 31576 8016 31628 8022
rect 31576 7958 31628 7964
rect 31444 7500 31524 7528
rect 31392 7482 31444 7488
rect 31392 7404 31444 7410
rect 31392 7346 31444 7352
rect 31404 6458 31432 7346
rect 31496 7206 31524 7500
rect 31588 7342 31616 7958
rect 31772 7410 31800 8298
rect 31864 7478 31892 8502
rect 31944 7812 31996 7818
rect 31944 7754 31996 7760
rect 31956 7478 31984 7754
rect 31852 7472 31904 7478
rect 31852 7414 31904 7420
rect 31944 7472 31996 7478
rect 31944 7414 31996 7420
rect 31760 7404 31812 7410
rect 31760 7346 31812 7352
rect 31576 7336 31628 7342
rect 31576 7278 31628 7284
rect 31864 7274 31892 7414
rect 31852 7268 31904 7274
rect 31852 7210 31904 7216
rect 31484 7200 31536 7206
rect 31484 7142 31536 7148
rect 31956 6730 31984 7414
rect 32220 7404 32272 7410
rect 32220 7346 32272 7352
rect 32036 7200 32088 7206
rect 32036 7142 32088 7148
rect 31944 6724 31996 6730
rect 31944 6666 31996 6672
rect 32048 6662 32076 7142
rect 32232 6866 32260 7346
rect 32404 7336 32456 7342
rect 32404 7278 32456 7284
rect 32416 7206 32444 7278
rect 32312 7200 32364 7206
rect 32312 7142 32364 7148
rect 32404 7200 32456 7206
rect 32404 7142 32456 7148
rect 32220 6860 32272 6866
rect 32220 6802 32272 6808
rect 32036 6656 32088 6662
rect 32036 6598 32088 6604
rect 31392 6452 31444 6458
rect 31392 6394 31444 6400
rect 32324 6322 32352 7142
rect 32416 6934 32444 7142
rect 32404 6928 32456 6934
rect 32404 6870 32456 6876
rect 32312 6316 32364 6322
rect 32312 6258 32364 6264
rect 31208 4140 31260 4146
rect 31208 4082 31260 4088
rect 31220 3534 31248 4082
rect 31208 3528 31260 3534
rect 31208 3470 31260 3476
rect 32508 2650 32536 8871
rect 32968 8090 32996 9522
rect 33428 8401 33456 9522
rect 35176 9178 35204 9590
rect 35164 9172 35216 9178
rect 35164 9114 35216 9120
rect 35808 9104 35860 9110
rect 35808 9046 35860 9052
rect 35256 9036 35308 9042
rect 35256 8978 35308 8984
rect 34152 8968 34204 8974
rect 34152 8910 34204 8916
rect 33790 8732 34098 8741
rect 33790 8730 33796 8732
rect 33852 8730 33876 8732
rect 33932 8730 33956 8732
rect 34012 8730 34036 8732
rect 34092 8730 34098 8732
rect 33852 8678 33854 8730
rect 34034 8678 34036 8730
rect 33790 8676 33796 8678
rect 33852 8676 33876 8678
rect 33932 8676 33956 8678
rect 34012 8676 34036 8678
rect 34092 8676 34098 8678
rect 33790 8667 34098 8676
rect 33414 8392 33470 8401
rect 34164 8362 34192 8910
rect 35072 8900 35124 8906
rect 35072 8842 35124 8848
rect 34518 8528 34574 8537
rect 34518 8463 34574 8472
rect 34532 8430 34560 8463
rect 34520 8424 34572 8430
rect 34520 8366 34572 8372
rect 33414 8327 33470 8336
rect 34152 8356 34204 8362
rect 34152 8298 34204 8304
rect 32956 8084 33008 8090
rect 32956 8026 33008 8032
rect 32954 7984 33010 7993
rect 32954 7919 33010 7928
rect 34336 7948 34388 7954
rect 32588 7880 32640 7886
rect 32588 7822 32640 7828
rect 32600 7410 32628 7822
rect 32968 7546 32996 7919
rect 34336 7890 34388 7896
rect 33790 7644 34098 7653
rect 33790 7642 33796 7644
rect 33852 7642 33876 7644
rect 33932 7642 33956 7644
rect 34012 7642 34036 7644
rect 34092 7642 34098 7644
rect 33852 7590 33854 7642
rect 34034 7590 34036 7642
rect 33790 7588 33796 7590
rect 33852 7588 33876 7590
rect 33932 7588 33956 7590
rect 34012 7588 34036 7590
rect 34092 7588 34098 7590
rect 33790 7579 34098 7588
rect 34348 7546 34376 7890
rect 35084 7886 35112 8842
rect 35072 7880 35124 7886
rect 35072 7822 35124 7828
rect 35164 7880 35216 7886
rect 35164 7822 35216 7828
rect 34428 7744 34480 7750
rect 34428 7686 34480 7692
rect 32956 7540 33008 7546
rect 32956 7482 33008 7488
rect 34336 7540 34388 7546
rect 34336 7482 34388 7488
rect 32968 7410 32996 7482
rect 33784 7472 33836 7478
rect 33784 7414 33836 7420
rect 32588 7404 32640 7410
rect 32588 7346 32640 7352
rect 32680 7404 32732 7410
rect 32680 7346 32732 7352
rect 32772 7404 32824 7410
rect 32772 7346 32824 7352
rect 32956 7404 33008 7410
rect 32956 7346 33008 7352
rect 33048 7404 33100 7410
rect 33048 7346 33100 7352
rect 33692 7404 33744 7410
rect 33692 7346 33744 7352
rect 32588 7268 32640 7274
rect 32588 7210 32640 7216
rect 32600 6934 32628 7210
rect 32588 6928 32640 6934
rect 32588 6870 32640 6876
rect 32600 6798 32628 6870
rect 32588 6792 32640 6798
rect 32588 6734 32640 6740
rect 32692 6662 32720 7346
rect 32784 7002 32812 7346
rect 32772 6996 32824 7002
rect 32772 6938 32824 6944
rect 33060 6866 33088 7346
rect 33048 6860 33100 6866
rect 33048 6802 33100 6808
rect 32680 6656 32732 6662
rect 32680 6598 32732 6604
rect 33704 6254 33732 7346
rect 33796 7206 33824 7414
rect 34336 7404 34388 7410
rect 34336 7346 34388 7352
rect 34244 7268 34296 7274
rect 34244 7210 34296 7216
rect 33784 7200 33836 7206
rect 33784 7142 33836 7148
rect 33796 6798 33824 7142
rect 33784 6792 33836 6798
rect 33784 6734 33836 6740
rect 34152 6656 34204 6662
rect 34152 6598 34204 6604
rect 33790 6556 34098 6565
rect 33790 6554 33796 6556
rect 33852 6554 33876 6556
rect 33932 6554 33956 6556
rect 34012 6554 34036 6556
rect 34092 6554 34098 6556
rect 33852 6502 33854 6554
rect 34034 6502 34036 6554
rect 33790 6500 33796 6502
rect 33852 6500 33876 6502
rect 33932 6500 33956 6502
rect 34012 6500 34036 6502
rect 34092 6500 34098 6502
rect 33790 6491 34098 6500
rect 33876 6452 33928 6458
rect 33876 6394 33928 6400
rect 33888 6322 33916 6394
rect 33876 6316 33928 6322
rect 33876 6258 33928 6264
rect 34060 6316 34112 6322
rect 34164 6304 34192 6598
rect 34112 6276 34192 6304
rect 34060 6258 34112 6264
rect 33692 6248 33744 6254
rect 33692 6190 33744 6196
rect 33416 6112 33468 6118
rect 33416 6054 33468 6060
rect 33428 5234 33456 6054
rect 34072 5710 34100 6258
rect 34256 5914 34284 7210
rect 34348 5914 34376 7346
rect 34440 6905 34468 7686
rect 35084 7274 35112 7822
rect 35072 7268 35124 7274
rect 35072 7210 35124 7216
rect 34796 7200 34848 7206
rect 34796 7142 34848 7148
rect 34426 6896 34482 6905
rect 34426 6831 34482 6840
rect 34428 6452 34480 6458
rect 34428 6394 34480 6400
rect 34244 5908 34296 5914
rect 34244 5850 34296 5856
rect 34336 5908 34388 5914
rect 34336 5850 34388 5856
rect 34440 5710 34468 6394
rect 34520 6248 34572 6254
rect 34520 6190 34572 6196
rect 34532 6089 34560 6190
rect 34518 6080 34574 6089
rect 34518 6015 34574 6024
rect 34808 5710 34836 7142
rect 34888 6792 34940 6798
rect 34888 6734 34940 6740
rect 34060 5704 34112 5710
rect 34060 5646 34112 5652
rect 34428 5704 34480 5710
rect 34428 5646 34480 5652
rect 34796 5704 34848 5710
rect 34900 5681 34928 6734
rect 35084 6390 35112 7210
rect 35176 6866 35204 7822
rect 35268 7342 35296 8978
rect 35624 8968 35676 8974
rect 35452 8928 35624 8956
rect 35452 8498 35480 8928
rect 35624 8910 35676 8916
rect 35624 8832 35676 8838
rect 35624 8774 35676 8780
rect 35716 8832 35768 8838
rect 35716 8774 35768 8780
rect 35636 8634 35664 8774
rect 35624 8628 35676 8634
rect 35624 8570 35676 8576
rect 35728 8566 35756 8774
rect 35716 8560 35768 8566
rect 35716 8502 35768 8508
rect 35820 8498 35848 9046
rect 36084 8560 36136 8566
rect 36084 8502 36136 8508
rect 35440 8492 35492 8498
rect 35440 8434 35492 8440
rect 35808 8492 35860 8498
rect 35808 8434 35860 8440
rect 35992 8424 36044 8430
rect 35992 8366 36044 8372
rect 36004 7410 36032 8366
rect 36096 7993 36124 8502
rect 36188 8294 36216 11086
rect 36372 10266 36400 11698
rect 36464 11694 36492 13806
rect 36636 13728 36688 13734
rect 36636 13670 36688 13676
rect 36648 13326 36676 13670
rect 37844 13530 37872 14010
rect 38212 13870 38240 14418
rect 38856 14385 38884 16934
rect 39264 16892 39572 16901
rect 39264 16890 39270 16892
rect 39326 16890 39350 16892
rect 39406 16890 39430 16892
rect 39486 16890 39510 16892
rect 39566 16890 39572 16892
rect 39326 16838 39328 16890
rect 39508 16838 39510 16890
rect 39264 16836 39270 16838
rect 39326 16836 39350 16838
rect 39406 16836 39430 16838
rect 39486 16836 39510 16838
rect 39566 16836 39572 16838
rect 39264 16827 39572 16836
rect 40604 16046 40632 19200
rect 41892 19106 41920 19200
rect 41880 19100 41932 19106
rect 41880 19042 41932 19048
rect 42800 19100 42852 19106
rect 42800 19042 42852 19048
rect 42812 17202 42840 19042
rect 43444 18080 43496 18086
rect 43444 18022 43496 18028
rect 43456 17202 43484 18022
rect 43824 17202 43852 19200
rect 45006 19136 45062 19145
rect 45006 19071 45062 19080
rect 45020 18086 45048 19071
rect 45008 18080 45060 18086
rect 45008 18022 45060 18028
rect 45006 17776 45062 17785
rect 45006 17711 45062 17720
rect 45020 17542 45048 17711
rect 43996 17536 44048 17542
rect 43996 17478 44048 17484
rect 45008 17536 45060 17542
rect 45008 17478 45060 17484
rect 42800 17196 42852 17202
rect 42800 17138 42852 17144
rect 43444 17196 43496 17202
rect 43444 17138 43496 17144
rect 43812 17196 43864 17202
rect 43812 17138 43864 17144
rect 41604 16108 41656 16114
rect 41604 16050 41656 16056
rect 40592 16040 40644 16046
rect 40592 15982 40644 15988
rect 41512 16040 41564 16046
rect 41512 15982 41564 15988
rect 39264 15804 39572 15813
rect 39264 15802 39270 15804
rect 39326 15802 39350 15804
rect 39406 15802 39430 15804
rect 39486 15802 39510 15804
rect 39566 15802 39572 15804
rect 39326 15750 39328 15802
rect 39508 15750 39510 15802
rect 39264 15748 39270 15750
rect 39326 15748 39350 15750
rect 39406 15748 39430 15750
rect 39486 15748 39510 15750
rect 39566 15748 39572 15750
rect 39264 15739 39572 15748
rect 41420 15496 41472 15502
rect 41420 15438 41472 15444
rect 40132 15020 40184 15026
rect 40132 14962 40184 14968
rect 38936 14952 38988 14958
rect 38936 14894 38988 14900
rect 38842 14376 38898 14385
rect 38842 14311 38898 14320
rect 38856 13938 38884 14311
rect 38384 13932 38436 13938
rect 38384 13874 38436 13880
rect 38844 13932 38896 13938
rect 38844 13874 38896 13880
rect 37924 13864 37976 13870
rect 37924 13806 37976 13812
rect 38200 13864 38252 13870
rect 38200 13806 38252 13812
rect 37832 13524 37884 13530
rect 37832 13466 37884 13472
rect 36636 13320 36688 13326
rect 36636 13262 36688 13268
rect 37096 13252 37148 13258
rect 37096 13194 37148 13200
rect 36544 12640 36596 12646
rect 36544 12582 36596 12588
rect 36556 12170 36584 12582
rect 36544 12164 36596 12170
rect 36544 12106 36596 12112
rect 36636 12096 36688 12102
rect 36636 12038 36688 12044
rect 36452 11688 36504 11694
rect 36452 11630 36504 11636
rect 36648 11558 36676 12038
rect 37108 11830 37136 13194
rect 37648 12844 37700 12850
rect 37648 12786 37700 12792
rect 37464 12640 37516 12646
rect 37464 12582 37516 12588
rect 37476 12170 37504 12582
rect 37464 12164 37516 12170
rect 37464 12106 37516 12112
rect 37660 11898 37688 12786
rect 37648 11892 37700 11898
rect 37648 11834 37700 11840
rect 37096 11824 37148 11830
rect 37096 11766 37148 11772
rect 37188 11824 37240 11830
rect 37188 11766 37240 11772
rect 36636 11552 36688 11558
rect 36636 11494 36688 11500
rect 37200 11150 37228 11766
rect 37280 11756 37332 11762
rect 37280 11698 37332 11704
rect 37292 11150 37320 11698
rect 37936 11558 37964 13806
rect 38108 13184 38160 13190
rect 38108 13126 38160 13132
rect 38120 12170 38148 13126
rect 38212 12986 38240 13806
rect 38396 13462 38424 13874
rect 38948 13734 38976 14894
rect 39672 14816 39724 14822
rect 39672 14758 39724 14764
rect 39264 14716 39572 14725
rect 39264 14714 39270 14716
rect 39326 14714 39350 14716
rect 39406 14714 39430 14716
rect 39486 14714 39510 14716
rect 39566 14714 39572 14716
rect 39326 14662 39328 14714
rect 39508 14662 39510 14714
rect 39264 14660 39270 14662
rect 39326 14660 39350 14662
rect 39406 14660 39430 14662
rect 39486 14660 39510 14662
rect 39566 14660 39572 14662
rect 39264 14651 39572 14660
rect 39684 14414 39712 14758
rect 39672 14408 39724 14414
rect 39672 14350 39724 14356
rect 40040 14408 40092 14414
rect 40040 14350 40092 14356
rect 40052 14006 40080 14350
rect 40144 14074 40172 14962
rect 41432 14074 41460 15438
rect 40132 14068 40184 14074
rect 40132 14010 40184 14016
rect 41420 14068 41472 14074
rect 41420 14010 41472 14016
rect 40040 14000 40092 14006
rect 40040 13942 40092 13948
rect 38936 13728 38988 13734
rect 38936 13670 38988 13676
rect 38384 13456 38436 13462
rect 38384 13398 38436 13404
rect 38200 12980 38252 12986
rect 38200 12922 38252 12928
rect 38396 12850 38424 13398
rect 38948 12918 38976 13670
rect 39264 13628 39572 13637
rect 39264 13626 39270 13628
rect 39326 13626 39350 13628
rect 39406 13626 39430 13628
rect 39486 13626 39510 13628
rect 39566 13626 39572 13628
rect 39326 13574 39328 13626
rect 39508 13574 39510 13626
rect 39264 13572 39270 13574
rect 39326 13572 39350 13574
rect 39406 13572 39430 13574
rect 39486 13572 39510 13574
rect 39566 13572 39572 13574
rect 39264 13563 39572 13572
rect 38936 12912 38988 12918
rect 38936 12854 38988 12860
rect 40040 12912 40092 12918
rect 40040 12854 40092 12860
rect 38384 12844 38436 12850
rect 38384 12786 38436 12792
rect 38396 12434 38424 12786
rect 38660 12776 38712 12782
rect 38660 12718 38712 12724
rect 38672 12442 38700 12718
rect 39264 12540 39572 12549
rect 39264 12538 39270 12540
rect 39326 12538 39350 12540
rect 39406 12538 39430 12540
rect 39486 12538 39510 12540
rect 39566 12538 39572 12540
rect 39326 12486 39328 12538
rect 39508 12486 39510 12538
rect 39264 12484 39270 12486
rect 39326 12484 39350 12486
rect 39406 12484 39430 12486
rect 39486 12484 39510 12486
rect 39566 12484 39572 12486
rect 39264 12475 39572 12484
rect 40052 12442 40080 12854
rect 41052 12844 41104 12850
rect 41052 12786 41104 12792
rect 40960 12640 41012 12646
rect 40960 12582 41012 12588
rect 38212 12406 38424 12434
rect 38660 12436 38712 12442
rect 38212 12306 38240 12406
rect 38660 12378 38712 12384
rect 40040 12436 40092 12442
rect 40040 12378 40092 12384
rect 38200 12300 38252 12306
rect 38200 12242 38252 12248
rect 38108 12164 38160 12170
rect 38108 12106 38160 12112
rect 38212 11762 38240 12242
rect 40224 12232 40276 12238
rect 40224 12174 40276 12180
rect 39120 12096 39172 12102
rect 39120 12038 39172 12044
rect 38200 11756 38252 11762
rect 38200 11698 38252 11704
rect 38660 11756 38712 11762
rect 38660 11698 38712 11704
rect 37464 11552 37516 11558
rect 37464 11494 37516 11500
rect 37924 11552 37976 11558
rect 37924 11494 37976 11500
rect 37188 11144 37240 11150
rect 37188 11086 37240 11092
rect 37280 11144 37332 11150
rect 37280 11086 37332 11092
rect 36820 11008 36872 11014
rect 36820 10950 36872 10956
rect 36360 10260 36412 10266
rect 36360 10202 36412 10208
rect 36372 9722 36400 10202
rect 36728 10056 36780 10062
rect 36728 9998 36780 10004
rect 36360 9716 36412 9722
rect 36360 9658 36412 9664
rect 36740 9586 36768 9998
rect 36832 9586 36860 10950
rect 37200 10690 37228 11086
rect 37292 10810 37320 11086
rect 37476 11082 37504 11494
rect 38672 11354 38700 11698
rect 38660 11348 38712 11354
rect 38660 11290 38712 11296
rect 37556 11280 37608 11286
rect 37556 11222 37608 11228
rect 37372 11076 37424 11082
rect 37372 11018 37424 11024
rect 37464 11076 37516 11082
rect 37464 11018 37516 11024
rect 37280 10804 37332 10810
rect 37280 10746 37332 10752
rect 37200 10662 37320 10690
rect 37292 10606 37320 10662
rect 37280 10600 37332 10606
rect 37280 10542 37332 10548
rect 37384 10146 37412 11018
rect 37568 10674 37596 11222
rect 39132 11150 39160 12038
rect 39264 11452 39572 11461
rect 39264 11450 39270 11452
rect 39326 11450 39350 11452
rect 39406 11450 39430 11452
rect 39486 11450 39510 11452
rect 39566 11450 39572 11452
rect 39326 11398 39328 11450
rect 39508 11398 39510 11450
rect 39264 11396 39270 11398
rect 39326 11396 39350 11398
rect 39406 11396 39430 11398
rect 39486 11396 39510 11398
rect 39566 11396 39572 11398
rect 39264 11387 39572 11396
rect 40236 11286 40264 12174
rect 40972 11830 41000 12582
rect 40960 11824 41012 11830
rect 40960 11766 41012 11772
rect 40684 11756 40736 11762
rect 40684 11698 40736 11704
rect 40224 11280 40276 11286
rect 40224 11222 40276 11228
rect 39120 11144 39172 11150
rect 39120 11086 39172 11092
rect 39764 11076 39816 11082
rect 39764 11018 39816 11024
rect 38108 11008 38160 11014
rect 38108 10950 38160 10956
rect 38120 10810 38148 10950
rect 38108 10804 38160 10810
rect 38108 10746 38160 10752
rect 37556 10668 37608 10674
rect 37556 10610 37608 10616
rect 37188 10124 37240 10130
rect 37188 10066 37240 10072
rect 37292 10118 37412 10146
rect 37556 10124 37608 10130
rect 36728 9580 36780 9586
rect 36728 9522 36780 9528
rect 36820 9580 36872 9586
rect 36820 9522 36872 9528
rect 36360 9512 36412 9518
rect 36360 9454 36412 9460
rect 36372 8498 36400 9454
rect 37004 9376 37056 9382
rect 37004 9318 37056 9324
rect 37016 8974 37044 9318
rect 37004 8968 37056 8974
rect 37004 8910 37056 8916
rect 36360 8492 36412 8498
rect 36360 8434 36412 8440
rect 36544 8424 36596 8430
rect 36544 8366 36596 8372
rect 36268 8356 36320 8362
rect 36268 8298 36320 8304
rect 36176 8288 36228 8294
rect 36176 8230 36228 8236
rect 36176 8016 36228 8022
rect 36082 7984 36138 7993
rect 36138 7964 36176 7970
rect 36138 7958 36228 7964
rect 36138 7942 36216 7958
rect 36082 7919 36138 7928
rect 36280 7750 36308 8298
rect 36452 8288 36504 8294
rect 36452 8230 36504 8236
rect 36464 8090 36492 8230
rect 36556 8090 36584 8366
rect 37016 8090 37044 8910
rect 36452 8084 36504 8090
rect 36452 8026 36504 8032
rect 36544 8084 36596 8090
rect 36544 8026 36596 8032
rect 37004 8084 37056 8090
rect 37004 8026 37056 8032
rect 36268 7744 36320 7750
rect 36268 7686 36320 7692
rect 35348 7404 35400 7410
rect 35992 7404 36044 7410
rect 35400 7364 35480 7392
rect 35348 7346 35400 7352
rect 35256 7336 35308 7342
rect 35256 7278 35308 7284
rect 35164 6860 35216 6866
rect 35164 6802 35216 6808
rect 35072 6384 35124 6390
rect 35072 6326 35124 6332
rect 34980 6112 35032 6118
rect 34980 6054 35032 6060
rect 34796 5646 34848 5652
rect 34886 5672 34942 5681
rect 34886 5607 34888 5616
rect 34940 5607 34942 5616
rect 34888 5578 34940 5584
rect 33790 5468 34098 5477
rect 33790 5466 33796 5468
rect 33852 5466 33876 5468
rect 33932 5466 33956 5468
rect 34012 5466 34036 5468
rect 34092 5466 34098 5468
rect 33852 5414 33854 5466
rect 34034 5414 34036 5466
rect 33790 5412 33796 5414
rect 33852 5412 33876 5414
rect 33932 5412 33956 5414
rect 34012 5412 34036 5414
rect 34092 5412 34098 5414
rect 33790 5403 34098 5412
rect 33416 5228 33468 5234
rect 33416 5170 33468 5176
rect 34992 5030 35020 6054
rect 35176 5914 35204 6802
rect 35348 6656 35400 6662
rect 35348 6598 35400 6604
rect 35360 6322 35388 6598
rect 35452 6322 35480 7364
rect 35992 7346 36044 7352
rect 36280 7342 36308 7686
rect 35624 7336 35676 7342
rect 35624 7278 35676 7284
rect 36268 7336 36320 7342
rect 36268 7278 36320 7284
rect 36728 7336 36780 7342
rect 36728 7278 36780 7284
rect 35636 6746 35664 7278
rect 36636 7200 36688 7206
rect 36636 7142 36688 7148
rect 36648 6798 36676 7142
rect 35808 6792 35860 6798
rect 35636 6740 35808 6746
rect 35636 6734 35860 6740
rect 36544 6792 36596 6798
rect 36544 6734 36596 6740
rect 36636 6792 36688 6798
rect 36636 6734 36688 6740
rect 35532 6724 35584 6730
rect 35532 6666 35584 6672
rect 35636 6718 35848 6734
rect 35992 6724 36044 6730
rect 35348 6316 35400 6322
rect 35348 6258 35400 6264
rect 35440 6316 35492 6322
rect 35440 6258 35492 6264
rect 35452 6118 35480 6258
rect 35348 6112 35400 6118
rect 35348 6054 35400 6060
rect 35440 6112 35492 6118
rect 35440 6054 35492 6060
rect 35164 5908 35216 5914
rect 35164 5850 35216 5856
rect 35176 5234 35204 5850
rect 35360 5642 35388 6054
rect 35544 5914 35572 6666
rect 35636 6186 35664 6718
rect 35992 6666 36044 6672
rect 36360 6724 36412 6730
rect 36412 6684 36492 6712
rect 36360 6666 36412 6672
rect 36004 6322 36032 6666
rect 36268 6656 36320 6662
rect 36268 6598 36320 6604
rect 36280 6390 36308 6598
rect 36464 6458 36492 6684
rect 36452 6452 36504 6458
rect 36452 6394 36504 6400
rect 36268 6384 36320 6390
rect 36268 6326 36320 6332
rect 35992 6316 36044 6322
rect 35992 6258 36044 6264
rect 35624 6180 35676 6186
rect 35624 6122 35676 6128
rect 36268 6112 36320 6118
rect 36268 6054 36320 6060
rect 35532 5908 35584 5914
rect 35532 5850 35584 5856
rect 35348 5636 35400 5642
rect 35348 5578 35400 5584
rect 35164 5228 35216 5234
rect 35164 5170 35216 5176
rect 35532 5228 35584 5234
rect 35532 5170 35584 5176
rect 34980 5024 35032 5030
rect 34980 4966 35032 4972
rect 35544 4826 35572 5170
rect 35532 4820 35584 4826
rect 35532 4762 35584 4768
rect 36280 4622 36308 6054
rect 36556 5914 36584 6734
rect 36544 5908 36596 5914
rect 36544 5850 36596 5856
rect 36740 5642 36768 7278
rect 37016 7002 37044 8026
rect 37200 7886 37228 10066
rect 37292 9042 37320 10118
rect 37556 10066 37608 10072
rect 37464 9580 37516 9586
rect 37464 9522 37516 9528
rect 37280 9036 37332 9042
rect 37280 8978 37332 8984
rect 37372 9036 37424 9042
rect 37372 8978 37424 8984
rect 37384 8945 37412 8978
rect 37370 8936 37426 8945
rect 37370 8871 37426 8880
rect 37476 8634 37504 9522
rect 37568 9518 37596 10066
rect 38120 10062 38148 10746
rect 39672 10736 39724 10742
rect 39672 10678 39724 10684
rect 39264 10364 39572 10373
rect 39264 10362 39270 10364
rect 39326 10362 39350 10364
rect 39406 10362 39430 10364
rect 39486 10362 39510 10364
rect 39566 10362 39572 10364
rect 39326 10310 39328 10362
rect 39508 10310 39510 10362
rect 39264 10308 39270 10310
rect 39326 10308 39350 10310
rect 39406 10308 39430 10310
rect 39486 10308 39510 10310
rect 39566 10308 39572 10310
rect 39264 10299 39572 10308
rect 37648 10056 37700 10062
rect 37648 9998 37700 10004
rect 38108 10056 38160 10062
rect 38108 9998 38160 10004
rect 37556 9512 37608 9518
rect 37556 9454 37608 9460
rect 37568 9382 37596 9454
rect 37660 9450 37688 9998
rect 39684 9722 39712 10678
rect 39776 10266 39804 11018
rect 40696 10674 40724 11698
rect 41064 11354 41092 12786
rect 41524 12306 41552 15982
rect 41616 14618 41644 16050
rect 44008 15570 44036 17478
rect 44737 17436 45045 17445
rect 44737 17434 44743 17436
rect 44799 17434 44823 17436
rect 44879 17434 44903 17436
rect 44959 17434 44983 17436
rect 45039 17434 45045 17436
rect 44799 17382 44801 17434
rect 44981 17382 44983 17434
rect 44737 17380 44743 17382
rect 44799 17380 44823 17382
rect 44879 17380 44903 17382
rect 44959 17380 44983 17382
rect 45039 17380 45045 17382
rect 44737 17371 45045 17380
rect 45112 16794 45140 19200
rect 45100 16788 45152 16794
rect 45100 16730 45152 16736
rect 44737 16348 45045 16357
rect 44737 16346 44743 16348
rect 44799 16346 44823 16348
rect 44879 16346 44903 16348
rect 44959 16346 44983 16348
rect 45039 16346 45045 16348
rect 44799 16294 44801 16346
rect 44981 16294 44983 16346
rect 44737 16292 44743 16294
rect 44799 16292 44823 16294
rect 44879 16292 44903 16294
rect 44959 16292 44983 16294
rect 45039 16292 45045 16294
rect 44737 16283 45045 16292
rect 44364 15904 44416 15910
rect 44364 15846 44416 15852
rect 44376 15745 44404 15846
rect 44362 15736 44418 15745
rect 44362 15671 44418 15680
rect 43996 15564 44048 15570
rect 43996 15506 44048 15512
rect 44737 15260 45045 15269
rect 44737 15258 44743 15260
rect 44799 15258 44823 15260
rect 44879 15258 44903 15260
rect 44959 15258 44983 15260
rect 45039 15258 45045 15260
rect 44799 15206 44801 15258
rect 44981 15206 44983 15258
rect 44737 15204 44743 15206
rect 44799 15204 44823 15206
rect 44879 15204 44903 15206
rect 44959 15204 44983 15206
rect 45039 15204 45045 15206
rect 44737 15195 45045 15204
rect 41604 14612 41656 14618
rect 41604 14554 41656 14560
rect 41696 14408 41748 14414
rect 41696 14350 41748 14356
rect 45006 14376 45062 14385
rect 41708 14006 41736 14350
rect 45006 14311 45008 14320
rect 45060 14311 45062 14320
rect 45008 14282 45060 14288
rect 44737 14172 45045 14181
rect 44737 14170 44743 14172
rect 44799 14170 44823 14172
rect 44879 14170 44903 14172
rect 44959 14170 44983 14172
rect 45039 14170 45045 14172
rect 44799 14118 44801 14170
rect 44981 14118 44983 14170
rect 44737 14116 44743 14118
rect 44799 14116 44823 14118
rect 44879 14116 44903 14118
rect 44959 14116 44983 14118
rect 45039 14116 45045 14118
rect 44737 14107 45045 14116
rect 41696 14000 41748 14006
rect 41694 13968 41696 13977
rect 41748 13968 41750 13977
rect 41694 13903 41750 13912
rect 41788 13864 41840 13870
rect 41788 13806 41840 13812
rect 41512 12300 41564 12306
rect 41512 12242 41564 12248
rect 41420 12232 41472 12238
rect 41420 12174 41472 12180
rect 41432 11354 41460 12174
rect 41800 11801 41828 13806
rect 41972 13796 42024 13802
rect 41972 13738 42024 13744
rect 41786 11792 41842 11801
rect 41786 11727 41842 11736
rect 41880 11552 41932 11558
rect 41880 11494 41932 11500
rect 41052 11348 41104 11354
rect 41052 11290 41104 11296
rect 41420 11348 41472 11354
rect 41420 11290 41472 11296
rect 41892 11218 41920 11494
rect 41984 11218 42012 13738
rect 44737 13084 45045 13093
rect 44737 13082 44743 13084
rect 44799 13082 44823 13084
rect 44879 13082 44903 13084
rect 44959 13082 44983 13084
rect 45039 13082 45045 13084
rect 44799 13030 44801 13082
rect 44981 13030 44983 13082
rect 44737 13028 44743 13030
rect 44799 13028 44823 13030
rect 44879 13028 44903 13030
rect 44959 13028 44983 13030
rect 45039 13028 45045 13030
rect 44737 13019 45045 13028
rect 45008 12640 45060 12646
rect 45008 12582 45060 12588
rect 45020 12345 45048 12582
rect 45006 12336 45062 12345
rect 45006 12271 45062 12280
rect 44737 11996 45045 12005
rect 44737 11994 44743 11996
rect 44799 11994 44823 11996
rect 44879 11994 44903 11996
rect 44959 11994 44983 11996
rect 45039 11994 45045 11996
rect 44799 11942 44801 11994
rect 44981 11942 44983 11994
rect 44737 11940 44743 11942
rect 44799 11940 44823 11942
rect 44879 11940 44903 11942
rect 44959 11940 44983 11942
rect 45039 11940 45045 11942
rect 44737 11931 45045 11940
rect 41880 11212 41932 11218
rect 41880 11154 41932 11160
rect 41972 11212 42024 11218
rect 41972 11154 42024 11160
rect 45008 11144 45060 11150
rect 45006 11112 45008 11121
rect 45060 11112 45062 11121
rect 41788 11076 41840 11082
rect 45006 11047 45062 11056
rect 41788 11018 41840 11024
rect 39948 10668 40000 10674
rect 39948 10610 40000 10616
rect 40684 10668 40736 10674
rect 40684 10610 40736 10616
rect 39856 10464 39908 10470
rect 39856 10406 39908 10412
rect 39764 10260 39816 10266
rect 39764 10202 39816 10208
rect 39672 9716 39724 9722
rect 39672 9658 39724 9664
rect 39776 9586 39804 10202
rect 39868 10130 39896 10406
rect 39960 10266 39988 10610
rect 40592 10532 40644 10538
rect 40592 10474 40644 10480
rect 40408 10464 40460 10470
rect 40408 10406 40460 10412
rect 39948 10260 40000 10266
rect 39948 10202 40000 10208
rect 40316 10260 40368 10266
rect 40316 10202 40368 10208
rect 39856 10124 39908 10130
rect 39856 10066 39908 10072
rect 40224 10056 40276 10062
rect 40224 9998 40276 10004
rect 40040 9920 40092 9926
rect 40040 9862 40092 9868
rect 39948 9716 40000 9722
rect 39948 9658 40000 9664
rect 39960 9586 39988 9658
rect 39764 9580 39816 9586
rect 39764 9522 39816 9528
rect 39948 9580 40000 9586
rect 39948 9522 40000 9528
rect 37648 9444 37700 9450
rect 37648 9386 37700 9392
rect 39672 9444 39724 9450
rect 39672 9386 39724 9392
rect 37556 9376 37608 9382
rect 37556 9318 37608 9324
rect 39264 9276 39572 9285
rect 39264 9274 39270 9276
rect 39326 9274 39350 9276
rect 39406 9274 39430 9276
rect 39486 9274 39510 9276
rect 39566 9274 39572 9276
rect 39326 9222 39328 9274
rect 39508 9222 39510 9274
rect 39264 9220 39270 9222
rect 39326 9220 39350 9222
rect 39406 9220 39430 9222
rect 39486 9220 39510 9222
rect 39566 9220 39572 9222
rect 39264 9211 39572 9220
rect 39396 8968 39448 8974
rect 39210 8936 39266 8945
rect 38936 8900 38988 8906
rect 39396 8910 39448 8916
rect 39210 8871 39212 8880
rect 38936 8842 38988 8848
rect 39264 8871 39266 8880
rect 39212 8842 39264 8848
rect 38476 8832 38528 8838
rect 38528 8780 38792 8786
rect 38476 8774 38792 8780
rect 38488 8758 38792 8774
rect 37464 8628 37516 8634
rect 37464 8570 37516 8576
rect 38764 8566 38792 8758
rect 37372 8560 37424 8566
rect 37372 8502 37424 8508
rect 38752 8560 38804 8566
rect 38752 8502 38804 8508
rect 37384 8090 37412 8502
rect 38568 8492 38620 8498
rect 38568 8434 38620 8440
rect 38474 8392 38530 8401
rect 38016 8356 38068 8362
rect 38474 8327 38530 8336
rect 38016 8298 38068 8304
rect 37372 8084 37424 8090
rect 37372 8026 37424 8032
rect 38028 7886 38056 8298
rect 37096 7880 37148 7886
rect 37096 7822 37148 7828
rect 37188 7880 37240 7886
rect 37188 7822 37240 7828
rect 38016 7880 38068 7886
rect 38016 7822 38068 7828
rect 37108 7546 37136 7822
rect 37188 7744 37240 7750
rect 37188 7686 37240 7692
rect 37096 7540 37148 7546
rect 37096 7482 37148 7488
rect 37200 7342 37228 7686
rect 38488 7426 38516 8327
rect 38580 7546 38608 8434
rect 38660 8288 38712 8294
rect 38660 8230 38712 8236
rect 38672 7954 38700 8230
rect 38660 7948 38712 7954
rect 38660 7890 38712 7896
rect 38764 7886 38792 8502
rect 38752 7880 38804 7886
rect 38752 7822 38804 7828
rect 38568 7540 38620 7546
rect 38568 7482 38620 7488
rect 38488 7398 38608 7426
rect 37188 7336 37240 7342
rect 37188 7278 37240 7284
rect 37004 6996 37056 7002
rect 37004 6938 37056 6944
rect 36910 6896 36966 6905
rect 36910 6831 36966 6840
rect 36924 6798 36952 6831
rect 36912 6792 36964 6798
rect 36912 6734 36964 6740
rect 37372 6656 37424 6662
rect 37372 6598 37424 6604
rect 37648 6656 37700 6662
rect 37648 6598 37700 6604
rect 37384 6322 37412 6598
rect 37556 6452 37608 6458
rect 37556 6394 37608 6400
rect 37372 6316 37424 6322
rect 37372 6258 37424 6264
rect 37280 6248 37332 6254
rect 37280 6190 37332 6196
rect 36912 6112 36964 6118
rect 36912 6054 36964 6060
rect 37094 6080 37150 6089
rect 36924 5681 36952 6054
rect 37094 6015 37150 6024
rect 36910 5672 36966 5681
rect 36728 5636 36780 5642
rect 36910 5607 36912 5616
rect 36728 5578 36780 5584
rect 36964 5607 36966 5616
rect 36912 5578 36964 5584
rect 36740 4622 36768 5578
rect 37108 5574 37136 6015
rect 37292 5914 37320 6190
rect 37188 5908 37240 5914
rect 37188 5850 37240 5856
rect 37280 5908 37332 5914
rect 37280 5850 37332 5856
rect 37096 5568 37148 5574
rect 37096 5510 37148 5516
rect 37200 5234 37228 5850
rect 37384 5642 37412 6258
rect 37372 5636 37424 5642
rect 37372 5578 37424 5584
rect 37568 5302 37596 6394
rect 37660 6322 37688 6598
rect 37648 6316 37700 6322
rect 37648 6258 37700 6264
rect 37660 5778 37688 6258
rect 38580 6186 38608 7398
rect 38660 6316 38712 6322
rect 38660 6258 38712 6264
rect 38568 6180 38620 6186
rect 38568 6122 38620 6128
rect 37648 5772 37700 5778
rect 37648 5714 37700 5720
rect 38580 5710 38608 6122
rect 38672 5710 38700 6258
rect 38752 6112 38804 6118
rect 38752 6054 38804 6060
rect 38016 5704 38068 5710
rect 38016 5646 38068 5652
rect 38568 5704 38620 5710
rect 38568 5646 38620 5652
rect 38660 5704 38712 5710
rect 38660 5646 38712 5652
rect 37556 5296 37608 5302
rect 37556 5238 37608 5244
rect 37188 5228 37240 5234
rect 37188 5170 37240 5176
rect 37200 5030 37228 5170
rect 37188 5024 37240 5030
rect 37188 4966 37240 4972
rect 37200 4690 37228 4966
rect 38028 4826 38056 5646
rect 38660 5568 38712 5574
rect 38660 5510 38712 5516
rect 38672 5302 38700 5510
rect 38764 5302 38792 6054
rect 38660 5296 38712 5302
rect 38660 5238 38712 5244
rect 38752 5296 38804 5302
rect 38752 5238 38804 5244
rect 38568 5160 38620 5166
rect 38568 5102 38620 5108
rect 38580 4826 38608 5102
rect 38948 5098 38976 8842
rect 39408 8634 39436 8910
rect 39684 8838 39712 9386
rect 39776 8974 39804 9522
rect 40052 9450 40080 9862
rect 40132 9512 40184 9518
rect 40132 9454 40184 9460
rect 40040 9444 40092 9450
rect 40040 9386 40092 9392
rect 39856 9104 39908 9110
rect 39856 9046 39908 9052
rect 39764 8968 39816 8974
rect 39764 8910 39816 8916
rect 39672 8832 39724 8838
rect 39672 8774 39724 8780
rect 39396 8628 39448 8634
rect 39396 8570 39448 8576
rect 39776 8498 39804 8910
rect 39868 8650 39896 9046
rect 40052 8974 40080 9386
rect 40040 8968 40092 8974
rect 40040 8910 40092 8916
rect 39868 8622 39988 8650
rect 39960 8498 39988 8622
rect 40144 8566 40172 9454
rect 40236 9178 40264 9998
rect 40224 9172 40276 9178
rect 40224 9114 40276 9120
rect 40328 8974 40356 10202
rect 40420 10062 40448 10406
rect 40500 10192 40552 10198
rect 40500 10134 40552 10140
rect 40512 10062 40540 10134
rect 40408 10056 40460 10062
rect 40408 9998 40460 10004
rect 40500 10056 40552 10062
rect 40500 9998 40552 10004
rect 40512 9926 40540 9998
rect 40500 9920 40552 9926
rect 40500 9862 40552 9868
rect 40512 9722 40540 9862
rect 40500 9716 40552 9722
rect 40500 9658 40552 9664
rect 40408 9580 40460 9586
rect 40408 9522 40460 9528
rect 40316 8968 40368 8974
rect 40314 8936 40316 8945
rect 40368 8936 40370 8945
rect 40314 8871 40370 8880
rect 40132 8560 40184 8566
rect 40132 8502 40184 8508
rect 39764 8492 39816 8498
rect 39764 8434 39816 8440
rect 39948 8492 40000 8498
rect 39948 8434 40000 8440
rect 39264 8188 39572 8197
rect 39264 8186 39270 8188
rect 39326 8186 39350 8188
rect 39406 8186 39430 8188
rect 39486 8186 39510 8188
rect 39566 8186 39572 8188
rect 39326 8134 39328 8186
rect 39508 8134 39510 8186
rect 39264 8132 39270 8134
rect 39326 8132 39350 8134
rect 39406 8132 39430 8134
rect 39486 8132 39510 8134
rect 39566 8132 39572 8134
rect 39264 8123 39572 8132
rect 39396 8084 39448 8090
rect 39396 8026 39448 8032
rect 39304 7880 39356 7886
rect 39304 7822 39356 7828
rect 39316 7546 39344 7822
rect 39304 7540 39356 7546
rect 39304 7482 39356 7488
rect 39408 7342 39436 8026
rect 39580 7812 39632 7818
rect 39580 7754 39632 7760
rect 39592 7546 39620 7754
rect 39580 7540 39632 7546
rect 39580 7482 39632 7488
rect 39776 7342 39804 8434
rect 39396 7336 39448 7342
rect 39396 7278 39448 7284
rect 39764 7336 39816 7342
rect 39764 7278 39816 7284
rect 39264 7100 39572 7109
rect 39264 7098 39270 7100
rect 39326 7098 39350 7100
rect 39406 7098 39430 7100
rect 39486 7098 39510 7100
rect 39566 7098 39572 7100
rect 39326 7046 39328 7098
rect 39508 7046 39510 7098
rect 39264 7044 39270 7046
rect 39326 7044 39350 7046
rect 39406 7044 39430 7046
rect 39486 7044 39510 7046
rect 39566 7044 39572 7046
rect 39264 7035 39572 7044
rect 39776 6934 39804 7278
rect 40328 7274 40356 8871
rect 40420 8294 40448 9522
rect 40604 9518 40632 10474
rect 40696 10130 40724 10610
rect 40684 10124 40736 10130
rect 40684 10066 40736 10072
rect 40960 9920 41012 9926
rect 40960 9862 41012 9868
rect 40592 9512 40644 9518
rect 40592 9454 40644 9460
rect 40500 8968 40552 8974
rect 40500 8910 40552 8916
rect 40408 8288 40460 8294
rect 40408 8230 40460 8236
rect 40512 7954 40540 8910
rect 40684 8628 40736 8634
rect 40684 8570 40736 8576
rect 40500 7948 40552 7954
rect 40500 7890 40552 7896
rect 40224 7268 40276 7274
rect 40224 7210 40276 7216
rect 40316 7268 40368 7274
rect 40316 7210 40368 7216
rect 40132 7200 40184 7206
rect 40132 7142 40184 7148
rect 39764 6928 39816 6934
rect 39764 6870 39816 6876
rect 40144 6798 40172 7142
rect 40236 7002 40264 7210
rect 40224 6996 40276 7002
rect 40224 6938 40276 6944
rect 40236 6798 40264 6938
rect 40132 6792 40184 6798
rect 40132 6734 40184 6740
rect 40224 6792 40276 6798
rect 40224 6734 40276 6740
rect 39028 6316 39080 6322
rect 39028 6258 39080 6264
rect 39040 5778 39068 6258
rect 39264 6012 39572 6021
rect 39264 6010 39270 6012
rect 39326 6010 39350 6012
rect 39406 6010 39430 6012
rect 39486 6010 39510 6012
rect 39566 6010 39572 6012
rect 39326 5958 39328 6010
rect 39508 5958 39510 6010
rect 39264 5956 39270 5958
rect 39326 5956 39350 5958
rect 39406 5956 39430 5958
rect 39486 5956 39510 5958
rect 39566 5956 39572 5958
rect 39264 5947 39572 5956
rect 40328 5914 40356 7210
rect 40512 6882 40540 7890
rect 40420 6866 40540 6882
rect 40408 6860 40540 6866
rect 40460 6854 40540 6860
rect 40408 6802 40460 6808
rect 40696 6798 40724 8570
rect 40972 8498 41000 9862
rect 41604 9580 41656 9586
rect 41604 9522 41656 9528
rect 41052 9512 41104 9518
rect 41052 9454 41104 9460
rect 41064 8838 41092 9454
rect 41328 9376 41380 9382
rect 41328 9318 41380 9324
rect 41052 8832 41104 8838
rect 41052 8774 41104 8780
rect 40960 8492 41012 8498
rect 40960 8434 41012 8440
rect 41064 8430 41092 8774
rect 41340 8498 41368 9318
rect 41616 9178 41644 9522
rect 41800 9450 41828 11018
rect 44737 10908 45045 10917
rect 44737 10906 44743 10908
rect 44799 10906 44823 10908
rect 44879 10906 44903 10908
rect 44959 10906 44983 10908
rect 45039 10906 45045 10908
rect 44799 10854 44801 10906
rect 44981 10854 44983 10906
rect 44737 10852 44743 10854
rect 44799 10852 44823 10854
rect 44879 10852 44903 10854
rect 44959 10852 44983 10854
rect 45039 10852 45045 10854
rect 44737 10843 45045 10852
rect 42800 10668 42852 10674
rect 42800 10610 42852 10616
rect 42812 10266 42840 10610
rect 42800 10260 42852 10266
rect 42800 10202 42852 10208
rect 42892 10056 42944 10062
rect 42892 9998 42944 10004
rect 42904 9654 42932 9998
rect 44737 9820 45045 9829
rect 44737 9818 44743 9820
rect 44799 9818 44823 9820
rect 44879 9818 44903 9820
rect 44959 9818 44983 9820
rect 45039 9818 45045 9820
rect 44799 9766 44801 9818
rect 44981 9766 44983 9818
rect 44737 9764 44743 9766
rect 44799 9764 44823 9766
rect 44879 9764 44903 9766
rect 44959 9764 44983 9766
rect 45039 9764 45045 9766
rect 44737 9755 45045 9764
rect 42892 9648 42944 9654
rect 42892 9590 42944 9596
rect 42616 9580 42668 9586
rect 42616 9522 42668 9528
rect 42708 9580 42760 9586
rect 42708 9522 42760 9528
rect 41972 9512 42024 9518
rect 41972 9454 42024 9460
rect 41788 9444 41840 9450
rect 41788 9386 41840 9392
rect 41604 9172 41656 9178
rect 41604 9114 41656 9120
rect 41696 8628 41748 8634
rect 41696 8570 41748 8576
rect 41708 8498 41736 8570
rect 41328 8492 41380 8498
rect 41328 8434 41380 8440
rect 41696 8492 41748 8498
rect 41696 8434 41748 8440
rect 41052 8424 41104 8430
rect 41052 8366 41104 8372
rect 41052 8288 41104 8294
rect 41052 8230 41104 8236
rect 41064 7886 41092 8230
rect 41052 7880 41104 7886
rect 41052 7822 41104 7828
rect 41064 7392 41092 7822
rect 41420 7812 41472 7818
rect 41420 7754 41472 7760
rect 41432 7546 41460 7754
rect 41604 7744 41656 7750
rect 41604 7686 41656 7692
rect 41420 7540 41472 7546
rect 41420 7482 41472 7488
rect 41616 7410 41644 7686
rect 40972 7364 41092 7392
rect 41604 7404 41656 7410
rect 40776 7336 40828 7342
rect 40776 7278 40828 7284
rect 40868 7336 40920 7342
rect 40868 7278 40920 7284
rect 40788 7002 40816 7278
rect 40776 6996 40828 7002
rect 40776 6938 40828 6944
rect 40880 6934 40908 7278
rect 40868 6928 40920 6934
rect 40868 6870 40920 6876
rect 40500 6792 40552 6798
rect 40500 6734 40552 6740
rect 40684 6792 40736 6798
rect 40684 6734 40736 6740
rect 40776 6792 40828 6798
rect 40776 6734 40828 6740
rect 40316 5908 40368 5914
rect 40316 5850 40368 5856
rect 40512 5846 40540 6734
rect 40696 6254 40724 6734
rect 40684 6248 40736 6254
rect 40684 6190 40736 6196
rect 40500 5840 40552 5846
rect 40500 5782 40552 5788
rect 40788 5778 40816 6734
rect 40972 6254 41000 7364
rect 41604 7346 41656 7352
rect 41420 7336 41472 7342
rect 41420 7278 41472 7284
rect 41432 6662 41460 7278
rect 41420 6656 41472 6662
rect 41420 6598 41472 6604
rect 41512 6316 41564 6322
rect 41512 6258 41564 6264
rect 40960 6248 41012 6254
rect 40960 6190 41012 6196
rect 41524 6186 41552 6258
rect 41984 6225 42012 9454
rect 42628 9382 42656 9522
rect 42616 9376 42668 9382
rect 42616 9318 42668 9324
rect 42720 8838 42748 9522
rect 44180 9444 44232 9450
rect 44180 9386 44232 9392
rect 42892 9376 42944 9382
rect 42892 9318 42944 9324
rect 42800 8900 42852 8906
rect 42800 8842 42852 8848
rect 42708 8832 42760 8838
rect 42708 8774 42760 8780
rect 42720 8634 42748 8774
rect 42708 8628 42760 8634
rect 42708 8570 42760 8576
rect 42812 8090 42840 8842
rect 42904 8634 42932 9318
rect 44192 8634 44220 9386
rect 44362 8936 44418 8945
rect 44362 8871 44418 8880
rect 42892 8628 42944 8634
rect 42892 8570 42944 8576
rect 44180 8628 44232 8634
rect 44180 8570 44232 8576
rect 44376 8498 44404 8871
rect 44737 8732 45045 8741
rect 44737 8730 44743 8732
rect 44799 8730 44823 8732
rect 44879 8730 44903 8732
rect 44959 8730 44983 8732
rect 45039 8730 45045 8732
rect 44799 8678 44801 8730
rect 44981 8678 44983 8730
rect 44737 8676 44743 8678
rect 44799 8676 44823 8678
rect 44879 8676 44903 8678
rect 44959 8676 44983 8678
rect 45039 8676 45045 8678
rect 44737 8667 45045 8676
rect 44364 8492 44416 8498
rect 44364 8434 44416 8440
rect 43168 8288 43220 8294
rect 43168 8230 43220 8236
rect 42800 8084 42852 8090
rect 42800 8026 42852 8032
rect 43180 7886 43208 8230
rect 43168 7880 43220 7886
rect 44364 7880 44416 7886
rect 43168 7822 43220 7828
rect 44362 7848 44364 7857
rect 44416 7848 44418 7857
rect 44362 7783 44418 7792
rect 43444 7744 43496 7750
rect 43444 7686 43496 7692
rect 43456 6866 43484 7686
rect 44737 7644 45045 7653
rect 44737 7642 44743 7644
rect 44799 7642 44823 7644
rect 44879 7642 44903 7644
rect 44959 7642 44983 7644
rect 45039 7642 45045 7644
rect 44799 7590 44801 7642
rect 44981 7590 44983 7642
rect 44737 7588 44743 7590
rect 44799 7588 44823 7590
rect 44879 7588 44903 7590
rect 44959 7588 44983 7590
rect 45039 7588 45045 7590
rect 44737 7579 45045 7588
rect 43444 6860 43496 6866
rect 43444 6802 43496 6808
rect 43720 6656 43772 6662
rect 43720 6598 43772 6604
rect 43732 6458 43760 6598
rect 44737 6556 45045 6565
rect 44737 6554 44743 6556
rect 44799 6554 44823 6556
rect 44879 6554 44903 6556
rect 44959 6554 44983 6556
rect 45039 6554 45045 6556
rect 44799 6502 44801 6554
rect 44981 6502 44983 6554
rect 44737 6500 44743 6502
rect 44799 6500 44823 6502
rect 44879 6500 44903 6502
rect 44959 6500 44983 6502
rect 45039 6500 45045 6502
rect 44737 6491 45045 6500
rect 43720 6452 43772 6458
rect 43720 6394 43772 6400
rect 41970 6216 42026 6225
rect 41512 6180 41564 6186
rect 41970 6151 42026 6160
rect 41512 6122 41564 6128
rect 39028 5772 39080 5778
rect 39028 5714 39080 5720
rect 40776 5772 40828 5778
rect 40776 5714 40828 5720
rect 41524 5370 41552 6122
rect 42616 6112 42668 6118
rect 42616 6054 42668 6060
rect 42628 5710 42656 6054
rect 42616 5704 42668 5710
rect 42616 5646 42668 5652
rect 43904 5636 43956 5642
rect 43904 5578 43956 5584
rect 41696 5568 41748 5574
rect 41696 5510 41748 5516
rect 41512 5364 41564 5370
rect 41512 5306 41564 5312
rect 41418 5264 41474 5273
rect 41708 5234 41736 5510
rect 41418 5199 41420 5208
rect 41472 5199 41474 5208
rect 41696 5228 41748 5234
rect 41420 5170 41472 5176
rect 41696 5170 41748 5176
rect 42800 5228 42852 5234
rect 42800 5170 42852 5176
rect 42812 5137 42840 5170
rect 42798 5128 42854 5137
rect 38936 5092 38988 5098
rect 42798 5063 42854 5072
rect 38936 5034 38988 5040
rect 39264 4924 39572 4933
rect 39264 4922 39270 4924
rect 39326 4922 39350 4924
rect 39406 4922 39430 4924
rect 39486 4922 39510 4924
rect 39566 4922 39572 4924
rect 39326 4870 39328 4922
rect 39508 4870 39510 4922
rect 39264 4868 39270 4870
rect 39326 4868 39350 4870
rect 39406 4868 39430 4870
rect 39486 4868 39510 4870
rect 39566 4868 39572 4870
rect 39264 4859 39572 4868
rect 38016 4820 38068 4826
rect 38016 4762 38068 4768
rect 38568 4820 38620 4826
rect 38568 4762 38620 4768
rect 37188 4684 37240 4690
rect 37188 4626 37240 4632
rect 36268 4616 36320 4622
rect 36268 4558 36320 4564
rect 36728 4616 36780 4622
rect 36728 4558 36780 4564
rect 37464 4616 37516 4622
rect 37464 4558 37516 4564
rect 33790 4380 34098 4389
rect 33790 4378 33796 4380
rect 33852 4378 33876 4380
rect 33932 4378 33956 4380
rect 34012 4378 34036 4380
rect 34092 4378 34098 4380
rect 33852 4326 33854 4378
rect 34034 4326 34036 4378
rect 33790 4324 33796 4326
rect 33852 4324 33876 4326
rect 33932 4324 33956 4326
rect 34012 4324 34036 4326
rect 34092 4324 34098 4326
rect 33790 4315 34098 4324
rect 33508 3460 33560 3466
rect 33508 3402 33560 3408
rect 32496 2644 32548 2650
rect 32496 2586 32548 2592
rect 32220 2372 32272 2378
rect 32220 2314 32272 2320
rect 30656 2304 30708 2310
rect 30656 2246 30708 2252
rect 30300 870 30420 898
rect 30300 800 30328 870
rect 32232 800 32260 2314
rect 33520 800 33548 3402
rect 33790 3292 34098 3301
rect 33790 3290 33796 3292
rect 33852 3290 33876 3292
rect 33932 3290 33956 3292
rect 34012 3290 34036 3292
rect 34092 3290 34098 3292
rect 33852 3238 33854 3290
rect 34034 3238 34036 3290
rect 33790 3236 33796 3238
rect 33852 3236 33876 3238
rect 33932 3236 33956 3238
rect 34012 3236 34036 3238
rect 34092 3236 34098 3238
rect 33790 3227 34098 3236
rect 35440 2984 35492 2990
rect 35440 2926 35492 2932
rect 33790 2204 34098 2213
rect 33790 2202 33796 2204
rect 33852 2202 33876 2204
rect 33932 2202 33956 2204
rect 34012 2202 34036 2204
rect 34092 2202 34098 2204
rect 33852 2150 33854 2202
rect 34034 2150 34036 2202
rect 33790 2148 33796 2150
rect 33852 2148 33876 2150
rect 33932 2148 33956 2150
rect 34012 2148 34036 2150
rect 34092 2148 34098 2150
rect 33790 2139 34098 2148
rect 35452 800 35480 2926
rect 37476 2650 37504 4558
rect 41420 4072 41472 4078
rect 41420 4014 41472 4020
rect 39264 3836 39572 3845
rect 39264 3834 39270 3836
rect 39326 3834 39350 3836
rect 39406 3834 39430 3836
rect 39486 3834 39510 3836
rect 39566 3834 39572 3836
rect 39326 3782 39328 3834
rect 39508 3782 39510 3834
rect 39264 3780 39270 3782
rect 39326 3780 39350 3782
rect 39406 3780 39430 3782
rect 39486 3780 39510 3782
rect 39566 3780 39572 3782
rect 39264 3771 39572 3780
rect 39264 2748 39572 2757
rect 39264 2746 39270 2748
rect 39326 2746 39350 2748
rect 39406 2746 39430 2748
rect 39486 2746 39510 2748
rect 39566 2746 39572 2748
rect 39326 2694 39328 2746
rect 39508 2694 39510 2746
rect 39264 2692 39270 2694
rect 39326 2692 39350 2694
rect 39406 2692 39430 2694
rect 39486 2692 39510 2694
rect 39566 2692 39572 2694
rect 39264 2683 39572 2692
rect 37464 2644 37516 2650
rect 37464 2586 37516 2592
rect 37648 2440 37700 2446
rect 37648 2382 37700 2388
rect 38660 2440 38712 2446
rect 38660 2382 38712 2388
rect 40040 2440 40092 2446
rect 41432 2417 41460 4014
rect 43916 2650 43944 5578
rect 44737 5468 45045 5477
rect 44737 5466 44743 5468
rect 44799 5466 44823 5468
rect 44879 5466 44903 5468
rect 44959 5466 44983 5468
rect 45039 5466 45045 5468
rect 44799 5414 44801 5466
rect 44981 5414 44983 5466
rect 44737 5412 44743 5414
rect 44799 5412 44823 5414
rect 44879 5412 44903 5414
rect 44959 5412 44983 5414
rect 45039 5412 45045 5414
rect 44737 5403 45045 5412
rect 44640 5160 44692 5166
rect 44640 5102 44692 5108
rect 44180 4684 44232 4690
rect 44180 4626 44232 4632
rect 44192 3194 44220 4626
rect 44652 4185 44680 5102
rect 44737 4380 45045 4389
rect 44737 4378 44743 4380
rect 44799 4378 44823 4380
rect 44879 4378 44903 4380
rect 44959 4378 44983 4380
rect 45039 4378 45045 4380
rect 44799 4326 44801 4378
rect 44981 4326 44983 4378
rect 44737 4324 44743 4326
rect 44799 4324 44823 4326
rect 44879 4324 44903 4326
rect 44959 4324 44983 4326
rect 45039 4324 45045 4326
rect 44737 4315 45045 4324
rect 44638 4176 44694 4185
rect 44638 4111 44694 4120
rect 44640 3528 44692 3534
rect 44640 3470 44692 3476
rect 44180 3188 44232 3194
rect 44180 3130 44232 3136
rect 43904 2644 43956 2650
rect 43904 2586 43956 2592
rect 43812 2440 43864 2446
rect 40040 2382 40092 2388
rect 41418 2408 41474 2417
rect 37660 950 37688 2382
rect 36728 944 36780 950
rect 36728 886 36780 892
rect 37648 944 37700 950
rect 37648 886 37700 892
rect 36740 800 36768 886
rect 38672 800 38700 2382
rect 40052 898 40080 2382
rect 43812 2382 43864 2388
rect 41418 2343 41474 2352
rect 41880 2372 41932 2378
rect 41880 2314 41932 2320
rect 39960 870 40080 898
rect 39960 800 39988 870
rect 41892 800 41920 2314
rect 43824 800 43852 2382
rect -10 0 102 800
rect 1278 0 1390 800
rect 3210 0 3322 800
rect 4498 0 4610 800
rect 6430 0 6542 800
rect 7718 0 7830 800
rect 9650 0 9762 800
rect 10938 0 11050 800
rect 12870 0 12982 800
rect 14158 0 14270 800
rect 16090 0 16202 800
rect 17378 0 17490 800
rect 19310 0 19422 800
rect 20598 0 20710 800
rect 22530 0 22642 800
rect 23818 0 23930 800
rect 25750 0 25862 800
rect 27038 0 27150 800
rect 28970 0 29082 800
rect 30258 0 30370 800
rect 32190 0 32302 800
rect 33478 0 33590 800
rect 35410 0 35522 800
rect 36698 0 36810 800
rect 38630 0 38742 800
rect 39918 0 40030 800
rect 41850 0 41962 800
rect 43782 0 43894 800
rect 44652 785 44680 3470
rect 44737 3292 45045 3301
rect 44737 3290 44743 3292
rect 44799 3290 44823 3292
rect 44879 3290 44903 3292
rect 44959 3290 44983 3292
rect 45039 3290 45045 3292
rect 44799 3238 44801 3290
rect 44981 3238 44983 3290
rect 44737 3236 44743 3238
rect 44799 3236 44823 3238
rect 44879 3236 44903 3238
rect 44959 3236 44983 3238
rect 45039 3236 45045 3238
rect 44737 3227 45045 3236
rect 45100 3052 45152 3058
rect 45100 2994 45152 3000
rect 44737 2204 45045 2213
rect 44737 2202 44743 2204
rect 44799 2202 44823 2204
rect 44879 2202 44903 2204
rect 44959 2202 44983 2204
rect 45039 2202 45045 2204
rect 44799 2150 44801 2202
rect 44981 2150 44983 2202
rect 44737 2148 44743 2150
rect 44799 2148 44823 2150
rect 44879 2148 44903 2150
rect 44959 2148 44983 2150
rect 45039 2148 45045 2150
rect 44737 2139 45045 2148
rect 45112 800 45140 2994
rect 44638 776 44694 785
rect 44638 711 44694 720
rect 45070 0 45182 800
<< via2 >>
rect 1030 18400 1086 18456
rect 938 17040 994 17096
rect 11902 17434 11958 17436
rect 11982 17434 12038 17436
rect 12062 17434 12118 17436
rect 12142 17434 12198 17436
rect 11902 17382 11948 17434
rect 11948 17382 11958 17434
rect 11982 17382 12012 17434
rect 12012 17382 12024 17434
rect 12024 17382 12038 17434
rect 12062 17382 12076 17434
rect 12076 17382 12088 17434
rect 12088 17382 12118 17434
rect 12142 17382 12152 17434
rect 12152 17382 12198 17434
rect 11902 17380 11958 17382
rect 11982 17380 12038 17382
rect 12062 17380 12118 17382
rect 12142 17380 12198 17382
rect 1030 15000 1086 15056
rect 938 13640 994 13696
rect 938 10240 994 10296
rect 2134 12144 2190 12200
rect 1766 9424 1822 9480
rect 938 8200 994 8256
rect 6429 16890 6485 16892
rect 6509 16890 6565 16892
rect 6589 16890 6645 16892
rect 6669 16890 6725 16892
rect 6429 16838 6475 16890
rect 6475 16838 6485 16890
rect 6509 16838 6539 16890
rect 6539 16838 6551 16890
rect 6551 16838 6565 16890
rect 6589 16838 6603 16890
rect 6603 16838 6615 16890
rect 6615 16838 6645 16890
rect 6669 16838 6679 16890
rect 6679 16838 6725 16890
rect 6429 16836 6485 16838
rect 6509 16836 6565 16838
rect 6589 16836 6645 16838
rect 6669 16836 6725 16838
rect 4066 11600 4122 11656
rect 6429 15802 6485 15804
rect 6509 15802 6565 15804
rect 6589 15802 6645 15804
rect 6669 15802 6725 15804
rect 6429 15750 6475 15802
rect 6475 15750 6485 15802
rect 6509 15750 6539 15802
rect 6539 15750 6551 15802
rect 6551 15750 6565 15802
rect 6589 15750 6603 15802
rect 6603 15750 6615 15802
rect 6615 15750 6645 15802
rect 6669 15750 6679 15802
rect 6679 15750 6725 15802
rect 6429 15748 6485 15750
rect 6509 15748 6565 15750
rect 6589 15748 6645 15750
rect 6669 15748 6725 15750
rect 6429 14714 6485 14716
rect 6509 14714 6565 14716
rect 6589 14714 6645 14716
rect 6669 14714 6725 14716
rect 6429 14662 6475 14714
rect 6475 14662 6485 14714
rect 6509 14662 6539 14714
rect 6539 14662 6551 14714
rect 6551 14662 6565 14714
rect 6589 14662 6603 14714
rect 6603 14662 6615 14714
rect 6615 14662 6645 14714
rect 6669 14662 6679 14714
rect 6679 14662 6725 14714
rect 6429 14660 6485 14662
rect 6509 14660 6565 14662
rect 6589 14660 6645 14662
rect 6669 14660 6725 14662
rect 6429 13626 6485 13628
rect 6509 13626 6565 13628
rect 6589 13626 6645 13628
rect 6669 13626 6725 13628
rect 6429 13574 6475 13626
rect 6475 13574 6485 13626
rect 6509 13574 6539 13626
rect 6539 13574 6551 13626
rect 6551 13574 6565 13626
rect 6589 13574 6603 13626
rect 6603 13574 6615 13626
rect 6615 13574 6645 13626
rect 6669 13574 6679 13626
rect 6679 13574 6725 13626
rect 6429 13572 6485 13574
rect 6509 13572 6565 13574
rect 6589 13572 6645 13574
rect 6669 13572 6725 13574
rect 6429 12538 6485 12540
rect 6509 12538 6565 12540
rect 6589 12538 6645 12540
rect 6669 12538 6725 12540
rect 6429 12486 6475 12538
rect 6475 12486 6485 12538
rect 6509 12486 6539 12538
rect 6539 12486 6551 12538
rect 6551 12486 6565 12538
rect 6589 12486 6603 12538
rect 6603 12486 6615 12538
rect 6615 12486 6645 12538
rect 6669 12486 6679 12538
rect 6679 12486 6725 12538
rect 6429 12484 6485 12486
rect 6509 12484 6565 12486
rect 6589 12484 6645 12486
rect 6669 12484 6725 12486
rect 6918 11756 6974 11792
rect 6918 11736 6920 11756
rect 6920 11736 6972 11756
rect 6972 11736 6974 11756
rect 6429 11450 6485 11452
rect 6509 11450 6565 11452
rect 6589 11450 6645 11452
rect 6669 11450 6725 11452
rect 6429 11398 6475 11450
rect 6475 11398 6485 11450
rect 6509 11398 6539 11450
rect 6539 11398 6551 11450
rect 6551 11398 6565 11450
rect 6589 11398 6603 11450
rect 6603 11398 6615 11450
rect 6615 11398 6645 11450
rect 6669 11398 6679 11450
rect 6679 11398 6725 11450
rect 6429 11396 6485 11398
rect 6509 11396 6565 11398
rect 6589 11396 6645 11398
rect 6669 11396 6725 11398
rect 5354 10668 5410 10704
rect 5354 10648 5356 10668
rect 5356 10648 5408 10668
rect 5408 10648 5410 10668
rect 3606 8472 3662 8528
rect 938 6840 994 6896
rect 6429 10362 6485 10364
rect 6509 10362 6565 10364
rect 6589 10362 6645 10364
rect 6669 10362 6725 10364
rect 6429 10310 6475 10362
rect 6475 10310 6485 10362
rect 6509 10310 6539 10362
rect 6539 10310 6551 10362
rect 6551 10310 6565 10362
rect 6589 10310 6603 10362
rect 6603 10310 6615 10362
rect 6615 10310 6645 10362
rect 6669 10310 6679 10362
rect 6679 10310 6725 10362
rect 6429 10308 6485 10310
rect 6509 10308 6565 10310
rect 6589 10308 6645 10310
rect 6669 10308 6725 10310
rect 938 4800 994 4856
rect 6429 9274 6485 9276
rect 6509 9274 6565 9276
rect 6589 9274 6645 9276
rect 6669 9274 6725 9276
rect 6429 9222 6475 9274
rect 6475 9222 6485 9274
rect 6509 9222 6539 9274
rect 6539 9222 6551 9274
rect 6551 9222 6565 9274
rect 6589 9222 6603 9274
rect 6603 9222 6615 9274
rect 6615 9222 6645 9274
rect 6669 9222 6679 9274
rect 6679 9222 6725 9274
rect 6429 9220 6485 9222
rect 6509 9220 6565 9222
rect 6589 9220 6645 9222
rect 6669 9220 6725 9222
rect 11902 16346 11958 16348
rect 11982 16346 12038 16348
rect 12062 16346 12118 16348
rect 12142 16346 12198 16348
rect 11902 16294 11948 16346
rect 11948 16294 11958 16346
rect 11982 16294 12012 16346
rect 12012 16294 12024 16346
rect 12024 16294 12038 16346
rect 12062 16294 12076 16346
rect 12076 16294 12088 16346
rect 12088 16294 12118 16346
rect 12142 16294 12152 16346
rect 12152 16294 12198 16346
rect 11902 16292 11958 16294
rect 11982 16292 12038 16294
rect 12062 16292 12118 16294
rect 12142 16292 12198 16294
rect 11902 15258 11958 15260
rect 11982 15258 12038 15260
rect 12062 15258 12118 15260
rect 12142 15258 12198 15260
rect 11902 15206 11948 15258
rect 11948 15206 11958 15258
rect 11982 15206 12012 15258
rect 12012 15206 12024 15258
rect 12024 15206 12038 15258
rect 12062 15206 12076 15258
rect 12076 15206 12088 15258
rect 12088 15206 12118 15258
rect 12142 15206 12152 15258
rect 12152 15206 12198 15258
rect 11902 15204 11958 15206
rect 11982 15204 12038 15206
rect 12062 15204 12118 15206
rect 12142 15204 12198 15206
rect 11902 14170 11958 14172
rect 11982 14170 12038 14172
rect 12062 14170 12118 14172
rect 12142 14170 12198 14172
rect 11902 14118 11948 14170
rect 11948 14118 11958 14170
rect 11982 14118 12012 14170
rect 12012 14118 12024 14170
rect 12024 14118 12038 14170
rect 12062 14118 12076 14170
rect 12076 14118 12088 14170
rect 12088 14118 12118 14170
rect 12142 14118 12152 14170
rect 12152 14118 12198 14170
rect 11902 14116 11958 14118
rect 11982 14116 12038 14118
rect 12062 14116 12118 14118
rect 12142 14116 12198 14118
rect 11902 13082 11958 13084
rect 11982 13082 12038 13084
rect 12062 13082 12118 13084
rect 12142 13082 12198 13084
rect 11902 13030 11948 13082
rect 11948 13030 11958 13082
rect 11982 13030 12012 13082
rect 12012 13030 12024 13082
rect 12024 13030 12038 13082
rect 12062 13030 12076 13082
rect 12076 13030 12088 13082
rect 12088 13030 12118 13082
rect 12142 13030 12152 13082
rect 12152 13030 12198 13082
rect 11902 13028 11958 13030
rect 11982 13028 12038 13030
rect 12062 13028 12118 13030
rect 12142 13028 12198 13030
rect 6429 8186 6485 8188
rect 6509 8186 6565 8188
rect 6589 8186 6645 8188
rect 6669 8186 6725 8188
rect 6429 8134 6475 8186
rect 6475 8134 6485 8186
rect 6509 8134 6539 8186
rect 6539 8134 6551 8186
rect 6551 8134 6565 8186
rect 6589 8134 6603 8186
rect 6603 8134 6615 8186
rect 6615 8134 6645 8186
rect 6669 8134 6679 8186
rect 6679 8134 6725 8186
rect 6429 8132 6485 8134
rect 6509 8132 6565 8134
rect 6589 8132 6645 8134
rect 6669 8132 6725 8134
rect 6429 7098 6485 7100
rect 6509 7098 6565 7100
rect 6589 7098 6645 7100
rect 6669 7098 6725 7100
rect 6429 7046 6475 7098
rect 6475 7046 6485 7098
rect 6509 7046 6539 7098
rect 6539 7046 6551 7098
rect 6551 7046 6565 7098
rect 6589 7046 6603 7098
rect 6603 7046 6615 7098
rect 6615 7046 6645 7098
rect 6669 7046 6679 7098
rect 6679 7046 6725 7098
rect 6429 7044 6485 7046
rect 6509 7044 6565 7046
rect 6589 7044 6645 7046
rect 6669 7044 6725 7046
rect 6429 6010 6485 6012
rect 6509 6010 6565 6012
rect 6589 6010 6645 6012
rect 6669 6010 6725 6012
rect 6429 5958 6475 6010
rect 6475 5958 6485 6010
rect 6509 5958 6539 6010
rect 6539 5958 6551 6010
rect 6551 5958 6565 6010
rect 6589 5958 6603 6010
rect 6603 5958 6615 6010
rect 6615 5958 6645 6010
rect 6669 5958 6679 6010
rect 6679 5958 6725 6010
rect 6429 5956 6485 5958
rect 6509 5956 6565 5958
rect 6589 5956 6645 5958
rect 6669 5956 6725 5958
rect 11902 11994 11958 11996
rect 11982 11994 12038 11996
rect 12062 11994 12118 11996
rect 12142 11994 12198 11996
rect 11902 11942 11948 11994
rect 11948 11942 11958 11994
rect 11982 11942 12012 11994
rect 12012 11942 12024 11994
rect 12024 11942 12038 11994
rect 12062 11942 12076 11994
rect 12076 11942 12088 11994
rect 12088 11942 12118 11994
rect 12142 11942 12152 11994
rect 12152 11942 12198 11994
rect 11902 11940 11958 11942
rect 11982 11940 12038 11942
rect 12062 11940 12118 11942
rect 12142 11940 12198 11942
rect 11902 10906 11958 10908
rect 11982 10906 12038 10908
rect 12062 10906 12118 10908
rect 12142 10906 12198 10908
rect 11902 10854 11948 10906
rect 11948 10854 11958 10906
rect 11982 10854 12012 10906
rect 12012 10854 12024 10906
rect 12024 10854 12038 10906
rect 12062 10854 12076 10906
rect 12076 10854 12088 10906
rect 12088 10854 12118 10906
rect 12142 10854 12152 10906
rect 12152 10854 12198 10906
rect 11902 10852 11958 10854
rect 11982 10852 12038 10854
rect 12062 10852 12118 10854
rect 12142 10852 12198 10854
rect 11902 9818 11958 9820
rect 11982 9818 12038 9820
rect 12062 9818 12118 9820
rect 12142 9818 12198 9820
rect 11902 9766 11948 9818
rect 11948 9766 11958 9818
rect 11982 9766 12012 9818
rect 12012 9766 12024 9818
rect 12024 9766 12038 9818
rect 12062 9766 12076 9818
rect 12076 9766 12088 9818
rect 12088 9766 12118 9818
rect 12142 9766 12152 9818
rect 12152 9766 12198 9818
rect 11902 9764 11958 9766
rect 11982 9764 12038 9766
rect 12062 9764 12118 9766
rect 12142 9764 12198 9766
rect 6182 5208 6238 5264
rect 8390 5752 8446 5808
rect 6429 4922 6485 4924
rect 6509 4922 6565 4924
rect 6589 4922 6645 4924
rect 6669 4922 6725 4924
rect 6429 4870 6475 4922
rect 6475 4870 6485 4922
rect 6509 4870 6539 4922
rect 6539 4870 6551 4922
rect 6551 4870 6565 4922
rect 6589 4870 6603 4922
rect 6603 4870 6615 4922
rect 6615 4870 6645 4922
rect 6669 4870 6679 4922
rect 6679 4870 6725 4922
rect 6429 4868 6485 4870
rect 6509 4868 6565 4870
rect 6589 4868 6645 4870
rect 6669 4868 6725 4870
rect 6429 3834 6485 3836
rect 6509 3834 6565 3836
rect 6589 3834 6645 3836
rect 6669 3834 6725 3836
rect 6429 3782 6475 3834
rect 6475 3782 6485 3834
rect 6509 3782 6539 3834
rect 6539 3782 6551 3834
rect 6551 3782 6565 3834
rect 6589 3782 6603 3834
rect 6603 3782 6615 3834
rect 6615 3782 6645 3834
rect 6669 3782 6679 3834
rect 6679 3782 6725 3834
rect 6429 3780 6485 3782
rect 6509 3780 6565 3782
rect 6589 3780 6645 3782
rect 6669 3780 6725 3782
rect 938 3476 940 3496
rect 940 3476 992 3496
rect 992 3476 994 3496
rect 938 3440 994 3476
rect 938 1400 994 1456
rect 11902 8730 11958 8732
rect 11982 8730 12038 8732
rect 12062 8730 12118 8732
rect 12142 8730 12198 8732
rect 11902 8678 11948 8730
rect 11948 8678 11958 8730
rect 11982 8678 12012 8730
rect 12012 8678 12024 8730
rect 12024 8678 12038 8730
rect 12062 8678 12076 8730
rect 12076 8678 12088 8730
rect 12088 8678 12118 8730
rect 12142 8678 12152 8730
rect 12152 8678 12198 8730
rect 11902 8676 11958 8678
rect 11982 8676 12038 8678
rect 12062 8676 12118 8678
rect 12142 8676 12198 8678
rect 11902 7642 11958 7644
rect 11982 7642 12038 7644
rect 12062 7642 12118 7644
rect 12142 7642 12198 7644
rect 11902 7590 11948 7642
rect 11948 7590 11958 7642
rect 11982 7590 12012 7642
rect 12012 7590 12024 7642
rect 12024 7590 12038 7642
rect 12062 7590 12076 7642
rect 12076 7590 12088 7642
rect 12088 7590 12118 7642
rect 12142 7590 12152 7642
rect 12152 7590 12198 7642
rect 11902 7588 11958 7590
rect 11982 7588 12038 7590
rect 12062 7588 12118 7590
rect 12142 7588 12198 7590
rect 11902 6554 11958 6556
rect 11982 6554 12038 6556
rect 12062 6554 12118 6556
rect 12142 6554 12198 6556
rect 11902 6502 11948 6554
rect 11948 6502 11958 6554
rect 11982 6502 12012 6554
rect 12012 6502 12024 6554
rect 12024 6502 12038 6554
rect 12062 6502 12076 6554
rect 12076 6502 12088 6554
rect 12088 6502 12118 6554
rect 12142 6502 12152 6554
rect 12152 6502 12198 6554
rect 11902 6500 11958 6502
rect 11982 6500 12038 6502
rect 12062 6500 12118 6502
rect 12142 6500 12198 6502
rect 11902 5466 11958 5468
rect 11982 5466 12038 5468
rect 12062 5466 12118 5468
rect 12142 5466 12198 5468
rect 11902 5414 11948 5466
rect 11948 5414 11958 5466
rect 11982 5414 12012 5466
rect 12012 5414 12024 5466
rect 12024 5414 12038 5466
rect 12062 5414 12076 5466
rect 12076 5414 12088 5466
rect 12088 5414 12118 5466
rect 12142 5414 12152 5466
rect 12152 5414 12198 5466
rect 11902 5412 11958 5414
rect 11982 5412 12038 5414
rect 12062 5412 12118 5414
rect 12142 5412 12198 5414
rect 17376 16890 17432 16892
rect 17456 16890 17512 16892
rect 17536 16890 17592 16892
rect 17616 16890 17672 16892
rect 17376 16838 17422 16890
rect 17422 16838 17432 16890
rect 17456 16838 17486 16890
rect 17486 16838 17498 16890
rect 17498 16838 17512 16890
rect 17536 16838 17550 16890
rect 17550 16838 17562 16890
rect 17562 16838 17592 16890
rect 17616 16838 17626 16890
rect 17626 16838 17672 16890
rect 17376 16836 17432 16838
rect 17456 16836 17512 16838
rect 17536 16836 17592 16838
rect 17616 16836 17672 16838
rect 22849 17434 22905 17436
rect 22929 17434 22985 17436
rect 23009 17434 23065 17436
rect 23089 17434 23145 17436
rect 22849 17382 22895 17434
rect 22895 17382 22905 17434
rect 22929 17382 22959 17434
rect 22959 17382 22971 17434
rect 22971 17382 22985 17434
rect 23009 17382 23023 17434
rect 23023 17382 23035 17434
rect 23035 17382 23065 17434
rect 23089 17382 23099 17434
rect 23099 17382 23145 17434
rect 22849 17380 22905 17382
rect 22929 17380 22985 17382
rect 23009 17380 23065 17382
rect 23089 17380 23145 17382
rect 33796 17434 33852 17436
rect 33876 17434 33932 17436
rect 33956 17434 34012 17436
rect 34036 17434 34092 17436
rect 33796 17382 33842 17434
rect 33842 17382 33852 17434
rect 33876 17382 33906 17434
rect 33906 17382 33918 17434
rect 33918 17382 33932 17434
rect 33956 17382 33970 17434
rect 33970 17382 33982 17434
rect 33982 17382 34012 17434
rect 34036 17382 34046 17434
rect 34046 17382 34092 17434
rect 33796 17380 33852 17382
rect 33876 17380 33932 17382
rect 33956 17380 34012 17382
rect 34036 17380 34092 17382
rect 17376 15802 17432 15804
rect 17456 15802 17512 15804
rect 17536 15802 17592 15804
rect 17616 15802 17672 15804
rect 17376 15750 17422 15802
rect 17422 15750 17432 15802
rect 17456 15750 17486 15802
rect 17486 15750 17498 15802
rect 17498 15750 17512 15802
rect 17536 15750 17550 15802
rect 17550 15750 17562 15802
rect 17562 15750 17592 15802
rect 17616 15750 17626 15802
rect 17626 15750 17672 15802
rect 17376 15748 17432 15750
rect 17456 15748 17512 15750
rect 17536 15748 17592 15750
rect 17616 15748 17672 15750
rect 22849 16346 22905 16348
rect 22929 16346 22985 16348
rect 23009 16346 23065 16348
rect 23089 16346 23145 16348
rect 22849 16294 22895 16346
rect 22895 16294 22905 16346
rect 22929 16294 22959 16346
rect 22959 16294 22971 16346
rect 22971 16294 22985 16346
rect 23009 16294 23023 16346
rect 23023 16294 23035 16346
rect 23035 16294 23065 16346
rect 23089 16294 23099 16346
rect 23099 16294 23145 16346
rect 22849 16292 22905 16294
rect 22929 16292 22985 16294
rect 23009 16292 23065 16294
rect 23089 16292 23145 16294
rect 16578 13912 16634 13968
rect 13358 5480 13414 5536
rect 11902 4378 11958 4380
rect 11982 4378 12038 4380
rect 12062 4378 12118 4380
rect 12142 4378 12198 4380
rect 11902 4326 11948 4378
rect 11948 4326 11958 4378
rect 11982 4326 12012 4378
rect 12012 4326 12024 4378
rect 12024 4326 12038 4378
rect 12062 4326 12076 4378
rect 12076 4326 12088 4378
rect 12088 4326 12118 4378
rect 12142 4326 12152 4378
rect 12152 4326 12198 4378
rect 11902 4324 11958 4326
rect 11982 4324 12038 4326
rect 12062 4324 12118 4326
rect 12142 4324 12198 4326
rect 11902 3290 11958 3292
rect 11982 3290 12038 3292
rect 12062 3290 12118 3292
rect 12142 3290 12198 3292
rect 11902 3238 11948 3290
rect 11948 3238 11958 3290
rect 11982 3238 12012 3290
rect 12012 3238 12024 3290
rect 12024 3238 12038 3290
rect 12062 3238 12076 3290
rect 12076 3238 12088 3290
rect 12088 3238 12118 3290
rect 12142 3238 12152 3290
rect 12152 3238 12198 3290
rect 11902 3236 11958 3238
rect 11982 3236 12038 3238
rect 12062 3236 12118 3238
rect 12142 3236 12198 3238
rect 6429 2746 6485 2748
rect 6509 2746 6565 2748
rect 6589 2746 6645 2748
rect 6669 2746 6725 2748
rect 6429 2694 6475 2746
rect 6475 2694 6485 2746
rect 6509 2694 6539 2746
rect 6539 2694 6551 2746
rect 6551 2694 6565 2746
rect 6589 2694 6603 2746
rect 6603 2694 6615 2746
rect 6615 2694 6645 2746
rect 6669 2694 6679 2746
rect 6679 2694 6725 2746
rect 6429 2692 6485 2694
rect 6509 2692 6565 2694
rect 6589 2692 6645 2694
rect 6669 2692 6725 2694
rect 11902 2202 11958 2204
rect 11982 2202 12038 2204
rect 12062 2202 12118 2204
rect 12142 2202 12198 2204
rect 11902 2150 11948 2202
rect 11948 2150 11958 2202
rect 11982 2150 12012 2202
rect 12012 2150 12024 2202
rect 12024 2150 12038 2202
rect 12062 2150 12076 2202
rect 12076 2150 12088 2202
rect 12088 2150 12118 2202
rect 12142 2150 12152 2202
rect 12152 2150 12198 2202
rect 11902 2148 11958 2150
rect 11982 2148 12038 2150
rect 12062 2148 12118 2150
rect 12142 2148 12198 2150
rect 14462 5616 14518 5672
rect 17376 14714 17432 14716
rect 17456 14714 17512 14716
rect 17536 14714 17592 14716
rect 17616 14714 17672 14716
rect 17376 14662 17422 14714
rect 17422 14662 17432 14714
rect 17456 14662 17486 14714
rect 17486 14662 17498 14714
rect 17498 14662 17512 14714
rect 17536 14662 17550 14714
rect 17550 14662 17562 14714
rect 17562 14662 17592 14714
rect 17616 14662 17626 14714
rect 17626 14662 17672 14714
rect 17376 14660 17432 14662
rect 17456 14660 17512 14662
rect 17536 14660 17592 14662
rect 17616 14660 17672 14662
rect 22849 15258 22905 15260
rect 22929 15258 22985 15260
rect 23009 15258 23065 15260
rect 23089 15258 23145 15260
rect 22849 15206 22895 15258
rect 22895 15206 22905 15258
rect 22929 15206 22959 15258
rect 22959 15206 22971 15258
rect 22971 15206 22985 15258
rect 23009 15206 23023 15258
rect 23023 15206 23035 15258
rect 23035 15206 23065 15258
rect 23089 15206 23099 15258
rect 23099 15206 23145 15258
rect 22849 15204 22905 15206
rect 22929 15204 22985 15206
rect 23009 15204 23065 15206
rect 23089 15204 23145 15206
rect 17376 13626 17432 13628
rect 17456 13626 17512 13628
rect 17536 13626 17592 13628
rect 17616 13626 17672 13628
rect 17376 13574 17422 13626
rect 17422 13574 17432 13626
rect 17456 13574 17486 13626
rect 17486 13574 17498 13626
rect 17498 13574 17512 13626
rect 17536 13574 17550 13626
rect 17550 13574 17562 13626
rect 17562 13574 17592 13626
rect 17616 13574 17626 13626
rect 17626 13574 17672 13626
rect 17376 13572 17432 13574
rect 17456 13572 17512 13574
rect 17536 13572 17592 13574
rect 17616 13572 17672 13574
rect 17376 12538 17432 12540
rect 17456 12538 17512 12540
rect 17536 12538 17592 12540
rect 17616 12538 17672 12540
rect 17376 12486 17422 12538
rect 17422 12486 17432 12538
rect 17456 12486 17486 12538
rect 17486 12486 17498 12538
rect 17498 12486 17512 12538
rect 17536 12486 17550 12538
rect 17550 12486 17562 12538
rect 17562 12486 17592 12538
rect 17616 12486 17626 12538
rect 17626 12486 17672 12538
rect 17376 12484 17432 12486
rect 17456 12484 17512 12486
rect 17536 12484 17592 12486
rect 17616 12484 17672 12486
rect 17376 11450 17432 11452
rect 17456 11450 17512 11452
rect 17536 11450 17592 11452
rect 17616 11450 17672 11452
rect 17376 11398 17422 11450
rect 17422 11398 17432 11450
rect 17456 11398 17486 11450
rect 17486 11398 17498 11450
rect 17498 11398 17512 11450
rect 17536 11398 17550 11450
rect 17550 11398 17562 11450
rect 17562 11398 17592 11450
rect 17616 11398 17626 11450
rect 17626 11398 17672 11450
rect 17376 11396 17432 11398
rect 17456 11396 17512 11398
rect 17536 11396 17592 11398
rect 17616 11396 17672 11398
rect 17958 10512 18014 10568
rect 17376 10362 17432 10364
rect 17456 10362 17512 10364
rect 17536 10362 17592 10364
rect 17616 10362 17672 10364
rect 17376 10310 17422 10362
rect 17422 10310 17432 10362
rect 17456 10310 17486 10362
rect 17486 10310 17498 10362
rect 17498 10310 17512 10362
rect 17536 10310 17550 10362
rect 17550 10310 17562 10362
rect 17562 10310 17592 10362
rect 17616 10310 17626 10362
rect 17626 10310 17672 10362
rect 17376 10308 17432 10310
rect 17456 10308 17512 10310
rect 17536 10308 17592 10310
rect 17616 10308 17672 10310
rect 17376 9274 17432 9276
rect 17456 9274 17512 9276
rect 17536 9274 17592 9276
rect 17616 9274 17672 9276
rect 17376 9222 17422 9274
rect 17422 9222 17432 9274
rect 17456 9222 17486 9274
rect 17486 9222 17498 9274
rect 17498 9222 17512 9274
rect 17536 9222 17550 9274
rect 17550 9222 17562 9274
rect 17562 9222 17592 9274
rect 17616 9222 17626 9274
rect 17626 9222 17672 9274
rect 17376 9220 17432 9222
rect 17456 9220 17512 9222
rect 17536 9220 17592 9222
rect 17616 9220 17672 9222
rect 17376 8186 17432 8188
rect 17456 8186 17512 8188
rect 17536 8186 17592 8188
rect 17616 8186 17672 8188
rect 17376 8134 17422 8186
rect 17422 8134 17432 8186
rect 17456 8134 17486 8186
rect 17486 8134 17498 8186
rect 17498 8134 17512 8186
rect 17536 8134 17550 8186
rect 17550 8134 17562 8186
rect 17562 8134 17592 8186
rect 17616 8134 17626 8186
rect 17626 8134 17672 8186
rect 17376 8132 17432 8134
rect 17456 8132 17512 8134
rect 17536 8132 17592 8134
rect 17616 8132 17672 8134
rect 19706 10004 19708 10024
rect 19708 10004 19760 10024
rect 19760 10004 19762 10024
rect 19706 9968 19762 10004
rect 22006 9716 22062 9752
rect 22006 9696 22008 9716
rect 22008 9696 22060 9716
rect 22060 9696 22062 9716
rect 17376 7098 17432 7100
rect 17456 7098 17512 7100
rect 17536 7098 17592 7100
rect 17616 7098 17672 7100
rect 17376 7046 17422 7098
rect 17422 7046 17432 7098
rect 17456 7046 17486 7098
rect 17486 7046 17498 7098
rect 17498 7046 17512 7098
rect 17536 7046 17550 7098
rect 17550 7046 17562 7098
rect 17562 7046 17592 7098
rect 17616 7046 17626 7098
rect 17626 7046 17672 7098
rect 17376 7044 17432 7046
rect 17456 7044 17512 7046
rect 17536 7044 17592 7046
rect 17616 7044 17672 7046
rect 17376 6010 17432 6012
rect 17456 6010 17512 6012
rect 17536 6010 17592 6012
rect 17616 6010 17672 6012
rect 17376 5958 17422 6010
rect 17422 5958 17432 6010
rect 17456 5958 17486 6010
rect 17486 5958 17498 6010
rect 17498 5958 17512 6010
rect 17536 5958 17550 6010
rect 17550 5958 17562 6010
rect 17562 5958 17592 6010
rect 17616 5958 17626 6010
rect 17626 5958 17672 6010
rect 17376 5956 17432 5958
rect 17456 5956 17512 5958
rect 17536 5956 17592 5958
rect 17616 5956 17672 5958
rect 15842 5108 15844 5128
rect 15844 5108 15896 5128
rect 15896 5108 15898 5128
rect 15842 5072 15898 5108
rect 17376 4922 17432 4924
rect 17456 4922 17512 4924
rect 17536 4922 17592 4924
rect 17616 4922 17672 4924
rect 17376 4870 17422 4922
rect 17422 4870 17432 4922
rect 17456 4870 17486 4922
rect 17486 4870 17498 4922
rect 17498 4870 17512 4922
rect 17536 4870 17550 4922
rect 17550 4870 17562 4922
rect 17562 4870 17592 4922
rect 17616 4870 17626 4922
rect 17626 4870 17672 4922
rect 17376 4868 17432 4870
rect 17456 4868 17512 4870
rect 17536 4868 17592 4870
rect 17616 4868 17672 4870
rect 17376 3834 17432 3836
rect 17456 3834 17512 3836
rect 17536 3834 17592 3836
rect 17616 3834 17672 3836
rect 17376 3782 17422 3834
rect 17422 3782 17432 3834
rect 17456 3782 17486 3834
rect 17486 3782 17498 3834
rect 17498 3782 17512 3834
rect 17536 3782 17550 3834
rect 17550 3782 17562 3834
rect 17562 3782 17592 3834
rect 17616 3782 17626 3834
rect 17626 3782 17672 3834
rect 17376 3780 17432 3782
rect 17456 3780 17512 3782
rect 17536 3780 17592 3782
rect 17616 3780 17672 3782
rect 17376 2746 17432 2748
rect 17456 2746 17512 2748
rect 17536 2746 17592 2748
rect 17616 2746 17672 2748
rect 17376 2694 17422 2746
rect 17422 2694 17432 2746
rect 17456 2694 17486 2746
rect 17486 2694 17498 2746
rect 17498 2694 17512 2746
rect 17536 2694 17550 2746
rect 17550 2694 17562 2746
rect 17562 2694 17592 2746
rect 17616 2694 17626 2746
rect 17626 2694 17672 2746
rect 17376 2692 17432 2694
rect 17456 2692 17512 2694
rect 17536 2692 17592 2694
rect 17616 2692 17672 2694
rect 28323 16890 28379 16892
rect 28403 16890 28459 16892
rect 28483 16890 28539 16892
rect 28563 16890 28619 16892
rect 28323 16838 28369 16890
rect 28369 16838 28379 16890
rect 28403 16838 28433 16890
rect 28433 16838 28445 16890
rect 28445 16838 28459 16890
rect 28483 16838 28497 16890
rect 28497 16838 28509 16890
rect 28509 16838 28539 16890
rect 28563 16838 28573 16890
rect 28573 16838 28619 16890
rect 28323 16836 28379 16838
rect 28403 16836 28459 16838
rect 28483 16836 28539 16838
rect 28563 16836 28619 16838
rect 28323 15802 28379 15804
rect 28403 15802 28459 15804
rect 28483 15802 28539 15804
rect 28563 15802 28619 15804
rect 28323 15750 28369 15802
rect 28369 15750 28379 15802
rect 28403 15750 28433 15802
rect 28433 15750 28445 15802
rect 28445 15750 28459 15802
rect 28483 15750 28497 15802
rect 28497 15750 28509 15802
rect 28509 15750 28539 15802
rect 28563 15750 28573 15802
rect 28573 15750 28619 15802
rect 28323 15748 28379 15750
rect 28403 15748 28459 15750
rect 28483 15748 28539 15750
rect 28563 15748 28619 15750
rect 23662 14340 23718 14376
rect 23662 14320 23664 14340
rect 23664 14320 23716 14340
rect 23716 14320 23718 14340
rect 22849 14170 22905 14172
rect 22929 14170 22985 14172
rect 23009 14170 23065 14172
rect 23089 14170 23145 14172
rect 22849 14118 22895 14170
rect 22895 14118 22905 14170
rect 22929 14118 22959 14170
rect 22959 14118 22971 14170
rect 22971 14118 22985 14170
rect 23009 14118 23023 14170
rect 23023 14118 23035 14170
rect 23035 14118 23065 14170
rect 23089 14118 23099 14170
rect 23099 14118 23145 14170
rect 22849 14116 22905 14118
rect 22929 14116 22985 14118
rect 23009 14116 23065 14118
rect 23089 14116 23145 14118
rect 22282 9696 22338 9752
rect 18510 5480 18566 5536
rect 17958 5108 17960 5128
rect 17960 5108 18012 5128
rect 18012 5108 18014 5128
rect 17958 5072 18014 5108
rect 22849 13082 22905 13084
rect 22929 13082 22985 13084
rect 23009 13082 23065 13084
rect 23089 13082 23145 13084
rect 22849 13030 22895 13082
rect 22895 13030 22905 13082
rect 22929 13030 22959 13082
rect 22959 13030 22971 13082
rect 22971 13030 22985 13082
rect 23009 13030 23023 13082
rect 23023 13030 23035 13082
rect 23035 13030 23065 13082
rect 23089 13030 23099 13082
rect 23099 13030 23145 13082
rect 22849 13028 22905 13030
rect 22929 13028 22985 13030
rect 23009 13028 23065 13030
rect 23089 13028 23145 13030
rect 22849 11994 22905 11996
rect 22929 11994 22985 11996
rect 23009 11994 23065 11996
rect 23089 11994 23145 11996
rect 22849 11942 22895 11994
rect 22895 11942 22905 11994
rect 22929 11942 22959 11994
rect 22959 11942 22971 11994
rect 22971 11942 22985 11994
rect 23009 11942 23023 11994
rect 23023 11942 23035 11994
rect 23035 11942 23065 11994
rect 23089 11942 23099 11994
rect 23099 11942 23145 11994
rect 22849 11940 22905 11942
rect 22929 11940 22985 11942
rect 23009 11940 23065 11942
rect 23089 11940 23145 11942
rect 22849 10906 22905 10908
rect 22929 10906 22985 10908
rect 23009 10906 23065 10908
rect 23089 10906 23145 10908
rect 22849 10854 22895 10906
rect 22895 10854 22905 10906
rect 22929 10854 22959 10906
rect 22959 10854 22971 10906
rect 22971 10854 22985 10906
rect 23009 10854 23023 10906
rect 23023 10854 23035 10906
rect 23035 10854 23065 10906
rect 23089 10854 23099 10906
rect 23099 10854 23145 10906
rect 22849 10852 22905 10854
rect 22929 10852 22985 10854
rect 23009 10852 23065 10854
rect 23089 10852 23145 10854
rect 23662 10512 23718 10568
rect 22849 9818 22905 9820
rect 22929 9818 22985 9820
rect 23009 9818 23065 9820
rect 23089 9818 23145 9820
rect 22849 9766 22895 9818
rect 22895 9766 22905 9818
rect 22929 9766 22959 9818
rect 22959 9766 22971 9818
rect 22971 9766 22985 9818
rect 23009 9766 23023 9818
rect 23023 9766 23035 9818
rect 23035 9766 23065 9818
rect 23089 9766 23099 9818
rect 23099 9766 23145 9818
rect 22849 9764 22905 9766
rect 22929 9764 22985 9766
rect 23009 9764 23065 9766
rect 23089 9764 23145 9766
rect 22849 8730 22905 8732
rect 22929 8730 22985 8732
rect 23009 8730 23065 8732
rect 23089 8730 23145 8732
rect 22849 8678 22895 8730
rect 22895 8678 22905 8730
rect 22929 8678 22959 8730
rect 22959 8678 22971 8730
rect 22971 8678 22985 8730
rect 23009 8678 23023 8730
rect 23023 8678 23035 8730
rect 23035 8678 23065 8730
rect 23089 8678 23099 8730
rect 23099 8678 23145 8730
rect 22849 8676 22905 8678
rect 22929 8676 22985 8678
rect 23009 8676 23065 8678
rect 23089 8676 23145 8678
rect 22849 7642 22905 7644
rect 22929 7642 22985 7644
rect 23009 7642 23065 7644
rect 23089 7642 23145 7644
rect 22849 7590 22895 7642
rect 22895 7590 22905 7642
rect 22929 7590 22959 7642
rect 22959 7590 22971 7642
rect 22971 7590 22985 7642
rect 23009 7590 23023 7642
rect 23023 7590 23035 7642
rect 23035 7590 23065 7642
rect 23089 7590 23099 7642
rect 23099 7590 23145 7642
rect 22849 7588 22905 7590
rect 22929 7588 22985 7590
rect 23009 7588 23065 7590
rect 23089 7588 23145 7590
rect 22849 6554 22905 6556
rect 22929 6554 22985 6556
rect 23009 6554 23065 6556
rect 23089 6554 23145 6556
rect 22849 6502 22895 6554
rect 22895 6502 22905 6554
rect 22929 6502 22959 6554
rect 22959 6502 22971 6554
rect 22971 6502 22985 6554
rect 23009 6502 23023 6554
rect 23023 6502 23035 6554
rect 23035 6502 23065 6554
rect 23089 6502 23099 6554
rect 23099 6502 23145 6554
rect 22849 6500 22905 6502
rect 22929 6500 22985 6502
rect 23009 6500 23065 6502
rect 23089 6500 23145 6502
rect 22849 5466 22905 5468
rect 22929 5466 22985 5468
rect 23009 5466 23065 5468
rect 23089 5466 23145 5468
rect 22849 5414 22895 5466
rect 22895 5414 22905 5466
rect 22929 5414 22959 5466
rect 22959 5414 22971 5466
rect 22971 5414 22985 5466
rect 23009 5414 23023 5466
rect 23023 5414 23035 5466
rect 23035 5414 23065 5466
rect 23089 5414 23099 5466
rect 23099 5414 23145 5466
rect 22849 5412 22905 5414
rect 22929 5412 22985 5414
rect 23009 5412 23065 5414
rect 23089 5412 23145 5414
rect 22849 4378 22905 4380
rect 22929 4378 22985 4380
rect 23009 4378 23065 4380
rect 23089 4378 23145 4380
rect 22849 4326 22895 4378
rect 22895 4326 22905 4378
rect 22929 4326 22959 4378
rect 22959 4326 22971 4378
rect 22971 4326 22985 4378
rect 23009 4326 23023 4378
rect 23023 4326 23035 4378
rect 23035 4326 23065 4378
rect 23089 4326 23099 4378
rect 23099 4326 23145 4378
rect 22849 4324 22905 4326
rect 22929 4324 22985 4326
rect 23009 4324 23065 4326
rect 23089 4324 23145 4326
rect 23846 9596 23848 9616
rect 23848 9596 23900 9616
rect 23900 9596 23902 9616
rect 23846 9560 23902 9596
rect 24766 9968 24822 10024
rect 23938 5752 23994 5808
rect 25870 5652 25872 5672
rect 25872 5652 25924 5672
rect 25924 5652 25926 5672
rect 25870 5616 25926 5652
rect 28323 14714 28379 14716
rect 28403 14714 28459 14716
rect 28483 14714 28539 14716
rect 28563 14714 28619 14716
rect 28323 14662 28369 14714
rect 28369 14662 28379 14714
rect 28403 14662 28433 14714
rect 28433 14662 28445 14714
rect 28445 14662 28459 14714
rect 28483 14662 28497 14714
rect 28497 14662 28509 14714
rect 28509 14662 28539 14714
rect 28563 14662 28573 14714
rect 28573 14662 28619 14714
rect 28323 14660 28379 14662
rect 28403 14660 28459 14662
rect 28483 14660 28539 14662
rect 28563 14660 28619 14662
rect 28323 13626 28379 13628
rect 28403 13626 28459 13628
rect 28483 13626 28539 13628
rect 28563 13626 28619 13628
rect 28323 13574 28369 13626
rect 28369 13574 28379 13626
rect 28403 13574 28433 13626
rect 28433 13574 28445 13626
rect 28445 13574 28459 13626
rect 28483 13574 28497 13626
rect 28497 13574 28509 13626
rect 28509 13574 28539 13626
rect 28563 13574 28573 13626
rect 28573 13574 28619 13626
rect 28323 13572 28379 13574
rect 28403 13572 28459 13574
rect 28483 13572 28539 13574
rect 28563 13572 28619 13574
rect 28323 12538 28379 12540
rect 28403 12538 28459 12540
rect 28483 12538 28539 12540
rect 28563 12538 28619 12540
rect 28323 12486 28369 12538
rect 28369 12486 28379 12538
rect 28403 12486 28433 12538
rect 28433 12486 28445 12538
rect 28445 12486 28459 12538
rect 28483 12486 28497 12538
rect 28497 12486 28509 12538
rect 28509 12486 28539 12538
rect 28563 12486 28573 12538
rect 28573 12486 28619 12538
rect 28323 12484 28379 12486
rect 28403 12484 28459 12486
rect 28483 12484 28539 12486
rect 28563 12484 28619 12486
rect 28323 11450 28379 11452
rect 28403 11450 28459 11452
rect 28483 11450 28539 11452
rect 28563 11450 28619 11452
rect 28323 11398 28369 11450
rect 28369 11398 28379 11450
rect 28403 11398 28433 11450
rect 28433 11398 28445 11450
rect 28445 11398 28459 11450
rect 28483 11398 28497 11450
rect 28497 11398 28509 11450
rect 28509 11398 28539 11450
rect 28563 11398 28573 11450
rect 28573 11398 28619 11450
rect 28323 11396 28379 11398
rect 28403 11396 28459 11398
rect 28483 11396 28539 11398
rect 28563 11396 28619 11398
rect 27894 11056 27950 11112
rect 28078 10648 28134 10704
rect 27894 9560 27950 9616
rect 29090 10648 29146 10704
rect 28323 10362 28379 10364
rect 28403 10362 28459 10364
rect 28483 10362 28539 10364
rect 28563 10362 28619 10364
rect 28323 10310 28369 10362
rect 28369 10310 28379 10362
rect 28403 10310 28433 10362
rect 28433 10310 28445 10362
rect 28445 10310 28459 10362
rect 28483 10310 28497 10362
rect 28497 10310 28509 10362
rect 28509 10310 28539 10362
rect 28563 10310 28573 10362
rect 28573 10310 28619 10362
rect 28323 10308 28379 10310
rect 28403 10308 28459 10310
rect 28483 10308 28539 10310
rect 28563 10308 28619 10310
rect 28323 9274 28379 9276
rect 28403 9274 28459 9276
rect 28483 9274 28539 9276
rect 28563 9274 28619 9276
rect 28323 9222 28369 9274
rect 28369 9222 28379 9274
rect 28403 9222 28433 9274
rect 28433 9222 28445 9274
rect 28445 9222 28459 9274
rect 28483 9222 28497 9274
rect 28497 9222 28509 9274
rect 28509 9222 28539 9274
rect 28563 9222 28573 9274
rect 28573 9222 28619 9274
rect 28323 9220 28379 9222
rect 28403 9220 28459 9222
rect 28483 9220 28539 9222
rect 28563 9220 28619 9222
rect 31022 12144 31078 12200
rect 33796 16346 33852 16348
rect 33876 16346 33932 16348
rect 33956 16346 34012 16348
rect 34036 16346 34092 16348
rect 33796 16294 33842 16346
rect 33842 16294 33852 16346
rect 33876 16294 33906 16346
rect 33906 16294 33918 16346
rect 33918 16294 33932 16346
rect 33956 16294 33970 16346
rect 33970 16294 33982 16346
rect 33982 16294 34012 16346
rect 34036 16294 34046 16346
rect 34046 16294 34092 16346
rect 33796 16292 33852 16294
rect 33876 16292 33932 16294
rect 33956 16292 34012 16294
rect 34036 16292 34092 16294
rect 33796 15258 33852 15260
rect 33876 15258 33932 15260
rect 33956 15258 34012 15260
rect 34036 15258 34092 15260
rect 33796 15206 33842 15258
rect 33842 15206 33852 15258
rect 33876 15206 33906 15258
rect 33906 15206 33918 15258
rect 33918 15206 33932 15258
rect 33956 15206 33970 15258
rect 33970 15206 33982 15258
rect 33982 15206 34012 15258
rect 34036 15206 34046 15258
rect 34046 15206 34092 15258
rect 33796 15204 33852 15206
rect 33876 15204 33932 15206
rect 33956 15204 34012 15206
rect 34036 15204 34092 15206
rect 33796 14170 33852 14172
rect 33876 14170 33932 14172
rect 33956 14170 34012 14172
rect 34036 14170 34092 14172
rect 33796 14118 33842 14170
rect 33842 14118 33852 14170
rect 33876 14118 33906 14170
rect 33906 14118 33918 14170
rect 33918 14118 33932 14170
rect 33956 14118 33970 14170
rect 33970 14118 33982 14170
rect 33982 14118 34012 14170
rect 34036 14118 34046 14170
rect 34046 14118 34092 14170
rect 33796 14116 33852 14118
rect 33876 14116 33932 14118
rect 33956 14116 34012 14118
rect 34036 14116 34092 14118
rect 30102 8900 30158 8936
rect 30102 8880 30104 8900
rect 30104 8880 30156 8900
rect 30156 8880 30158 8900
rect 28323 8186 28379 8188
rect 28403 8186 28459 8188
rect 28483 8186 28539 8188
rect 28563 8186 28619 8188
rect 28323 8134 28369 8186
rect 28369 8134 28379 8186
rect 28403 8134 28433 8186
rect 28433 8134 28445 8186
rect 28445 8134 28459 8186
rect 28483 8134 28497 8186
rect 28497 8134 28509 8186
rect 28509 8134 28539 8186
rect 28563 8134 28573 8186
rect 28573 8134 28619 8186
rect 28323 8132 28379 8134
rect 28403 8132 28459 8134
rect 28483 8132 28539 8134
rect 28563 8132 28619 8134
rect 28323 7098 28379 7100
rect 28403 7098 28459 7100
rect 28483 7098 28539 7100
rect 28563 7098 28619 7100
rect 28323 7046 28369 7098
rect 28369 7046 28379 7098
rect 28403 7046 28433 7098
rect 28433 7046 28445 7098
rect 28445 7046 28459 7098
rect 28483 7046 28497 7098
rect 28497 7046 28509 7098
rect 28509 7046 28539 7098
rect 28563 7046 28573 7098
rect 28573 7046 28619 7098
rect 28323 7044 28379 7046
rect 28403 7044 28459 7046
rect 28483 7044 28539 7046
rect 28563 7044 28619 7046
rect 27526 6160 27582 6216
rect 28323 6010 28379 6012
rect 28403 6010 28459 6012
rect 28483 6010 28539 6012
rect 28563 6010 28619 6012
rect 28323 5958 28369 6010
rect 28369 5958 28379 6010
rect 28403 5958 28433 6010
rect 28433 5958 28445 6010
rect 28445 5958 28459 6010
rect 28483 5958 28497 6010
rect 28497 5958 28509 6010
rect 28509 5958 28539 6010
rect 28563 5958 28573 6010
rect 28573 5958 28619 6010
rect 28323 5956 28379 5958
rect 28403 5956 28459 5958
rect 28483 5956 28539 5958
rect 28563 5956 28619 5958
rect 27526 5752 27582 5808
rect 22849 3290 22905 3292
rect 22929 3290 22985 3292
rect 23009 3290 23065 3292
rect 23089 3290 23145 3292
rect 22849 3238 22895 3290
rect 22895 3238 22905 3290
rect 22929 3238 22959 3290
rect 22959 3238 22971 3290
rect 22971 3238 22985 3290
rect 23009 3238 23023 3290
rect 23023 3238 23035 3290
rect 23035 3238 23065 3290
rect 23089 3238 23099 3290
rect 23099 3238 23145 3290
rect 22849 3236 22905 3238
rect 22929 3236 22985 3238
rect 23009 3236 23065 3238
rect 23089 3236 23145 3238
rect 28323 4922 28379 4924
rect 28403 4922 28459 4924
rect 28483 4922 28539 4924
rect 28563 4922 28619 4924
rect 28323 4870 28369 4922
rect 28369 4870 28379 4922
rect 28403 4870 28433 4922
rect 28433 4870 28445 4922
rect 28445 4870 28459 4922
rect 28483 4870 28497 4922
rect 28497 4870 28509 4922
rect 28509 4870 28539 4922
rect 28563 4870 28573 4922
rect 28573 4870 28619 4922
rect 28323 4868 28379 4870
rect 28403 4868 28459 4870
rect 28483 4868 28539 4870
rect 28563 4868 28619 4870
rect 28323 3834 28379 3836
rect 28403 3834 28459 3836
rect 28483 3834 28539 3836
rect 28563 3834 28619 3836
rect 28323 3782 28369 3834
rect 28369 3782 28379 3834
rect 28403 3782 28433 3834
rect 28433 3782 28445 3834
rect 28445 3782 28459 3834
rect 28483 3782 28497 3834
rect 28497 3782 28509 3834
rect 28509 3782 28539 3834
rect 28563 3782 28573 3834
rect 28573 3782 28619 3834
rect 28323 3780 28379 3782
rect 28403 3780 28459 3782
rect 28483 3780 28539 3782
rect 28563 3780 28619 3782
rect 28323 2746 28379 2748
rect 28403 2746 28459 2748
rect 28483 2746 28539 2748
rect 28563 2746 28619 2748
rect 28323 2694 28369 2746
rect 28369 2694 28379 2746
rect 28403 2694 28433 2746
rect 28433 2694 28445 2746
rect 28445 2694 28459 2746
rect 28483 2694 28497 2746
rect 28497 2694 28509 2746
rect 28509 2694 28539 2746
rect 28563 2694 28573 2746
rect 28573 2694 28619 2746
rect 28323 2692 28379 2694
rect 28403 2692 28459 2694
rect 28483 2692 28539 2694
rect 28563 2692 28619 2694
rect 22849 2202 22905 2204
rect 22929 2202 22985 2204
rect 23009 2202 23065 2204
rect 23089 2202 23145 2204
rect 22849 2150 22895 2202
rect 22895 2150 22905 2202
rect 22929 2150 22959 2202
rect 22959 2150 22971 2202
rect 22971 2150 22985 2202
rect 23009 2150 23023 2202
rect 23023 2150 23035 2202
rect 23035 2150 23065 2202
rect 23089 2150 23099 2202
rect 23099 2150 23145 2202
rect 22849 2148 22905 2150
rect 22929 2148 22985 2150
rect 23009 2148 23065 2150
rect 23089 2148 23145 2150
rect 33796 13082 33852 13084
rect 33876 13082 33932 13084
rect 33956 13082 34012 13084
rect 34036 13082 34092 13084
rect 33796 13030 33842 13082
rect 33842 13030 33852 13082
rect 33876 13030 33906 13082
rect 33906 13030 33918 13082
rect 33918 13030 33932 13082
rect 33956 13030 33970 13082
rect 33970 13030 33982 13082
rect 33982 13030 34012 13082
rect 34036 13030 34046 13082
rect 34046 13030 34092 13082
rect 33796 13028 33852 13030
rect 33876 13028 33932 13030
rect 33956 13028 34012 13030
rect 34036 13028 34092 13030
rect 33796 11994 33852 11996
rect 33876 11994 33932 11996
rect 33956 11994 34012 11996
rect 34036 11994 34092 11996
rect 33796 11942 33842 11994
rect 33842 11942 33852 11994
rect 33876 11942 33906 11994
rect 33906 11942 33918 11994
rect 33918 11942 33932 11994
rect 33956 11942 33970 11994
rect 33970 11942 33982 11994
rect 33982 11942 34012 11994
rect 34036 11942 34046 11994
rect 34046 11942 34092 11994
rect 33796 11940 33852 11942
rect 33876 11940 33932 11942
rect 33956 11940 34012 11942
rect 34036 11940 34092 11942
rect 33796 10906 33852 10908
rect 33876 10906 33932 10908
rect 33956 10906 34012 10908
rect 34036 10906 34092 10908
rect 33796 10854 33842 10906
rect 33842 10854 33852 10906
rect 33876 10854 33906 10906
rect 33906 10854 33918 10906
rect 33918 10854 33932 10906
rect 33956 10854 33970 10906
rect 33970 10854 33982 10906
rect 33982 10854 34012 10906
rect 34036 10854 34046 10906
rect 34046 10854 34092 10906
rect 33796 10852 33852 10854
rect 33876 10852 33932 10854
rect 33956 10852 34012 10854
rect 34036 10852 34092 10854
rect 35070 11092 35072 11112
rect 35072 11092 35124 11112
rect 35124 11092 35126 11112
rect 35070 11056 35126 11092
rect 33796 9818 33852 9820
rect 33876 9818 33932 9820
rect 33956 9818 34012 9820
rect 34036 9818 34092 9820
rect 33796 9766 33842 9818
rect 33842 9766 33852 9818
rect 33876 9766 33906 9818
rect 33906 9766 33918 9818
rect 33918 9766 33932 9818
rect 33956 9766 33970 9818
rect 33970 9766 33982 9818
rect 33982 9766 34012 9818
rect 34036 9766 34046 9818
rect 34046 9766 34092 9818
rect 33796 9764 33852 9766
rect 33876 9764 33932 9766
rect 33956 9764 34012 9766
rect 34036 9764 34092 9766
rect 32862 9424 32918 9480
rect 32494 8880 32550 8936
rect 33796 8730 33852 8732
rect 33876 8730 33932 8732
rect 33956 8730 34012 8732
rect 34036 8730 34092 8732
rect 33796 8678 33842 8730
rect 33842 8678 33852 8730
rect 33876 8678 33906 8730
rect 33906 8678 33918 8730
rect 33918 8678 33932 8730
rect 33956 8678 33970 8730
rect 33970 8678 33982 8730
rect 33982 8678 34012 8730
rect 34036 8678 34046 8730
rect 34046 8678 34092 8730
rect 33796 8676 33852 8678
rect 33876 8676 33932 8678
rect 33956 8676 34012 8678
rect 34036 8676 34092 8678
rect 33414 8336 33470 8392
rect 34518 8472 34574 8528
rect 32954 7928 33010 7984
rect 33796 7642 33852 7644
rect 33876 7642 33932 7644
rect 33956 7642 34012 7644
rect 34036 7642 34092 7644
rect 33796 7590 33842 7642
rect 33842 7590 33852 7642
rect 33876 7590 33906 7642
rect 33906 7590 33918 7642
rect 33918 7590 33932 7642
rect 33956 7590 33970 7642
rect 33970 7590 33982 7642
rect 33982 7590 34012 7642
rect 34036 7590 34046 7642
rect 34046 7590 34092 7642
rect 33796 7588 33852 7590
rect 33876 7588 33932 7590
rect 33956 7588 34012 7590
rect 34036 7588 34092 7590
rect 33796 6554 33852 6556
rect 33876 6554 33932 6556
rect 33956 6554 34012 6556
rect 34036 6554 34092 6556
rect 33796 6502 33842 6554
rect 33842 6502 33852 6554
rect 33876 6502 33906 6554
rect 33906 6502 33918 6554
rect 33918 6502 33932 6554
rect 33956 6502 33970 6554
rect 33970 6502 33982 6554
rect 33982 6502 34012 6554
rect 34036 6502 34046 6554
rect 34046 6502 34092 6554
rect 33796 6500 33852 6502
rect 33876 6500 33932 6502
rect 33956 6500 34012 6502
rect 34036 6500 34092 6502
rect 34426 6840 34482 6896
rect 34518 6024 34574 6080
rect 39270 16890 39326 16892
rect 39350 16890 39406 16892
rect 39430 16890 39486 16892
rect 39510 16890 39566 16892
rect 39270 16838 39316 16890
rect 39316 16838 39326 16890
rect 39350 16838 39380 16890
rect 39380 16838 39392 16890
rect 39392 16838 39406 16890
rect 39430 16838 39444 16890
rect 39444 16838 39456 16890
rect 39456 16838 39486 16890
rect 39510 16838 39520 16890
rect 39520 16838 39566 16890
rect 39270 16836 39326 16838
rect 39350 16836 39406 16838
rect 39430 16836 39486 16838
rect 39510 16836 39566 16838
rect 45006 19080 45062 19136
rect 45006 17720 45062 17776
rect 39270 15802 39326 15804
rect 39350 15802 39406 15804
rect 39430 15802 39486 15804
rect 39510 15802 39566 15804
rect 39270 15750 39316 15802
rect 39316 15750 39326 15802
rect 39350 15750 39380 15802
rect 39380 15750 39392 15802
rect 39392 15750 39406 15802
rect 39430 15750 39444 15802
rect 39444 15750 39456 15802
rect 39456 15750 39486 15802
rect 39510 15750 39520 15802
rect 39520 15750 39566 15802
rect 39270 15748 39326 15750
rect 39350 15748 39406 15750
rect 39430 15748 39486 15750
rect 39510 15748 39566 15750
rect 38842 14320 38898 14376
rect 39270 14714 39326 14716
rect 39350 14714 39406 14716
rect 39430 14714 39486 14716
rect 39510 14714 39566 14716
rect 39270 14662 39316 14714
rect 39316 14662 39326 14714
rect 39350 14662 39380 14714
rect 39380 14662 39392 14714
rect 39392 14662 39406 14714
rect 39430 14662 39444 14714
rect 39444 14662 39456 14714
rect 39456 14662 39486 14714
rect 39510 14662 39520 14714
rect 39520 14662 39566 14714
rect 39270 14660 39326 14662
rect 39350 14660 39406 14662
rect 39430 14660 39486 14662
rect 39510 14660 39566 14662
rect 39270 13626 39326 13628
rect 39350 13626 39406 13628
rect 39430 13626 39486 13628
rect 39510 13626 39566 13628
rect 39270 13574 39316 13626
rect 39316 13574 39326 13626
rect 39350 13574 39380 13626
rect 39380 13574 39392 13626
rect 39392 13574 39406 13626
rect 39430 13574 39444 13626
rect 39444 13574 39456 13626
rect 39456 13574 39486 13626
rect 39510 13574 39520 13626
rect 39520 13574 39566 13626
rect 39270 13572 39326 13574
rect 39350 13572 39406 13574
rect 39430 13572 39486 13574
rect 39510 13572 39566 13574
rect 39270 12538 39326 12540
rect 39350 12538 39406 12540
rect 39430 12538 39486 12540
rect 39510 12538 39566 12540
rect 39270 12486 39316 12538
rect 39316 12486 39326 12538
rect 39350 12486 39380 12538
rect 39380 12486 39392 12538
rect 39392 12486 39406 12538
rect 39430 12486 39444 12538
rect 39444 12486 39456 12538
rect 39456 12486 39486 12538
rect 39510 12486 39520 12538
rect 39520 12486 39566 12538
rect 39270 12484 39326 12486
rect 39350 12484 39406 12486
rect 39430 12484 39486 12486
rect 39510 12484 39566 12486
rect 39270 11450 39326 11452
rect 39350 11450 39406 11452
rect 39430 11450 39486 11452
rect 39510 11450 39566 11452
rect 39270 11398 39316 11450
rect 39316 11398 39326 11450
rect 39350 11398 39380 11450
rect 39380 11398 39392 11450
rect 39392 11398 39406 11450
rect 39430 11398 39444 11450
rect 39444 11398 39456 11450
rect 39456 11398 39486 11450
rect 39510 11398 39520 11450
rect 39520 11398 39566 11450
rect 39270 11396 39326 11398
rect 39350 11396 39406 11398
rect 39430 11396 39486 11398
rect 39510 11396 39566 11398
rect 36082 7928 36138 7984
rect 34886 5636 34942 5672
rect 34886 5616 34888 5636
rect 34888 5616 34940 5636
rect 34940 5616 34942 5636
rect 33796 5466 33852 5468
rect 33876 5466 33932 5468
rect 33956 5466 34012 5468
rect 34036 5466 34092 5468
rect 33796 5414 33842 5466
rect 33842 5414 33852 5466
rect 33876 5414 33906 5466
rect 33906 5414 33918 5466
rect 33918 5414 33932 5466
rect 33956 5414 33970 5466
rect 33970 5414 33982 5466
rect 33982 5414 34012 5466
rect 34036 5414 34046 5466
rect 34046 5414 34092 5466
rect 33796 5412 33852 5414
rect 33876 5412 33932 5414
rect 33956 5412 34012 5414
rect 34036 5412 34092 5414
rect 37370 8880 37426 8936
rect 39270 10362 39326 10364
rect 39350 10362 39406 10364
rect 39430 10362 39486 10364
rect 39510 10362 39566 10364
rect 39270 10310 39316 10362
rect 39316 10310 39326 10362
rect 39350 10310 39380 10362
rect 39380 10310 39392 10362
rect 39392 10310 39406 10362
rect 39430 10310 39444 10362
rect 39444 10310 39456 10362
rect 39456 10310 39486 10362
rect 39510 10310 39520 10362
rect 39520 10310 39566 10362
rect 39270 10308 39326 10310
rect 39350 10308 39406 10310
rect 39430 10308 39486 10310
rect 39510 10308 39566 10310
rect 44743 17434 44799 17436
rect 44823 17434 44879 17436
rect 44903 17434 44959 17436
rect 44983 17434 45039 17436
rect 44743 17382 44789 17434
rect 44789 17382 44799 17434
rect 44823 17382 44853 17434
rect 44853 17382 44865 17434
rect 44865 17382 44879 17434
rect 44903 17382 44917 17434
rect 44917 17382 44929 17434
rect 44929 17382 44959 17434
rect 44983 17382 44993 17434
rect 44993 17382 45039 17434
rect 44743 17380 44799 17382
rect 44823 17380 44879 17382
rect 44903 17380 44959 17382
rect 44983 17380 45039 17382
rect 44743 16346 44799 16348
rect 44823 16346 44879 16348
rect 44903 16346 44959 16348
rect 44983 16346 45039 16348
rect 44743 16294 44789 16346
rect 44789 16294 44799 16346
rect 44823 16294 44853 16346
rect 44853 16294 44865 16346
rect 44865 16294 44879 16346
rect 44903 16294 44917 16346
rect 44917 16294 44929 16346
rect 44929 16294 44959 16346
rect 44983 16294 44993 16346
rect 44993 16294 45039 16346
rect 44743 16292 44799 16294
rect 44823 16292 44879 16294
rect 44903 16292 44959 16294
rect 44983 16292 45039 16294
rect 44362 15680 44418 15736
rect 44743 15258 44799 15260
rect 44823 15258 44879 15260
rect 44903 15258 44959 15260
rect 44983 15258 45039 15260
rect 44743 15206 44789 15258
rect 44789 15206 44799 15258
rect 44823 15206 44853 15258
rect 44853 15206 44865 15258
rect 44865 15206 44879 15258
rect 44903 15206 44917 15258
rect 44917 15206 44929 15258
rect 44929 15206 44959 15258
rect 44983 15206 44993 15258
rect 44993 15206 45039 15258
rect 44743 15204 44799 15206
rect 44823 15204 44879 15206
rect 44903 15204 44959 15206
rect 44983 15204 45039 15206
rect 45006 14340 45062 14376
rect 45006 14320 45008 14340
rect 45008 14320 45060 14340
rect 45060 14320 45062 14340
rect 44743 14170 44799 14172
rect 44823 14170 44879 14172
rect 44903 14170 44959 14172
rect 44983 14170 45039 14172
rect 44743 14118 44789 14170
rect 44789 14118 44799 14170
rect 44823 14118 44853 14170
rect 44853 14118 44865 14170
rect 44865 14118 44879 14170
rect 44903 14118 44917 14170
rect 44917 14118 44929 14170
rect 44929 14118 44959 14170
rect 44983 14118 44993 14170
rect 44993 14118 45039 14170
rect 44743 14116 44799 14118
rect 44823 14116 44879 14118
rect 44903 14116 44959 14118
rect 44983 14116 45039 14118
rect 41694 13948 41696 13968
rect 41696 13948 41748 13968
rect 41748 13948 41750 13968
rect 41694 13912 41750 13948
rect 41786 11736 41842 11792
rect 44743 13082 44799 13084
rect 44823 13082 44879 13084
rect 44903 13082 44959 13084
rect 44983 13082 45039 13084
rect 44743 13030 44789 13082
rect 44789 13030 44799 13082
rect 44823 13030 44853 13082
rect 44853 13030 44865 13082
rect 44865 13030 44879 13082
rect 44903 13030 44917 13082
rect 44917 13030 44929 13082
rect 44929 13030 44959 13082
rect 44983 13030 44993 13082
rect 44993 13030 45039 13082
rect 44743 13028 44799 13030
rect 44823 13028 44879 13030
rect 44903 13028 44959 13030
rect 44983 13028 45039 13030
rect 45006 12280 45062 12336
rect 44743 11994 44799 11996
rect 44823 11994 44879 11996
rect 44903 11994 44959 11996
rect 44983 11994 45039 11996
rect 44743 11942 44789 11994
rect 44789 11942 44799 11994
rect 44823 11942 44853 11994
rect 44853 11942 44865 11994
rect 44865 11942 44879 11994
rect 44903 11942 44917 11994
rect 44917 11942 44929 11994
rect 44929 11942 44959 11994
rect 44983 11942 44993 11994
rect 44993 11942 45039 11994
rect 44743 11940 44799 11942
rect 44823 11940 44879 11942
rect 44903 11940 44959 11942
rect 44983 11940 45039 11942
rect 45006 11092 45008 11112
rect 45008 11092 45060 11112
rect 45060 11092 45062 11112
rect 45006 11056 45062 11092
rect 39270 9274 39326 9276
rect 39350 9274 39406 9276
rect 39430 9274 39486 9276
rect 39510 9274 39566 9276
rect 39270 9222 39316 9274
rect 39316 9222 39326 9274
rect 39350 9222 39380 9274
rect 39380 9222 39392 9274
rect 39392 9222 39406 9274
rect 39430 9222 39444 9274
rect 39444 9222 39456 9274
rect 39456 9222 39486 9274
rect 39510 9222 39520 9274
rect 39520 9222 39566 9274
rect 39270 9220 39326 9222
rect 39350 9220 39406 9222
rect 39430 9220 39486 9222
rect 39510 9220 39566 9222
rect 39210 8900 39266 8936
rect 39210 8880 39212 8900
rect 39212 8880 39264 8900
rect 39264 8880 39266 8900
rect 38474 8336 38530 8392
rect 36910 6840 36966 6896
rect 37094 6024 37150 6080
rect 36910 5636 36966 5672
rect 36910 5616 36912 5636
rect 36912 5616 36964 5636
rect 36964 5616 36966 5636
rect 40314 8916 40316 8936
rect 40316 8916 40368 8936
rect 40368 8916 40370 8936
rect 40314 8880 40370 8916
rect 39270 8186 39326 8188
rect 39350 8186 39406 8188
rect 39430 8186 39486 8188
rect 39510 8186 39566 8188
rect 39270 8134 39316 8186
rect 39316 8134 39326 8186
rect 39350 8134 39380 8186
rect 39380 8134 39392 8186
rect 39392 8134 39406 8186
rect 39430 8134 39444 8186
rect 39444 8134 39456 8186
rect 39456 8134 39486 8186
rect 39510 8134 39520 8186
rect 39520 8134 39566 8186
rect 39270 8132 39326 8134
rect 39350 8132 39406 8134
rect 39430 8132 39486 8134
rect 39510 8132 39566 8134
rect 39270 7098 39326 7100
rect 39350 7098 39406 7100
rect 39430 7098 39486 7100
rect 39510 7098 39566 7100
rect 39270 7046 39316 7098
rect 39316 7046 39326 7098
rect 39350 7046 39380 7098
rect 39380 7046 39392 7098
rect 39392 7046 39406 7098
rect 39430 7046 39444 7098
rect 39444 7046 39456 7098
rect 39456 7046 39486 7098
rect 39510 7046 39520 7098
rect 39520 7046 39566 7098
rect 39270 7044 39326 7046
rect 39350 7044 39406 7046
rect 39430 7044 39486 7046
rect 39510 7044 39566 7046
rect 39270 6010 39326 6012
rect 39350 6010 39406 6012
rect 39430 6010 39486 6012
rect 39510 6010 39566 6012
rect 39270 5958 39316 6010
rect 39316 5958 39326 6010
rect 39350 5958 39380 6010
rect 39380 5958 39392 6010
rect 39392 5958 39406 6010
rect 39430 5958 39444 6010
rect 39444 5958 39456 6010
rect 39456 5958 39486 6010
rect 39510 5958 39520 6010
rect 39520 5958 39566 6010
rect 39270 5956 39326 5958
rect 39350 5956 39406 5958
rect 39430 5956 39486 5958
rect 39510 5956 39566 5958
rect 44743 10906 44799 10908
rect 44823 10906 44879 10908
rect 44903 10906 44959 10908
rect 44983 10906 45039 10908
rect 44743 10854 44789 10906
rect 44789 10854 44799 10906
rect 44823 10854 44853 10906
rect 44853 10854 44865 10906
rect 44865 10854 44879 10906
rect 44903 10854 44917 10906
rect 44917 10854 44929 10906
rect 44929 10854 44959 10906
rect 44983 10854 44993 10906
rect 44993 10854 45039 10906
rect 44743 10852 44799 10854
rect 44823 10852 44879 10854
rect 44903 10852 44959 10854
rect 44983 10852 45039 10854
rect 44743 9818 44799 9820
rect 44823 9818 44879 9820
rect 44903 9818 44959 9820
rect 44983 9818 45039 9820
rect 44743 9766 44789 9818
rect 44789 9766 44799 9818
rect 44823 9766 44853 9818
rect 44853 9766 44865 9818
rect 44865 9766 44879 9818
rect 44903 9766 44917 9818
rect 44917 9766 44929 9818
rect 44929 9766 44959 9818
rect 44983 9766 44993 9818
rect 44993 9766 45039 9818
rect 44743 9764 44799 9766
rect 44823 9764 44879 9766
rect 44903 9764 44959 9766
rect 44983 9764 45039 9766
rect 44362 8880 44418 8936
rect 44743 8730 44799 8732
rect 44823 8730 44879 8732
rect 44903 8730 44959 8732
rect 44983 8730 45039 8732
rect 44743 8678 44789 8730
rect 44789 8678 44799 8730
rect 44823 8678 44853 8730
rect 44853 8678 44865 8730
rect 44865 8678 44879 8730
rect 44903 8678 44917 8730
rect 44917 8678 44929 8730
rect 44929 8678 44959 8730
rect 44983 8678 44993 8730
rect 44993 8678 45039 8730
rect 44743 8676 44799 8678
rect 44823 8676 44879 8678
rect 44903 8676 44959 8678
rect 44983 8676 45039 8678
rect 44362 7828 44364 7848
rect 44364 7828 44416 7848
rect 44416 7828 44418 7848
rect 44362 7792 44418 7828
rect 44743 7642 44799 7644
rect 44823 7642 44879 7644
rect 44903 7642 44959 7644
rect 44983 7642 45039 7644
rect 44743 7590 44789 7642
rect 44789 7590 44799 7642
rect 44823 7590 44853 7642
rect 44853 7590 44865 7642
rect 44865 7590 44879 7642
rect 44903 7590 44917 7642
rect 44917 7590 44929 7642
rect 44929 7590 44959 7642
rect 44983 7590 44993 7642
rect 44993 7590 45039 7642
rect 44743 7588 44799 7590
rect 44823 7588 44879 7590
rect 44903 7588 44959 7590
rect 44983 7588 45039 7590
rect 44743 6554 44799 6556
rect 44823 6554 44879 6556
rect 44903 6554 44959 6556
rect 44983 6554 45039 6556
rect 44743 6502 44789 6554
rect 44789 6502 44799 6554
rect 44823 6502 44853 6554
rect 44853 6502 44865 6554
rect 44865 6502 44879 6554
rect 44903 6502 44917 6554
rect 44917 6502 44929 6554
rect 44929 6502 44959 6554
rect 44983 6502 44993 6554
rect 44993 6502 45039 6554
rect 44743 6500 44799 6502
rect 44823 6500 44879 6502
rect 44903 6500 44959 6502
rect 44983 6500 45039 6502
rect 41970 6160 42026 6216
rect 41418 5228 41474 5264
rect 41418 5208 41420 5228
rect 41420 5208 41472 5228
rect 41472 5208 41474 5228
rect 42798 5072 42854 5128
rect 39270 4922 39326 4924
rect 39350 4922 39406 4924
rect 39430 4922 39486 4924
rect 39510 4922 39566 4924
rect 39270 4870 39316 4922
rect 39316 4870 39326 4922
rect 39350 4870 39380 4922
rect 39380 4870 39392 4922
rect 39392 4870 39406 4922
rect 39430 4870 39444 4922
rect 39444 4870 39456 4922
rect 39456 4870 39486 4922
rect 39510 4870 39520 4922
rect 39520 4870 39566 4922
rect 39270 4868 39326 4870
rect 39350 4868 39406 4870
rect 39430 4868 39486 4870
rect 39510 4868 39566 4870
rect 33796 4378 33852 4380
rect 33876 4378 33932 4380
rect 33956 4378 34012 4380
rect 34036 4378 34092 4380
rect 33796 4326 33842 4378
rect 33842 4326 33852 4378
rect 33876 4326 33906 4378
rect 33906 4326 33918 4378
rect 33918 4326 33932 4378
rect 33956 4326 33970 4378
rect 33970 4326 33982 4378
rect 33982 4326 34012 4378
rect 34036 4326 34046 4378
rect 34046 4326 34092 4378
rect 33796 4324 33852 4326
rect 33876 4324 33932 4326
rect 33956 4324 34012 4326
rect 34036 4324 34092 4326
rect 33796 3290 33852 3292
rect 33876 3290 33932 3292
rect 33956 3290 34012 3292
rect 34036 3290 34092 3292
rect 33796 3238 33842 3290
rect 33842 3238 33852 3290
rect 33876 3238 33906 3290
rect 33906 3238 33918 3290
rect 33918 3238 33932 3290
rect 33956 3238 33970 3290
rect 33970 3238 33982 3290
rect 33982 3238 34012 3290
rect 34036 3238 34046 3290
rect 34046 3238 34092 3290
rect 33796 3236 33852 3238
rect 33876 3236 33932 3238
rect 33956 3236 34012 3238
rect 34036 3236 34092 3238
rect 33796 2202 33852 2204
rect 33876 2202 33932 2204
rect 33956 2202 34012 2204
rect 34036 2202 34092 2204
rect 33796 2150 33842 2202
rect 33842 2150 33852 2202
rect 33876 2150 33906 2202
rect 33906 2150 33918 2202
rect 33918 2150 33932 2202
rect 33956 2150 33970 2202
rect 33970 2150 33982 2202
rect 33982 2150 34012 2202
rect 34036 2150 34046 2202
rect 34046 2150 34092 2202
rect 33796 2148 33852 2150
rect 33876 2148 33932 2150
rect 33956 2148 34012 2150
rect 34036 2148 34092 2150
rect 39270 3834 39326 3836
rect 39350 3834 39406 3836
rect 39430 3834 39486 3836
rect 39510 3834 39566 3836
rect 39270 3782 39316 3834
rect 39316 3782 39326 3834
rect 39350 3782 39380 3834
rect 39380 3782 39392 3834
rect 39392 3782 39406 3834
rect 39430 3782 39444 3834
rect 39444 3782 39456 3834
rect 39456 3782 39486 3834
rect 39510 3782 39520 3834
rect 39520 3782 39566 3834
rect 39270 3780 39326 3782
rect 39350 3780 39406 3782
rect 39430 3780 39486 3782
rect 39510 3780 39566 3782
rect 39270 2746 39326 2748
rect 39350 2746 39406 2748
rect 39430 2746 39486 2748
rect 39510 2746 39566 2748
rect 39270 2694 39316 2746
rect 39316 2694 39326 2746
rect 39350 2694 39380 2746
rect 39380 2694 39392 2746
rect 39392 2694 39406 2746
rect 39430 2694 39444 2746
rect 39444 2694 39456 2746
rect 39456 2694 39486 2746
rect 39510 2694 39520 2746
rect 39520 2694 39566 2746
rect 39270 2692 39326 2694
rect 39350 2692 39406 2694
rect 39430 2692 39486 2694
rect 39510 2692 39566 2694
rect 44743 5466 44799 5468
rect 44823 5466 44879 5468
rect 44903 5466 44959 5468
rect 44983 5466 45039 5468
rect 44743 5414 44789 5466
rect 44789 5414 44799 5466
rect 44823 5414 44853 5466
rect 44853 5414 44865 5466
rect 44865 5414 44879 5466
rect 44903 5414 44917 5466
rect 44917 5414 44929 5466
rect 44929 5414 44959 5466
rect 44983 5414 44993 5466
rect 44993 5414 45039 5466
rect 44743 5412 44799 5414
rect 44823 5412 44879 5414
rect 44903 5412 44959 5414
rect 44983 5412 45039 5414
rect 44743 4378 44799 4380
rect 44823 4378 44879 4380
rect 44903 4378 44959 4380
rect 44983 4378 45039 4380
rect 44743 4326 44789 4378
rect 44789 4326 44799 4378
rect 44823 4326 44853 4378
rect 44853 4326 44865 4378
rect 44865 4326 44879 4378
rect 44903 4326 44917 4378
rect 44917 4326 44929 4378
rect 44929 4326 44959 4378
rect 44983 4326 44993 4378
rect 44993 4326 45039 4378
rect 44743 4324 44799 4326
rect 44823 4324 44879 4326
rect 44903 4324 44959 4326
rect 44983 4324 45039 4326
rect 44638 4120 44694 4176
rect 41418 2352 41474 2408
rect 44743 3290 44799 3292
rect 44823 3290 44879 3292
rect 44903 3290 44959 3292
rect 44983 3290 45039 3292
rect 44743 3238 44789 3290
rect 44789 3238 44799 3290
rect 44823 3238 44853 3290
rect 44853 3238 44865 3290
rect 44865 3238 44879 3290
rect 44903 3238 44917 3290
rect 44917 3238 44929 3290
rect 44929 3238 44959 3290
rect 44983 3238 44993 3290
rect 44993 3238 45039 3290
rect 44743 3236 44799 3238
rect 44823 3236 44879 3238
rect 44903 3236 44959 3238
rect 44983 3236 45039 3238
rect 44743 2202 44799 2204
rect 44823 2202 44879 2204
rect 44903 2202 44959 2204
rect 44983 2202 45039 2204
rect 44743 2150 44789 2202
rect 44789 2150 44799 2202
rect 44823 2150 44853 2202
rect 44853 2150 44865 2202
rect 44865 2150 44879 2202
rect 44903 2150 44917 2202
rect 44917 2150 44929 2202
rect 44929 2150 44959 2202
rect 44983 2150 44993 2202
rect 44993 2150 45039 2202
rect 44743 2148 44799 2150
rect 44823 2148 44879 2150
rect 44903 2148 44959 2150
rect 44983 2148 45039 2150
rect 44638 720 44694 776
<< metal3 >>
rect 45001 19138 45067 19141
rect 45200 19138 46000 19228
rect 45001 19136 46000 19138
rect 45001 19080 45006 19136
rect 45062 19080 46000 19136
rect 45001 19078 46000 19080
rect 45001 19075 45067 19078
rect 45200 18988 46000 19078
rect 0 18458 800 18548
rect 1025 18458 1091 18461
rect 0 18456 1091 18458
rect 0 18400 1030 18456
rect 1086 18400 1091 18456
rect 0 18398 1091 18400
rect 0 18308 800 18398
rect 1025 18395 1091 18398
rect 45001 17778 45067 17781
rect 45200 17778 46000 17868
rect 45001 17776 46000 17778
rect 45001 17720 45006 17776
rect 45062 17720 46000 17776
rect 45001 17718 46000 17720
rect 45001 17715 45067 17718
rect 45200 17628 46000 17718
rect 11892 17440 12208 17441
rect 11892 17376 11898 17440
rect 11962 17376 11978 17440
rect 12042 17376 12058 17440
rect 12122 17376 12138 17440
rect 12202 17376 12208 17440
rect 11892 17375 12208 17376
rect 22839 17440 23155 17441
rect 22839 17376 22845 17440
rect 22909 17376 22925 17440
rect 22989 17376 23005 17440
rect 23069 17376 23085 17440
rect 23149 17376 23155 17440
rect 22839 17375 23155 17376
rect 33786 17440 34102 17441
rect 33786 17376 33792 17440
rect 33856 17376 33872 17440
rect 33936 17376 33952 17440
rect 34016 17376 34032 17440
rect 34096 17376 34102 17440
rect 33786 17375 34102 17376
rect 44733 17440 45049 17441
rect 44733 17376 44739 17440
rect 44803 17376 44819 17440
rect 44883 17376 44899 17440
rect 44963 17376 44979 17440
rect 45043 17376 45049 17440
rect 44733 17375 45049 17376
rect 0 17098 800 17188
rect 933 17098 999 17101
rect 0 17096 999 17098
rect 0 17040 938 17096
rect 994 17040 999 17096
rect 0 17038 999 17040
rect 0 16948 800 17038
rect 933 17035 999 17038
rect 6419 16896 6735 16897
rect 6419 16832 6425 16896
rect 6489 16832 6505 16896
rect 6569 16832 6585 16896
rect 6649 16832 6665 16896
rect 6729 16832 6735 16896
rect 6419 16831 6735 16832
rect 17366 16896 17682 16897
rect 17366 16832 17372 16896
rect 17436 16832 17452 16896
rect 17516 16832 17532 16896
rect 17596 16832 17612 16896
rect 17676 16832 17682 16896
rect 17366 16831 17682 16832
rect 28313 16896 28629 16897
rect 28313 16832 28319 16896
rect 28383 16832 28399 16896
rect 28463 16832 28479 16896
rect 28543 16832 28559 16896
rect 28623 16832 28629 16896
rect 28313 16831 28629 16832
rect 39260 16896 39576 16897
rect 39260 16832 39266 16896
rect 39330 16832 39346 16896
rect 39410 16832 39426 16896
rect 39490 16832 39506 16896
rect 39570 16832 39576 16896
rect 39260 16831 39576 16832
rect 11892 16352 12208 16353
rect 11892 16288 11898 16352
rect 11962 16288 11978 16352
rect 12042 16288 12058 16352
rect 12122 16288 12138 16352
rect 12202 16288 12208 16352
rect 11892 16287 12208 16288
rect 22839 16352 23155 16353
rect 22839 16288 22845 16352
rect 22909 16288 22925 16352
rect 22989 16288 23005 16352
rect 23069 16288 23085 16352
rect 23149 16288 23155 16352
rect 22839 16287 23155 16288
rect 33786 16352 34102 16353
rect 33786 16288 33792 16352
rect 33856 16288 33872 16352
rect 33936 16288 33952 16352
rect 34016 16288 34032 16352
rect 34096 16288 34102 16352
rect 33786 16287 34102 16288
rect 44733 16352 45049 16353
rect 44733 16288 44739 16352
rect 44803 16288 44819 16352
rect 44883 16288 44899 16352
rect 44963 16288 44979 16352
rect 45043 16288 45049 16352
rect 44733 16287 45049 16288
rect 6419 15808 6735 15809
rect 6419 15744 6425 15808
rect 6489 15744 6505 15808
rect 6569 15744 6585 15808
rect 6649 15744 6665 15808
rect 6729 15744 6735 15808
rect 6419 15743 6735 15744
rect 17366 15808 17682 15809
rect 17366 15744 17372 15808
rect 17436 15744 17452 15808
rect 17516 15744 17532 15808
rect 17596 15744 17612 15808
rect 17676 15744 17682 15808
rect 17366 15743 17682 15744
rect 28313 15808 28629 15809
rect 28313 15744 28319 15808
rect 28383 15744 28399 15808
rect 28463 15744 28479 15808
rect 28543 15744 28559 15808
rect 28623 15744 28629 15808
rect 28313 15743 28629 15744
rect 39260 15808 39576 15809
rect 39260 15744 39266 15808
rect 39330 15744 39346 15808
rect 39410 15744 39426 15808
rect 39490 15744 39506 15808
rect 39570 15744 39576 15808
rect 39260 15743 39576 15744
rect 44357 15738 44423 15741
rect 45200 15738 46000 15828
rect 44357 15736 46000 15738
rect 44357 15680 44362 15736
rect 44418 15680 46000 15736
rect 44357 15678 46000 15680
rect 44357 15675 44423 15678
rect 45200 15588 46000 15678
rect 11892 15264 12208 15265
rect 11892 15200 11898 15264
rect 11962 15200 11978 15264
rect 12042 15200 12058 15264
rect 12122 15200 12138 15264
rect 12202 15200 12208 15264
rect 11892 15199 12208 15200
rect 22839 15264 23155 15265
rect 22839 15200 22845 15264
rect 22909 15200 22925 15264
rect 22989 15200 23005 15264
rect 23069 15200 23085 15264
rect 23149 15200 23155 15264
rect 22839 15199 23155 15200
rect 33786 15264 34102 15265
rect 33786 15200 33792 15264
rect 33856 15200 33872 15264
rect 33936 15200 33952 15264
rect 34016 15200 34032 15264
rect 34096 15200 34102 15264
rect 33786 15199 34102 15200
rect 44733 15264 45049 15265
rect 44733 15200 44739 15264
rect 44803 15200 44819 15264
rect 44883 15200 44899 15264
rect 44963 15200 44979 15264
rect 45043 15200 45049 15264
rect 44733 15199 45049 15200
rect 0 15058 800 15148
rect 1025 15058 1091 15061
rect 0 15056 1091 15058
rect 0 15000 1030 15056
rect 1086 15000 1091 15056
rect 0 14998 1091 15000
rect 0 14908 800 14998
rect 1025 14995 1091 14998
rect 6419 14720 6735 14721
rect 6419 14656 6425 14720
rect 6489 14656 6505 14720
rect 6569 14656 6585 14720
rect 6649 14656 6665 14720
rect 6729 14656 6735 14720
rect 6419 14655 6735 14656
rect 17366 14720 17682 14721
rect 17366 14656 17372 14720
rect 17436 14656 17452 14720
rect 17516 14656 17532 14720
rect 17596 14656 17612 14720
rect 17676 14656 17682 14720
rect 17366 14655 17682 14656
rect 28313 14720 28629 14721
rect 28313 14656 28319 14720
rect 28383 14656 28399 14720
rect 28463 14656 28479 14720
rect 28543 14656 28559 14720
rect 28623 14656 28629 14720
rect 28313 14655 28629 14656
rect 39260 14720 39576 14721
rect 39260 14656 39266 14720
rect 39330 14656 39346 14720
rect 39410 14656 39426 14720
rect 39490 14656 39506 14720
rect 39570 14656 39576 14720
rect 39260 14655 39576 14656
rect 23657 14378 23723 14381
rect 38837 14378 38903 14381
rect 23657 14376 38903 14378
rect 23657 14320 23662 14376
rect 23718 14320 38842 14376
rect 38898 14320 38903 14376
rect 23657 14318 38903 14320
rect 23657 14315 23723 14318
rect 38837 14315 38903 14318
rect 45001 14378 45067 14381
rect 45200 14378 46000 14468
rect 45001 14376 46000 14378
rect 45001 14320 45006 14376
rect 45062 14320 46000 14376
rect 45001 14318 46000 14320
rect 45001 14315 45067 14318
rect 45200 14228 46000 14318
rect 11892 14176 12208 14177
rect 11892 14112 11898 14176
rect 11962 14112 11978 14176
rect 12042 14112 12058 14176
rect 12122 14112 12138 14176
rect 12202 14112 12208 14176
rect 11892 14111 12208 14112
rect 22839 14176 23155 14177
rect 22839 14112 22845 14176
rect 22909 14112 22925 14176
rect 22989 14112 23005 14176
rect 23069 14112 23085 14176
rect 23149 14112 23155 14176
rect 22839 14111 23155 14112
rect 33786 14176 34102 14177
rect 33786 14112 33792 14176
rect 33856 14112 33872 14176
rect 33936 14112 33952 14176
rect 34016 14112 34032 14176
rect 34096 14112 34102 14176
rect 33786 14111 34102 14112
rect 44733 14176 45049 14177
rect 44733 14112 44739 14176
rect 44803 14112 44819 14176
rect 44883 14112 44899 14176
rect 44963 14112 44979 14176
rect 45043 14112 45049 14176
rect 44733 14111 45049 14112
rect 16573 13970 16639 13973
rect 41689 13970 41755 13973
rect 16573 13968 41755 13970
rect 16573 13912 16578 13968
rect 16634 13912 41694 13968
rect 41750 13912 41755 13968
rect 16573 13910 41755 13912
rect 16573 13907 16639 13910
rect 41689 13907 41755 13910
rect 0 13698 800 13788
rect 933 13698 999 13701
rect 0 13696 999 13698
rect 0 13640 938 13696
rect 994 13640 999 13696
rect 0 13638 999 13640
rect 0 13548 800 13638
rect 933 13635 999 13638
rect 6419 13632 6735 13633
rect 6419 13568 6425 13632
rect 6489 13568 6505 13632
rect 6569 13568 6585 13632
rect 6649 13568 6665 13632
rect 6729 13568 6735 13632
rect 6419 13567 6735 13568
rect 17366 13632 17682 13633
rect 17366 13568 17372 13632
rect 17436 13568 17452 13632
rect 17516 13568 17532 13632
rect 17596 13568 17612 13632
rect 17676 13568 17682 13632
rect 17366 13567 17682 13568
rect 28313 13632 28629 13633
rect 28313 13568 28319 13632
rect 28383 13568 28399 13632
rect 28463 13568 28479 13632
rect 28543 13568 28559 13632
rect 28623 13568 28629 13632
rect 28313 13567 28629 13568
rect 39260 13632 39576 13633
rect 39260 13568 39266 13632
rect 39330 13568 39346 13632
rect 39410 13568 39426 13632
rect 39490 13568 39506 13632
rect 39570 13568 39576 13632
rect 39260 13567 39576 13568
rect 11892 13088 12208 13089
rect 11892 13024 11898 13088
rect 11962 13024 11978 13088
rect 12042 13024 12058 13088
rect 12122 13024 12138 13088
rect 12202 13024 12208 13088
rect 11892 13023 12208 13024
rect 22839 13088 23155 13089
rect 22839 13024 22845 13088
rect 22909 13024 22925 13088
rect 22989 13024 23005 13088
rect 23069 13024 23085 13088
rect 23149 13024 23155 13088
rect 22839 13023 23155 13024
rect 33786 13088 34102 13089
rect 33786 13024 33792 13088
rect 33856 13024 33872 13088
rect 33936 13024 33952 13088
rect 34016 13024 34032 13088
rect 34096 13024 34102 13088
rect 33786 13023 34102 13024
rect 44733 13088 45049 13089
rect 44733 13024 44739 13088
rect 44803 13024 44819 13088
rect 44883 13024 44899 13088
rect 44963 13024 44979 13088
rect 45043 13024 45049 13088
rect 44733 13023 45049 13024
rect 6419 12544 6735 12545
rect 6419 12480 6425 12544
rect 6489 12480 6505 12544
rect 6569 12480 6585 12544
rect 6649 12480 6665 12544
rect 6729 12480 6735 12544
rect 6419 12479 6735 12480
rect 17366 12544 17682 12545
rect 17366 12480 17372 12544
rect 17436 12480 17452 12544
rect 17516 12480 17532 12544
rect 17596 12480 17612 12544
rect 17676 12480 17682 12544
rect 17366 12479 17682 12480
rect 28313 12544 28629 12545
rect 28313 12480 28319 12544
rect 28383 12480 28399 12544
rect 28463 12480 28479 12544
rect 28543 12480 28559 12544
rect 28623 12480 28629 12544
rect 28313 12479 28629 12480
rect 39260 12544 39576 12545
rect 39260 12480 39266 12544
rect 39330 12480 39346 12544
rect 39410 12480 39426 12544
rect 39490 12480 39506 12544
rect 39570 12480 39576 12544
rect 39260 12479 39576 12480
rect 45001 12338 45067 12341
rect 45200 12338 46000 12428
rect 45001 12336 46000 12338
rect 45001 12280 45006 12336
rect 45062 12280 46000 12336
rect 45001 12278 46000 12280
rect 45001 12275 45067 12278
rect 2129 12202 2195 12205
rect 31017 12202 31083 12205
rect 2129 12200 31083 12202
rect 2129 12144 2134 12200
rect 2190 12144 31022 12200
rect 31078 12144 31083 12200
rect 45200 12188 46000 12278
rect 2129 12142 31083 12144
rect 2129 12139 2195 12142
rect 31017 12139 31083 12142
rect 11892 12000 12208 12001
rect 11892 11936 11898 12000
rect 11962 11936 11978 12000
rect 12042 11936 12058 12000
rect 12122 11936 12138 12000
rect 12202 11936 12208 12000
rect 11892 11935 12208 11936
rect 22839 12000 23155 12001
rect 22839 11936 22845 12000
rect 22909 11936 22925 12000
rect 22989 11936 23005 12000
rect 23069 11936 23085 12000
rect 23149 11936 23155 12000
rect 22839 11935 23155 11936
rect 33786 12000 34102 12001
rect 33786 11936 33792 12000
rect 33856 11936 33872 12000
rect 33936 11936 33952 12000
rect 34016 11936 34032 12000
rect 34096 11936 34102 12000
rect 33786 11935 34102 11936
rect 44733 12000 45049 12001
rect 44733 11936 44739 12000
rect 44803 11936 44819 12000
rect 44883 11936 44899 12000
rect 44963 11936 44979 12000
rect 45043 11936 45049 12000
rect 44733 11935 45049 11936
rect 6913 11794 6979 11797
rect 41781 11794 41847 11797
rect 6913 11792 41847 11794
rect 0 11658 800 11748
rect 6913 11736 6918 11792
rect 6974 11736 41786 11792
rect 41842 11736 41847 11792
rect 6913 11734 41847 11736
rect 6913 11731 6979 11734
rect 41781 11731 41847 11734
rect 4061 11658 4127 11661
rect 0 11656 4127 11658
rect 0 11600 4066 11656
rect 4122 11600 4127 11656
rect 0 11598 4127 11600
rect 0 11508 800 11598
rect 4061 11595 4127 11598
rect 6419 11456 6735 11457
rect 6419 11392 6425 11456
rect 6489 11392 6505 11456
rect 6569 11392 6585 11456
rect 6649 11392 6665 11456
rect 6729 11392 6735 11456
rect 6419 11391 6735 11392
rect 17366 11456 17682 11457
rect 17366 11392 17372 11456
rect 17436 11392 17452 11456
rect 17516 11392 17532 11456
rect 17596 11392 17612 11456
rect 17676 11392 17682 11456
rect 17366 11391 17682 11392
rect 28313 11456 28629 11457
rect 28313 11392 28319 11456
rect 28383 11392 28399 11456
rect 28463 11392 28479 11456
rect 28543 11392 28559 11456
rect 28623 11392 28629 11456
rect 28313 11391 28629 11392
rect 39260 11456 39576 11457
rect 39260 11392 39266 11456
rect 39330 11392 39346 11456
rect 39410 11392 39426 11456
rect 39490 11392 39506 11456
rect 39570 11392 39576 11456
rect 39260 11391 39576 11392
rect 27889 11114 27955 11117
rect 35065 11114 35131 11117
rect 27889 11112 35131 11114
rect 27889 11056 27894 11112
rect 27950 11056 35070 11112
rect 35126 11056 35131 11112
rect 27889 11054 35131 11056
rect 27889 11051 27955 11054
rect 35065 11051 35131 11054
rect 45001 11114 45067 11117
rect 45001 11112 45202 11114
rect 45001 11056 45006 11112
rect 45062 11068 45202 11112
rect 45062 11056 46000 11068
rect 45001 11054 46000 11056
rect 45001 11051 45067 11054
rect 45142 10918 46000 11054
rect 11892 10912 12208 10913
rect 11892 10848 11898 10912
rect 11962 10848 11978 10912
rect 12042 10848 12058 10912
rect 12122 10848 12138 10912
rect 12202 10848 12208 10912
rect 11892 10847 12208 10848
rect 22839 10912 23155 10913
rect 22839 10848 22845 10912
rect 22909 10848 22925 10912
rect 22989 10848 23005 10912
rect 23069 10848 23085 10912
rect 23149 10848 23155 10912
rect 22839 10847 23155 10848
rect 33786 10912 34102 10913
rect 33786 10848 33792 10912
rect 33856 10848 33872 10912
rect 33936 10848 33952 10912
rect 34016 10848 34032 10912
rect 34096 10848 34102 10912
rect 33786 10847 34102 10848
rect 44733 10912 45049 10913
rect 44733 10848 44739 10912
rect 44803 10848 44819 10912
rect 44883 10848 44899 10912
rect 44963 10848 44979 10912
rect 45043 10848 45049 10912
rect 44733 10847 45049 10848
rect 45200 10828 46000 10918
rect 5349 10706 5415 10709
rect 28073 10706 28139 10709
rect 29085 10706 29151 10709
rect 5349 10704 29151 10706
rect 5349 10648 5354 10704
rect 5410 10648 28078 10704
rect 28134 10648 29090 10704
rect 29146 10648 29151 10704
rect 5349 10646 29151 10648
rect 5349 10643 5415 10646
rect 28073 10643 28139 10646
rect 29085 10643 29151 10646
rect 17953 10570 18019 10573
rect 23657 10570 23723 10573
rect 17953 10568 23723 10570
rect 17953 10512 17958 10568
rect 18014 10512 23662 10568
rect 23718 10512 23723 10568
rect 17953 10510 23723 10512
rect 17953 10507 18019 10510
rect 23657 10507 23723 10510
rect 0 10298 800 10388
rect 6419 10368 6735 10369
rect 6419 10304 6425 10368
rect 6489 10304 6505 10368
rect 6569 10304 6585 10368
rect 6649 10304 6665 10368
rect 6729 10304 6735 10368
rect 6419 10303 6735 10304
rect 17366 10368 17682 10369
rect 17366 10304 17372 10368
rect 17436 10304 17452 10368
rect 17516 10304 17532 10368
rect 17596 10304 17612 10368
rect 17676 10304 17682 10368
rect 17366 10303 17682 10304
rect 28313 10368 28629 10369
rect 28313 10304 28319 10368
rect 28383 10304 28399 10368
rect 28463 10304 28479 10368
rect 28543 10304 28559 10368
rect 28623 10304 28629 10368
rect 28313 10303 28629 10304
rect 39260 10368 39576 10369
rect 39260 10304 39266 10368
rect 39330 10304 39346 10368
rect 39410 10304 39426 10368
rect 39490 10304 39506 10368
rect 39570 10304 39576 10368
rect 39260 10303 39576 10304
rect 933 10298 999 10301
rect 0 10296 999 10298
rect 0 10240 938 10296
rect 994 10240 999 10296
rect 0 10238 999 10240
rect 0 10148 800 10238
rect 933 10235 999 10238
rect 19701 10026 19767 10029
rect 24761 10026 24827 10029
rect 19701 10024 24827 10026
rect 19701 9968 19706 10024
rect 19762 9968 24766 10024
rect 24822 9968 24827 10024
rect 19701 9966 24827 9968
rect 19701 9963 19767 9966
rect 24761 9963 24827 9966
rect 11892 9824 12208 9825
rect 11892 9760 11898 9824
rect 11962 9760 11978 9824
rect 12042 9760 12058 9824
rect 12122 9760 12138 9824
rect 12202 9760 12208 9824
rect 11892 9759 12208 9760
rect 22839 9824 23155 9825
rect 22839 9760 22845 9824
rect 22909 9760 22925 9824
rect 22989 9760 23005 9824
rect 23069 9760 23085 9824
rect 23149 9760 23155 9824
rect 22839 9759 23155 9760
rect 33786 9824 34102 9825
rect 33786 9760 33792 9824
rect 33856 9760 33872 9824
rect 33936 9760 33952 9824
rect 34016 9760 34032 9824
rect 34096 9760 34102 9824
rect 33786 9759 34102 9760
rect 44733 9824 45049 9825
rect 44733 9760 44739 9824
rect 44803 9760 44819 9824
rect 44883 9760 44899 9824
rect 44963 9760 44979 9824
rect 45043 9760 45049 9824
rect 44733 9759 45049 9760
rect 22001 9754 22067 9757
rect 22277 9754 22343 9757
rect 22001 9752 22343 9754
rect 22001 9696 22006 9752
rect 22062 9696 22282 9752
rect 22338 9696 22343 9752
rect 22001 9694 22343 9696
rect 22001 9691 22067 9694
rect 22277 9691 22343 9694
rect 23841 9618 23907 9621
rect 27889 9618 27955 9621
rect 23841 9616 27955 9618
rect 23841 9560 23846 9616
rect 23902 9560 27894 9616
rect 27950 9560 27955 9616
rect 23841 9558 27955 9560
rect 23841 9555 23907 9558
rect 27889 9555 27955 9558
rect 1761 9482 1827 9485
rect 32857 9482 32923 9485
rect 1761 9480 32923 9482
rect 1761 9424 1766 9480
rect 1822 9424 32862 9480
rect 32918 9424 32923 9480
rect 1761 9422 32923 9424
rect 1761 9419 1827 9422
rect 32857 9419 32923 9422
rect 6419 9280 6735 9281
rect 6419 9216 6425 9280
rect 6489 9216 6505 9280
rect 6569 9216 6585 9280
rect 6649 9216 6665 9280
rect 6729 9216 6735 9280
rect 6419 9215 6735 9216
rect 17366 9280 17682 9281
rect 17366 9216 17372 9280
rect 17436 9216 17452 9280
rect 17516 9216 17532 9280
rect 17596 9216 17612 9280
rect 17676 9216 17682 9280
rect 17366 9215 17682 9216
rect 28313 9280 28629 9281
rect 28313 9216 28319 9280
rect 28383 9216 28399 9280
rect 28463 9216 28479 9280
rect 28543 9216 28559 9280
rect 28623 9216 28629 9280
rect 28313 9215 28629 9216
rect 39260 9280 39576 9281
rect 39260 9216 39266 9280
rect 39330 9216 39346 9280
rect 39410 9216 39426 9280
rect 39490 9216 39506 9280
rect 39570 9216 39576 9280
rect 39260 9215 39576 9216
rect 30097 8938 30163 8941
rect 32489 8938 32555 8941
rect 37365 8938 37431 8941
rect 30097 8936 37431 8938
rect 30097 8880 30102 8936
rect 30158 8880 32494 8936
rect 32550 8880 37370 8936
rect 37426 8880 37431 8936
rect 30097 8878 37431 8880
rect 30097 8875 30163 8878
rect 32489 8875 32555 8878
rect 37365 8875 37431 8878
rect 39205 8938 39271 8941
rect 40309 8938 40375 8941
rect 39205 8936 40375 8938
rect 39205 8880 39210 8936
rect 39266 8880 40314 8936
rect 40370 8880 40375 8936
rect 39205 8878 40375 8880
rect 39205 8875 39271 8878
rect 40309 8875 40375 8878
rect 44357 8938 44423 8941
rect 45200 8938 46000 9028
rect 44357 8936 46000 8938
rect 44357 8880 44362 8936
rect 44418 8880 46000 8936
rect 44357 8878 46000 8880
rect 44357 8875 44423 8878
rect 45200 8788 46000 8878
rect 11892 8736 12208 8737
rect 11892 8672 11898 8736
rect 11962 8672 11978 8736
rect 12042 8672 12058 8736
rect 12122 8672 12138 8736
rect 12202 8672 12208 8736
rect 11892 8671 12208 8672
rect 22839 8736 23155 8737
rect 22839 8672 22845 8736
rect 22909 8672 22925 8736
rect 22989 8672 23005 8736
rect 23069 8672 23085 8736
rect 23149 8672 23155 8736
rect 22839 8671 23155 8672
rect 33786 8736 34102 8737
rect 33786 8672 33792 8736
rect 33856 8672 33872 8736
rect 33936 8672 33952 8736
rect 34016 8672 34032 8736
rect 34096 8672 34102 8736
rect 33786 8671 34102 8672
rect 44733 8736 45049 8737
rect 44733 8672 44739 8736
rect 44803 8672 44819 8736
rect 44883 8672 44899 8736
rect 44963 8672 44979 8736
rect 45043 8672 45049 8736
rect 44733 8671 45049 8672
rect 3601 8530 3667 8533
rect 34513 8530 34579 8533
rect 3601 8528 34579 8530
rect 3601 8472 3606 8528
rect 3662 8472 34518 8528
rect 34574 8472 34579 8528
rect 3601 8470 34579 8472
rect 3601 8467 3667 8470
rect 34513 8467 34579 8470
rect 33409 8394 33475 8397
rect 38469 8394 38535 8397
rect 33409 8392 38535 8394
rect 0 8258 800 8348
rect 33409 8336 33414 8392
rect 33470 8336 38474 8392
rect 38530 8336 38535 8392
rect 33409 8334 38535 8336
rect 33409 8331 33475 8334
rect 38469 8331 38535 8334
rect 933 8258 999 8261
rect 0 8256 999 8258
rect 0 8200 938 8256
rect 994 8200 999 8256
rect 0 8198 999 8200
rect 0 8108 800 8198
rect 933 8195 999 8198
rect 6419 8192 6735 8193
rect 6419 8128 6425 8192
rect 6489 8128 6505 8192
rect 6569 8128 6585 8192
rect 6649 8128 6665 8192
rect 6729 8128 6735 8192
rect 6419 8127 6735 8128
rect 17366 8192 17682 8193
rect 17366 8128 17372 8192
rect 17436 8128 17452 8192
rect 17516 8128 17532 8192
rect 17596 8128 17612 8192
rect 17676 8128 17682 8192
rect 17366 8127 17682 8128
rect 28313 8192 28629 8193
rect 28313 8128 28319 8192
rect 28383 8128 28399 8192
rect 28463 8128 28479 8192
rect 28543 8128 28559 8192
rect 28623 8128 28629 8192
rect 28313 8127 28629 8128
rect 39260 8192 39576 8193
rect 39260 8128 39266 8192
rect 39330 8128 39346 8192
rect 39410 8128 39426 8192
rect 39490 8128 39506 8192
rect 39570 8128 39576 8192
rect 39260 8127 39576 8128
rect 32949 7986 33015 7989
rect 36077 7986 36143 7989
rect 32949 7984 36143 7986
rect 32949 7928 32954 7984
rect 33010 7928 36082 7984
rect 36138 7928 36143 7984
rect 32949 7926 36143 7928
rect 32949 7923 33015 7926
rect 36077 7923 36143 7926
rect 44357 7850 44423 7853
rect 44357 7848 45202 7850
rect 44357 7792 44362 7848
rect 44418 7792 45202 7848
rect 44357 7790 45202 7792
rect 44357 7787 44423 7790
rect 45142 7668 45202 7790
rect 11892 7648 12208 7649
rect 11892 7584 11898 7648
rect 11962 7584 11978 7648
rect 12042 7584 12058 7648
rect 12122 7584 12138 7648
rect 12202 7584 12208 7648
rect 11892 7583 12208 7584
rect 22839 7648 23155 7649
rect 22839 7584 22845 7648
rect 22909 7584 22925 7648
rect 22989 7584 23005 7648
rect 23069 7584 23085 7648
rect 23149 7584 23155 7648
rect 22839 7583 23155 7584
rect 33786 7648 34102 7649
rect 33786 7584 33792 7648
rect 33856 7584 33872 7648
rect 33936 7584 33952 7648
rect 34016 7584 34032 7648
rect 34096 7584 34102 7648
rect 33786 7583 34102 7584
rect 44733 7648 45049 7649
rect 44733 7584 44739 7648
rect 44803 7584 44819 7648
rect 44883 7584 44899 7648
rect 44963 7584 44979 7648
rect 45043 7584 45049 7648
rect 44733 7583 45049 7584
rect 45142 7518 46000 7668
rect 45200 7428 46000 7518
rect 6419 7104 6735 7105
rect 6419 7040 6425 7104
rect 6489 7040 6505 7104
rect 6569 7040 6585 7104
rect 6649 7040 6665 7104
rect 6729 7040 6735 7104
rect 6419 7039 6735 7040
rect 17366 7104 17682 7105
rect 17366 7040 17372 7104
rect 17436 7040 17452 7104
rect 17516 7040 17532 7104
rect 17596 7040 17612 7104
rect 17676 7040 17682 7104
rect 17366 7039 17682 7040
rect 28313 7104 28629 7105
rect 28313 7040 28319 7104
rect 28383 7040 28399 7104
rect 28463 7040 28479 7104
rect 28543 7040 28559 7104
rect 28623 7040 28629 7104
rect 28313 7039 28629 7040
rect 39260 7104 39576 7105
rect 39260 7040 39266 7104
rect 39330 7040 39346 7104
rect 39410 7040 39426 7104
rect 39490 7040 39506 7104
rect 39570 7040 39576 7104
rect 39260 7039 39576 7040
rect 0 6898 800 6988
rect 933 6898 999 6901
rect 0 6896 999 6898
rect 0 6840 938 6896
rect 994 6840 999 6896
rect 0 6838 999 6840
rect 0 6748 800 6838
rect 933 6835 999 6838
rect 34421 6898 34487 6901
rect 36905 6898 36971 6901
rect 34421 6896 36971 6898
rect 34421 6840 34426 6896
rect 34482 6840 36910 6896
rect 36966 6840 36971 6896
rect 34421 6838 36971 6840
rect 34421 6835 34487 6838
rect 36905 6835 36971 6838
rect 11892 6560 12208 6561
rect 11892 6496 11898 6560
rect 11962 6496 11978 6560
rect 12042 6496 12058 6560
rect 12122 6496 12138 6560
rect 12202 6496 12208 6560
rect 11892 6495 12208 6496
rect 22839 6560 23155 6561
rect 22839 6496 22845 6560
rect 22909 6496 22925 6560
rect 22989 6496 23005 6560
rect 23069 6496 23085 6560
rect 23149 6496 23155 6560
rect 22839 6495 23155 6496
rect 33786 6560 34102 6561
rect 33786 6496 33792 6560
rect 33856 6496 33872 6560
rect 33936 6496 33952 6560
rect 34016 6496 34032 6560
rect 34096 6496 34102 6560
rect 33786 6495 34102 6496
rect 44733 6560 45049 6561
rect 44733 6496 44739 6560
rect 44803 6496 44819 6560
rect 44883 6496 44899 6560
rect 44963 6496 44979 6560
rect 45043 6496 45049 6560
rect 44733 6495 45049 6496
rect 27521 6218 27587 6221
rect 41965 6218 42031 6221
rect 27521 6216 42031 6218
rect 27521 6160 27526 6216
rect 27582 6160 41970 6216
rect 42026 6160 42031 6216
rect 27521 6158 42031 6160
rect 27521 6155 27587 6158
rect 41965 6155 42031 6158
rect 34513 6082 34579 6085
rect 37089 6082 37155 6085
rect 34513 6080 37155 6082
rect 34513 6024 34518 6080
rect 34574 6024 37094 6080
rect 37150 6024 37155 6080
rect 34513 6022 37155 6024
rect 34513 6019 34579 6022
rect 37089 6019 37155 6022
rect 6419 6016 6735 6017
rect 6419 5952 6425 6016
rect 6489 5952 6505 6016
rect 6569 5952 6585 6016
rect 6649 5952 6665 6016
rect 6729 5952 6735 6016
rect 6419 5951 6735 5952
rect 17366 6016 17682 6017
rect 17366 5952 17372 6016
rect 17436 5952 17452 6016
rect 17516 5952 17532 6016
rect 17596 5952 17612 6016
rect 17676 5952 17682 6016
rect 17366 5951 17682 5952
rect 28313 6016 28629 6017
rect 28313 5952 28319 6016
rect 28383 5952 28399 6016
rect 28463 5952 28479 6016
rect 28543 5952 28559 6016
rect 28623 5952 28629 6016
rect 28313 5951 28629 5952
rect 39260 6016 39576 6017
rect 39260 5952 39266 6016
rect 39330 5952 39346 6016
rect 39410 5952 39426 6016
rect 39490 5952 39506 6016
rect 39570 5952 39576 6016
rect 39260 5951 39576 5952
rect 8385 5810 8451 5813
rect 23933 5810 23999 5813
rect 27521 5810 27587 5813
rect 8385 5808 27587 5810
rect 8385 5752 8390 5808
rect 8446 5752 23938 5808
rect 23994 5752 27526 5808
rect 27582 5752 27587 5808
rect 8385 5750 27587 5752
rect 8385 5747 8451 5750
rect 23933 5747 23999 5750
rect 27521 5747 27587 5750
rect 14457 5674 14523 5677
rect 25865 5674 25931 5677
rect 14457 5672 25931 5674
rect 14457 5616 14462 5672
rect 14518 5616 25870 5672
rect 25926 5616 25931 5672
rect 14457 5614 25931 5616
rect 14457 5611 14523 5614
rect 25865 5611 25931 5614
rect 34881 5674 34947 5677
rect 36905 5674 36971 5677
rect 34881 5672 36971 5674
rect 34881 5616 34886 5672
rect 34942 5616 36910 5672
rect 36966 5616 36971 5672
rect 34881 5614 36971 5616
rect 34881 5611 34947 5614
rect 36905 5611 36971 5614
rect 13353 5538 13419 5541
rect 18505 5538 18571 5541
rect 45200 5538 46000 5628
rect 13353 5536 18571 5538
rect 13353 5480 13358 5536
rect 13414 5480 18510 5536
rect 18566 5480 18571 5536
rect 13353 5478 18571 5480
rect 13353 5475 13419 5478
rect 18505 5475 18571 5478
rect 11892 5472 12208 5473
rect 11892 5408 11898 5472
rect 11962 5408 11978 5472
rect 12042 5408 12058 5472
rect 12122 5408 12138 5472
rect 12202 5408 12208 5472
rect 11892 5407 12208 5408
rect 22839 5472 23155 5473
rect 22839 5408 22845 5472
rect 22909 5408 22925 5472
rect 22989 5408 23005 5472
rect 23069 5408 23085 5472
rect 23149 5408 23155 5472
rect 22839 5407 23155 5408
rect 33786 5472 34102 5473
rect 33786 5408 33792 5472
rect 33856 5408 33872 5472
rect 33936 5408 33952 5472
rect 34016 5408 34032 5472
rect 34096 5408 34102 5472
rect 33786 5407 34102 5408
rect 44733 5472 45049 5473
rect 44733 5408 44739 5472
rect 44803 5408 44819 5472
rect 44883 5408 44899 5472
rect 44963 5408 44979 5472
rect 45043 5408 45049 5472
rect 44733 5407 45049 5408
rect 45142 5388 46000 5538
rect 6177 5266 6243 5269
rect 41413 5266 41479 5269
rect 45142 5266 45202 5388
rect 6177 5264 22110 5266
rect 6177 5208 6182 5264
rect 6238 5208 22110 5264
rect 6177 5206 22110 5208
rect 6177 5203 6243 5206
rect 15837 5130 15903 5133
rect 17953 5130 18019 5133
rect 15837 5128 18019 5130
rect 15837 5072 15842 5128
rect 15898 5072 17958 5128
rect 18014 5072 18019 5128
rect 15837 5070 18019 5072
rect 22050 5130 22110 5206
rect 41413 5264 45202 5266
rect 41413 5208 41418 5264
rect 41474 5208 45202 5264
rect 41413 5206 45202 5208
rect 41413 5203 41479 5206
rect 42793 5130 42859 5133
rect 22050 5128 42859 5130
rect 22050 5072 42798 5128
rect 42854 5072 42859 5128
rect 22050 5070 42859 5072
rect 15837 5067 15903 5070
rect 17953 5067 18019 5070
rect 42793 5067 42859 5070
rect 0 4858 800 4948
rect 6419 4928 6735 4929
rect 6419 4864 6425 4928
rect 6489 4864 6505 4928
rect 6569 4864 6585 4928
rect 6649 4864 6665 4928
rect 6729 4864 6735 4928
rect 6419 4863 6735 4864
rect 17366 4928 17682 4929
rect 17366 4864 17372 4928
rect 17436 4864 17452 4928
rect 17516 4864 17532 4928
rect 17596 4864 17612 4928
rect 17676 4864 17682 4928
rect 17366 4863 17682 4864
rect 28313 4928 28629 4929
rect 28313 4864 28319 4928
rect 28383 4864 28399 4928
rect 28463 4864 28479 4928
rect 28543 4864 28559 4928
rect 28623 4864 28629 4928
rect 28313 4863 28629 4864
rect 39260 4928 39576 4929
rect 39260 4864 39266 4928
rect 39330 4864 39346 4928
rect 39410 4864 39426 4928
rect 39490 4864 39506 4928
rect 39570 4864 39576 4928
rect 39260 4863 39576 4864
rect 933 4858 999 4861
rect 0 4856 999 4858
rect 0 4800 938 4856
rect 994 4800 999 4856
rect 0 4798 999 4800
rect 0 4708 800 4798
rect 933 4795 999 4798
rect 11892 4384 12208 4385
rect 11892 4320 11898 4384
rect 11962 4320 11978 4384
rect 12042 4320 12058 4384
rect 12122 4320 12138 4384
rect 12202 4320 12208 4384
rect 11892 4319 12208 4320
rect 22839 4384 23155 4385
rect 22839 4320 22845 4384
rect 22909 4320 22925 4384
rect 22989 4320 23005 4384
rect 23069 4320 23085 4384
rect 23149 4320 23155 4384
rect 22839 4319 23155 4320
rect 33786 4384 34102 4385
rect 33786 4320 33792 4384
rect 33856 4320 33872 4384
rect 33936 4320 33952 4384
rect 34016 4320 34032 4384
rect 34096 4320 34102 4384
rect 33786 4319 34102 4320
rect 44733 4384 45049 4385
rect 44733 4320 44739 4384
rect 44803 4320 44819 4384
rect 44883 4320 44899 4384
rect 44963 4320 44979 4384
rect 45043 4320 45049 4384
rect 44733 4319 45049 4320
rect 44633 4178 44699 4181
rect 45200 4178 46000 4268
rect 44633 4176 46000 4178
rect 44633 4120 44638 4176
rect 44694 4120 46000 4176
rect 44633 4118 46000 4120
rect 44633 4115 44699 4118
rect 45200 4028 46000 4118
rect 6419 3840 6735 3841
rect 6419 3776 6425 3840
rect 6489 3776 6505 3840
rect 6569 3776 6585 3840
rect 6649 3776 6665 3840
rect 6729 3776 6735 3840
rect 6419 3775 6735 3776
rect 17366 3840 17682 3841
rect 17366 3776 17372 3840
rect 17436 3776 17452 3840
rect 17516 3776 17532 3840
rect 17596 3776 17612 3840
rect 17676 3776 17682 3840
rect 17366 3775 17682 3776
rect 28313 3840 28629 3841
rect 28313 3776 28319 3840
rect 28383 3776 28399 3840
rect 28463 3776 28479 3840
rect 28543 3776 28559 3840
rect 28623 3776 28629 3840
rect 28313 3775 28629 3776
rect 39260 3840 39576 3841
rect 39260 3776 39266 3840
rect 39330 3776 39346 3840
rect 39410 3776 39426 3840
rect 39490 3776 39506 3840
rect 39570 3776 39576 3840
rect 39260 3775 39576 3776
rect 0 3498 800 3588
rect 933 3498 999 3501
rect 0 3496 999 3498
rect 0 3440 938 3496
rect 994 3440 999 3496
rect 0 3438 999 3440
rect 0 3348 800 3438
rect 933 3435 999 3438
rect 11892 3296 12208 3297
rect 11892 3232 11898 3296
rect 11962 3232 11978 3296
rect 12042 3232 12058 3296
rect 12122 3232 12138 3296
rect 12202 3232 12208 3296
rect 11892 3231 12208 3232
rect 22839 3296 23155 3297
rect 22839 3232 22845 3296
rect 22909 3232 22925 3296
rect 22989 3232 23005 3296
rect 23069 3232 23085 3296
rect 23149 3232 23155 3296
rect 22839 3231 23155 3232
rect 33786 3296 34102 3297
rect 33786 3232 33792 3296
rect 33856 3232 33872 3296
rect 33936 3232 33952 3296
rect 34016 3232 34032 3296
rect 34096 3232 34102 3296
rect 33786 3231 34102 3232
rect 44733 3296 45049 3297
rect 44733 3232 44739 3296
rect 44803 3232 44819 3296
rect 44883 3232 44899 3296
rect 44963 3232 44979 3296
rect 45043 3232 45049 3296
rect 44733 3231 45049 3232
rect 6419 2752 6735 2753
rect 6419 2688 6425 2752
rect 6489 2688 6505 2752
rect 6569 2688 6585 2752
rect 6649 2688 6665 2752
rect 6729 2688 6735 2752
rect 6419 2687 6735 2688
rect 17366 2752 17682 2753
rect 17366 2688 17372 2752
rect 17436 2688 17452 2752
rect 17516 2688 17532 2752
rect 17596 2688 17612 2752
rect 17676 2688 17682 2752
rect 17366 2687 17682 2688
rect 28313 2752 28629 2753
rect 28313 2688 28319 2752
rect 28383 2688 28399 2752
rect 28463 2688 28479 2752
rect 28543 2688 28559 2752
rect 28623 2688 28629 2752
rect 28313 2687 28629 2688
rect 39260 2752 39576 2753
rect 39260 2688 39266 2752
rect 39330 2688 39346 2752
rect 39410 2688 39426 2752
rect 39490 2688 39506 2752
rect 39570 2688 39576 2752
rect 39260 2687 39576 2688
rect 41413 2410 41479 2413
rect 41413 2408 45202 2410
rect 41413 2352 41418 2408
rect 41474 2352 45202 2408
rect 41413 2350 45202 2352
rect 41413 2347 41479 2350
rect 45142 2228 45202 2350
rect 11892 2208 12208 2209
rect 11892 2144 11898 2208
rect 11962 2144 11978 2208
rect 12042 2144 12058 2208
rect 12122 2144 12138 2208
rect 12202 2144 12208 2208
rect 11892 2143 12208 2144
rect 22839 2208 23155 2209
rect 22839 2144 22845 2208
rect 22909 2144 22925 2208
rect 22989 2144 23005 2208
rect 23069 2144 23085 2208
rect 23149 2144 23155 2208
rect 22839 2143 23155 2144
rect 33786 2208 34102 2209
rect 33786 2144 33792 2208
rect 33856 2144 33872 2208
rect 33936 2144 33952 2208
rect 34016 2144 34032 2208
rect 34096 2144 34102 2208
rect 33786 2143 34102 2144
rect 44733 2208 45049 2209
rect 44733 2144 44739 2208
rect 44803 2144 44819 2208
rect 44883 2144 44899 2208
rect 44963 2144 44979 2208
rect 45043 2144 45049 2208
rect 44733 2143 45049 2144
rect 45142 2078 46000 2228
rect 45200 1988 46000 2078
rect 0 1458 800 1548
rect 933 1458 999 1461
rect 0 1456 999 1458
rect 0 1400 938 1456
rect 994 1400 999 1456
rect 0 1398 999 1400
rect 0 1308 800 1398
rect 933 1395 999 1398
rect 44633 778 44699 781
rect 45200 778 46000 868
rect 44633 776 46000 778
rect 44633 720 44638 776
rect 44694 720 46000 776
rect 44633 718 46000 720
rect 44633 715 44699 718
rect 45200 628 46000 718
<< via3 >>
rect 11898 17436 11962 17440
rect 11898 17380 11902 17436
rect 11902 17380 11958 17436
rect 11958 17380 11962 17436
rect 11898 17376 11962 17380
rect 11978 17436 12042 17440
rect 11978 17380 11982 17436
rect 11982 17380 12038 17436
rect 12038 17380 12042 17436
rect 11978 17376 12042 17380
rect 12058 17436 12122 17440
rect 12058 17380 12062 17436
rect 12062 17380 12118 17436
rect 12118 17380 12122 17436
rect 12058 17376 12122 17380
rect 12138 17436 12202 17440
rect 12138 17380 12142 17436
rect 12142 17380 12198 17436
rect 12198 17380 12202 17436
rect 12138 17376 12202 17380
rect 22845 17436 22909 17440
rect 22845 17380 22849 17436
rect 22849 17380 22905 17436
rect 22905 17380 22909 17436
rect 22845 17376 22909 17380
rect 22925 17436 22989 17440
rect 22925 17380 22929 17436
rect 22929 17380 22985 17436
rect 22985 17380 22989 17436
rect 22925 17376 22989 17380
rect 23005 17436 23069 17440
rect 23005 17380 23009 17436
rect 23009 17380 23065 17436
rect 23065 17380 23069 17436
rect 23005 17376 23069 17380
rect 23085 17436 23149 17440
rect 23085 17380 23089 17436
rect 23089 17380 23145 17436
rect 23145 17380 23149 17436
rect 23085 17376 23149 17380
rect 33792 17436 33856 17440
rect 33792 17380 33796 17436
rect 33796 17380 33852 17436
rect 33852 17380 33856 17436
rect 33792 17376 33856 17380
rect 33872 17436 33936 17440
rect 33872 17380 33876 17436
rect 33876 17380 33932 17436
rect 33932 17380 33936 17436
rect 33872 17376 33936 17380
rect 33952 17436 34016 17440
rect 33952 17380 33956 17436
rect 33956 17380 34012 17436
rect 34012 17380 34016 17436
rect 33952 17376 34016 17380
rect 34032 17436 34096 17440
rect 34032 17380 34036 17436
rect 34036 17380 34092 17436
rect 34092 17380 34096 17436
rect 34032 17376 34096 17380
rect 44739 17436 44803 17440
rect 44739 17380 44743 17436
rect 44743 17380 44799 17436
rect 44799 17380 44803 17436
rect 44739 17376 44803 17380
rect 44819 17436 44883 17440
rect 44819 17380 44823 17436
rect 44823 17380 44879 17436
rect 44879 17380 44883 17436
rect 44819 17376 44883 17380
rect 44899 17436 44963 17440
rect 44899 17380 44903 17436
rect 44903 17380 44959 17436
rect 44959 17380 44963 17436
rect 44899 17376 44963 17380
rect 44979 17436 45043 17440
rect 44979 17380 44983 17436
rect 44983 17380 45039 17436
rect 45039 17380 45043 17436
rect 44979 17376 45043 17380
rect 6425 16892 6489 16896
rect 6425 16836 6429 16892
rect 6429 16836 6485 16892
rect 6485 16836 6489 16892
rect 6425 16832 6489 16836
rect 6505 16892 6569 16896
rect 6505 16836 6509 16892
rect 6509 16836 6565 16892
rect 6565 16836 6569 16892
rect 6505 16832 6569 16836
rect 6585 16892 6649 16896
rect 6585 16836 6589 16892
rect 6589 16836 6645 16892
rect 6645 16836 6649 16892
rect 6585 16832 6649 16836
rect 6665 16892 6729 16896
rect 6665 16836 6669 16892
rect 6669 16836 6725 16892
rect 6725 16836 6729 16892
rect 6665 16832 6729 16836
rect 17372 16892 17436 16896
rect 17372 16836 17376 16892
rect 17376 16836 17432 16892
rect 17432 16836 17436 16892
rect 17372 16832 17436 16836
rect 17452 16892 17516 16896
rect 17452 16836 17456 16892
rect 17456 16836 17512 16892
rect 17512 16836 17516 16892
rect 17452 16832 17516 16836
rect 17532 16892 17596 16896
rect 17532 16836 17536 16892
rect 17536 16836 17592 16892
rect 17592 16836 17596 16892
rect 17532 16832 17596 16836
rect 17612 16892 17676 16896
rect 17612 16836 17616 16892
rect 17616 16836 17672 16892
rect 17672 16836 17676 16892
rect 17612 16832 17676 16836
rect 28319 16892 28383 16896
rect 28319 16836 28323 16892
rect 28323 16836 28379 16892
rect 28379 16836 28383 16892
rect 28319 16832 28383 16836
rect 28399 16892 28463 16896
rect 28399 16836 28403 16892
rect 28403 16836 28459 16892
rect 28459 16836 28463 16892
rect 28399 16832 28463 16836
rect 28479 16892 28543 16896
rect 28479 16836 28483 16892
rect 28483 16836 28539 16892
rect 28539 16836 28543 16892
rect 28479 16832 28543 16836
rect 28559 16892 28623 16896
rect 28559 16836 28563 16892
rect 28563 16836 28619 16892
rect 28619 16836 28623 16892
rect 28559 16832 28623 16836
rect 39266 16892 39330 16896
rect 39266 16836 39270 16892
rect 39270 16836 39326 16892
rect 39326 16836 39330 16892
rect 39266 16832 39330 16836
rect 39346 16892 39410 16896
rect 39346 16836 39350 16892
rect 39350 16836 39406 16892
rect 39406 16836 39410 16892
rect 39346 16832 39410 16836
rect 39426 16892 39490 16896
rect 39426 16836 39430 16892
rect 39430 16836 39486 16892
rect 39486 16836 39490 16892
rect 39426 16832 39490 16836
rect 39506 16892 39570 16896
rect 39506 16836 39510 16892
rect 39510 16836 39566 16892
rect 39566 16836 39570 16892
rect 39506 16832 39570 16836
rect 11898 16348 11962 16352
rect 11898 16292 11902 16348
rect 11902 16292 11958 16348
rect 11958 16292 11962 16348
rect 11898 16288 11962 16292
rect 11978 16348 12042 16352
rect 11978 16292 11982 16348
rect 11982 16292 12038 16348
rect 12038 16292 12042 16348
rect 11978 16288 12042 16292
rect 12058 16348 12122 16352
rect 12058 16292 12062 16348
rect 12062 16292 12118 16348
rect 12118 16292 12122 16348
rect 12058 16288 12122 16292
rect 12138 16348 12202 16352
rect 12138 16292 12142 16348
rect 12142 16292 12198 16348
rect 12198 16292 12202 16348
rect 12138 16288 12202 16292
rect 22845 16348 22909 16352
rect 22845 16292 22849 16348
rect 22849 16292 22905 16348
rect 22905 16292 22909 16348
rect 22845 16288 22909 16292
rect 22925 16348 22989 16352
rect 22925 16292 22929 16348
rect 22929 16292 22985 16348
rect 22985 16292 22989 16348
rect 22925 16288 22989 16292
rect 23005 16348 23069 16352
rect 23005 16292 23009 16348
rect 23009 16292 23065 16348
rect 23065 16292 23069 16348
rect 23005 16288 23069 16292
rect 23085 16348 23149 16352
rect 23085 16292 23089 16348
rect 23089 16292 23145 16348
rect 23145 16292 23149 16348
rect 23085 16288 23149 16292
rect 33792 16348 33856 16352
rect 33792 16292 33796 16348
rect 33796 16292 33852 16348
rect 33852 16292 33856 16348
rect 33792 16288 33856 16292
rect 33872 16348 33936 16352
rect 33872 16292 33876 16348
rect 33876 16292 33932 16348
rect 33932 16292 33936 16348
rect 33872 16288 33936 16292
rect 33952 16348 34016 16352
rect 33952 16292 33956 16348
rect 33956 16292 34012 16348
rect 34012 16292 34016 16348
rect 33952 16288 34016 16292
rect 34032 16348 34096 16352
rect 34032 16292 34036 16348
rect 34036 16292 34092 16348
rect 34092 16292 34096 16348
rect 34032 16288 34096 16292
rect 44739 16348 44803 16352
rect 44739 16292 44743 16348
rect 44743 16292 44799 16348
rect 44799 16292 44803 16348
rect 44739 16288 44803 16292
rect 44819 16348 44883 16352
rect 44819 16292 44823 16348
rect 44823 16292 44879 16348
rect 44879 16292 44883 16348
rect 44819 16288 44883 16292
rect 44899 16348 44963 16352
rect 44899 16292 44903 16348
rect 44903 16292 44959 16348
rect 44959 16292 44963 16348
rect 44899 16288 44963 16292
rect 44979 16348 45043 16352
rect 44979 16292 44983 16348
rect 44983 16292 45039 16348
rect 45039 16292 45043 16348
rect 44979 16288 45043 16292
rect 6425 15804 6489 15808
rect 6425 15748 6429 15804
rect 6429 15748 6485 15804
rect 6485 15748 6489 15804
rect 6425 15744 6489 15748
rect 6505 15804 6569 15808
rect 6505 15748 6509 15804
rect 6509 15748 6565 15804
rect 6565 15748 6569 15804
rect 6505 15744 6569 15748
rect 6585 15804 6649 15808
rect 6585 15748 6589 15804
rect 6589 15748 6645 15804
rect 6645 15748 6649 15804
rect 6585 15744 6649 15748
rect 6665 15804 6729 15808
rect 6665 15748 6669 15804
rect 6669 15748 6725 15804
rect 6725 15748 6729 15804
rect 6665 15744 6729 15748
rect 17372 15804 17436 15808
rect 17372 15748 17376 15804
rect 17376 15748 17432 15804
rect 17432 15748 17436 15804
rect 17372 15744 17436 15748
rect 17452 15804 17516 15808
rect 17452 15748 17456 15804
rect 17456 15748 17512 15804
rect 17512 15748 17516 15804
rect 17452 15744 17516 15748
rect 17532 15804 17596 15808
rect 17532 15748 17536 15804
rect 17536 15748 17592 15804
rect 17592 15748 17596 15804
rect 17532 15744 17596 15748
rect 17612 15804 17676 15808
rect 17612 15748 17616 15804
rect 17616 15748 17672 15804
rect 17672 15748 17676 15804
rect 17612 15744 17676 15748
rect 28319 15804 28383 15808
rect 28319 15748 28323 15804
rect 28323 15748 28379 15804
rect 28379 15748 28383 15804
rect 28319 15744 28383 15748
rect 28399 15804 28463 15808
rect 28399 15748 28403 15804
rect 28403 15748 28459 15804
rect 28459 15748 28463 15804
rect 28399 15744 28463 15748
rect 28479 15804 28543 15808
rect 28479 15748 28483 15804
rect 28483 15748 28539 15804
rect 28539 15748 28543 15804
rect 28479 15744 28543 15748
rect 28559 15804 28623 15808
rect 28559 15748 28563 15804
rect 28563 15748 28619 15804
rect 28619 15748 28623 15804
rect 28559 15744 28623 15748
rect 39266 15804 39330 15808
rect 39266 15748 39270 15804
rect 39270 15748 39326 15804
rect 39326 15748 39330 15804
rect 39266 15744 39330 15748
rect 39346 15804 39410 15808
rect 39346 15748 39350 15804
rect 39350 15748 39406 15804
rect 39406 15748 39410 15804
rect 39346 15744 39410 15748
rect 39426 15804 39490 15808
rect 39426 15748 39430 15804
rect 39430 15748 39486 15804
rect 39486 15748 39490 15804
rect 39426 15744 39490 15748
rect 39506 15804 39570 15808
rect 39506 15748 39510 15804
rect 39510 15748 39566 15804
rect 39566 15748 39570 15804
rect 39506 15744 39570 15748
rect 11898 15260 11962 15264
rect 11898 15204 11902 15260
rect 11902 15204 11958 15260
rect 11958 15204 11962 15260
rect 11898 15200 11962 15204
rect 11978 15260 12042 15264
rect 11978 15204 11982 15260
rect 11982 15204 12038 15260
rect 12038 15204 12042 15260
rect 11978 15200 12042 15204
rect 12058 15260 12122 15264
rect 12058 15204 12062 15260
rect 12062 15204 12118 15260
rect 12118 15204 12122 15260
rect 12058 15200 12122 15204
rect 12138 15260 12202 15264
rect 12138 15204 12142 15260
rect 12142 15204 12198 15260
rect 12198 15204 12202 15260
rect 12138 15200 12202 15204
rect 22845 15260 22909 15264
rect 22845 15204 22849 15260
rect 22849 15204 22905 15260
rect 22905 15204 22909 15260
rect 22845 15200 22909 15204
rect 22925 15260 22989 15264
rect 22925 15204 22929 15260
rect 22929 15204 22985 15260
rect 22985 15204 22989 15260
rect 22925 15200 22989 15204
rect 23005 15260 23069 15264
rect 23005 15204 23009 15260
rect 23009 15204 23065 15260
rect 23065 15204 23069 15260
rect 23005 15200 23069 15204
rect 23085 15260 23149 15264
rect 23085 15204 23089 15260
rect 23089 15204 23145 15260
rect 23145 15204 23149 15260
rect 23085 15200 23149 15204
rect 33792 15260 33856 15264
rect 33792 15204 33796 15260
rect 33796 15204 33852 15260
rect 33852 15204 33856 15260
rect 33792 15200 33856 15204
rect 33872 15260 33936 15264
rect 33872 15204 33876 15260
rect 33876 15204 33932 15260
rect 33932 15204 33936 15260
rect 33872 15200 33936 15204
rect 33952 15260 34016 15264
rect 33952 15204 33956 15260
rect 33956 15204 34012 15260
rect 34012 15204 34016 15260
rect 33952 15200 34016 15204
rect 34032 15260 34096 15264
rect 34032 15204 34036 15260
rect 34036 15204 34092 15260
rect 34092 15204 34096 15260
rect 34032 15200 34096 15204
rect 44739 15260 44803 15264
rect 44739 15204 44743 15260
rect 44743 15204 44799 15260
rect 44799 15204 44803 15260
rect 44739 15200 44803 15204
rect 44819 15260 44883 15264
rect 44819 15204 44823 15260
rect 44823 15204 44879 15260
rect 44879 15204 44883 15260
rect 44819 15200 44883 15204
rect 44899 15260 44963 15264
rect 44899 15204 44903 15260
rect 44903 15204 44959 15260
rect 44959 15204 44963 15260
rect 44899 15200 44963 15204
rect 44979 15260 45043 15264
rect 44979 15204 44983 15260
rect 44983 15204 45039 15260
rect 45039 15204 45043 15260
rect 44979 15200 45043 15204
rect 6425 14716 6489 14720
rect 6425 14660 6429 14716
rect 6429 14660 6485 14716
rect 6485 14660 6489 14716
rect 6425 14656 6489 14660
rect 6505 14716 6569 14720
rect 6505 14660 6509 14716
rect 6509 14660 6565 14716
rect 6565 14660 6569 14716
rect 6505 14656 6569 14660
rect 6585 14716 6649 14720
rect 6585 14660 6589 14716
rect 6589 14660 6645 14716
rect 6645 14660 6649 14716
rect 6585 14656 6649 14660
rect 6665 14716 6729 14720
rect 6665 14660 6669 14716
rect 6669 14660 6725 14716
rect 6725 14660 6729 14716
rect 6665 14656 6729 14660
rect 17372 14716 17436 14720
rect 17372 14660 17376 14716
rect 17376 14660 17432 14716
rect 17432 14660 17436 14716
rect 17372 14656 17436 14660
rect 17452 14716 17516 14720
rect 17452 14660 17456 14716
rect 17456 14660 17512 14716
rect 17512 14660 17516 14716
rect 17452 14656 17516 14660
rect 17532 14716 17596 14720
rect 17532 14660 17536 14716
rect 17536 14660 17592 14716
rect 17592 14660 17596 14716
rect 17532 14656 17596 14660
rect 17612 14716 17676 14720
rect 17612 14660 17616 14716
rect 17616 14660 17672 14716
rect 17672 14660 17676 14716
rect 17612 14656 17676 14660
rect 28319 14716 28383 14720
rect 28319 14660 28323 14716
rect 28323 14660 28379 14716
rect 28379 14660 28383 14716
rect 28319 14656 28383 14660
rect 28399 14716 28463 14720
rect 28399 14660 28403 14716
rect 28403 14660 28459 14716
rect 28459 14660 28463 14716
rect 28399 14656 28463 14660
rect 28479 14716 28543 14720
rect 28479 14660 28483 14716
rect 28483 14660 28539 14716
rect 28539 14660 28543 14716
rect 28479 14656 28543 14660
rect 28559 14716 28623 14720
rect 28559 14660 28563 14716
rect 28563 14660 28619 14716
rect 28619 14660 28623 14716
rect 28559 14656 28623 14660
rect 39266 14716 39330 14720
rect 39266 14660 39270 14716
rect 39270 14660 39326 14716
rect 39326 14660 39330 14716
rect 39266 14656 39330 14660
rect 39346 14716 39410 14720
rect 39346 14660 39350 14716
rect 39350 14660 39406 14716
rect 39406 14660 39410 14716
rect 39346 14656 39410 14660
rect 39426 14716 39490 14720
rect 39426 14660 39430 14716
rect 39430 14660 39486 14716
rect 39486 14660 39490 14716
rect 39426 14656 39490 14660
rect 39506 14716 39570 14720
rect 39506 14660 39510 14716
rect 39510 14660 39566 14716
rect 39566 14660 39570 14716
rect 39506 14656 39570 14660
rect 11898 14172 11962 14176
rect 11898 14116 11902 14172
rect 11902 14116 11958 14172
rect 11958 14116 11962 14172
rect 11898 14112 11962 14116
rect 11978 14172 12042 14176
rect 11978 14116 11982 14172
rect 11982 14116 12038 14172
rect 12038 14116 12042 14172
rect 11978 14112 12042 14116
rect 12058 14172 12122 14176
rect 12058 14116 12062 14172
rect 12062 14116 12118 14172
rect 12118 14116 12122 14172
rect 12058 14112 12122 14116
rect 12138 14172 12202 14176
rect 12138 14116 12142 14172
rect 12142 14116 12198 14172
rect 12198 14116 12202 14172
rect 12138 14112 12202 14116
rect 22845 14172 22909 14176
rect 22845 14116 22849 14172
rect 22849 14116 22905 14172
rect 22905 14116 22909 14172
rect 22845 14112 22909 14116
rect 22925 14172 22989 14176
rect 22925 14116 22929 14172
rect 22929 14116 22985 14172
rect 22985 14116 22989 14172
rect 22925 14112 22989 14116
rect 23005 14172 23069 14176
rect 23005 14116 23009 14172
rect 23009 14116 23065 14172
rect 23065 14116 23069 14172
rect 23005 14112 23069 14116
rect 23085 14172 23149 14176
rect 23085 14116 23089 14172
rect 23089 14116 23145 14172
rect 23145 14116 23149 14172
rect 23085 14112 23149 14116
rect 33792 14172 33856 14176
rect 33792 14116 33796 14172
rect 33796 14116 33852 14172
rect 33852 14116 33856 14172
rect 33792 14112 33856 14116
rect 33872 14172 33936 14176
rect 33872 14116 33876 14172
rect 33876 14116 33932 14172
rect 33932 14116 33936 14172
rect 33872 14112 33936 14116
rect 33952 14172 34016 14176
rect 33952 14116 33956 14172
rect 33956 14116 34012 14172
rect 34012 14116 34016 14172
rect 33952 14112 34016 14116
rect 34032 14172 34096 14176
rect 34032 14116 34036 14172
rect 34036 14116 34092 14172
rect 34092 14116 34096 14172
rect 34032 14112 34096 14116
rect 44739 14172 44803 14176
rect 44739 14116 44743 14172
rect 44743 14116 44799 14172
rect 44799 14116 44803 14172
rect 44739 14112 44803 14116
rect 44819 14172 44883 14176
rect 44819 14116 44823 14172
rect 44823 14116 44879 14172
rect 44879 14116 44883 14172
rect 44819 14112 44883 14116
rect 44899 14172 44963 14176
rect 44899 14116 44903 14172
rect 44903 14116 44959 14172
rect 44959 14116 44963 14172
rect 44899 14112 44963 14116
rect 44979 14172 45043 14176
rect 44979 14116 44983 14172
rect 44983 14116 45039 14172
rect 45039 14116 45043 14172
rect 44979 14112 45043 14116
rect 6425 13628 6489 13632
rect 6425 13572 6429 13628
rect 6429 13572 6485 13628
rect 6485 13572 6489 13628
rect 6425 13568 6489 13572
rect 6505 13628 6569 13632
rect 6505 13572 6509 13628
rect 6509 13572 6565 13628
rect 6565 13572 6569 13628
rect 6505 13568 6569 13572
rect 6585 13628 6649 13632
rect 6585 13572 6589 13628
rect 6589 13572 6645 13628
rect 6645 13572 6649 13628
rect 6585 13568 6649 13572
rect 6665 13628 6729 13632
rect 6665 13572 6669 13628
rect 6669 13572 6725 13628
rect 6725 13572 6729 13628
rect 6665 13568 6729 13572
rect 17372 13628 17436 13632
rect 17372 13572 17376 13628
rect 17376 13572 17432 13628
rect 17432 13572 17436 13628
rect 17372 13568 17436 13572
rect 17452 13628 17516 13632
rect 17452 13572 17456 13628
rect 17456 13572 17512 13628
rect 17512 13572 17516 13628
rect 17452 13568 17516 13572
rect 17532 13628 17596 13632
rect 17532 13572 17536 13628
rect 17536 13572 17592 13628
rect 17592 13572 17596 13628
rect 17532 13568 17596 13572
rect 17612 13628 17676 13632
rect 17612 13572 17616 13628
rect 17616 13572 17672 13628
rect 17672 13572 17676 13628
rect 17612 13568 17676 13572
rect 28319 13628 28383 13632
rect 28319 13572 28323 13628
rect 28323 13572 28379 13628
rect 28379 13572 28383 13628
rect 28319 13568 28383 13572
rect 28399 13628 28463 13632
rect 28399 13572 28403 13628
rect 28403 13572 28459 13628
rect 28459 13572 28463 13628
rect 28399 13568 28463 13572
rect 28479 13628 28543 13632
rect 28479 13572 28483 13628
rect 28483 13572 28539 13628
rect 28539 13572 28543 13628
rect 28479 13568 28543 13572
rect 28559 13628 28623 13632
rect 28559 13572 28563 13628
rect 28563 13572 28619 13628
rect 28619 13572 28623 13628
rect 28559 13568 28623 13572
rect 39266 13628 39330 13632
rect 39266 13572 39270 13628
rect 39270 13572 39326 13628
rect 39326 13572 39330 13628
rect 39266 13568 39330 13572
rect 39346 13628 39410 13632
rect 39346 13572 39350 13628
rect 39350 13572 39406 13628
rect 39406 13572 39410 13628
rect 39346 13568 39410 13572
rect 39426 13628 39490 13632
rect 39426 13572 39430 13628
rect 39430 13572 39486 13628
rect 39486 13572 39490 13628
rect 39426 13568 39490 13572
rect 39506 13628 39570 13632
rect 39506 13572 39510 13628
rect 39510 13572 39566 13628
rect 39566 13572 39570 13628
rect 39506 13568 39570 13572
rect 11898 13084 11962 13088
rect 11898 13028 11902 13084
rect 11902 13028 11958 13084
rect 11958 13028 11962 13084
rect 11898 13024 11962 13028
rect 11978 13084 12042 13088
rect 11978 13028 11982 13084
rect 11982 13028 12038 13084
rect 12038 13028 12042 13084
rect 11978 13024 12042 13028
rect 12058 13084 12122 13088
rect 12058 13028 12062 13084
rect 12062 13028 12118 13084
rect 12118 13028 12122 13084
rect 12058 13024 12122 13028
rect 12138 13084 12202 13088
rect 12138 13028 12142 13084
rect 12142 13028 12198 13084
rect 12198 13028 12202 13084
rect 12138 13024 12202 13028
rect 22845 13084 22909 13088
rect 22845 13028 22849 13084
rect 22849 13028 22905 13084
rect 22905 13028 22909 13084
rect 22845 13024 22909 13028
rect 22925 13084 22989 13088
rect 22925 13028 22929 13084
rect 22929 13028 22985 13084
rect 22985 13028 22989 13084
rect 22925 13024 22989 13028
rect 23005 13084 23069 13088
rect 23005 13028 23009 13084
rect 23009 13028 23065 13084
rect 23065 13028 23069 13084
rect 23005 13024 23069 13028
rect 23085 13084 23149 13088
rect 23085 13028 23089 13084
rect 23089 13028 23145 13084
rect 23145 13028 23149 13084
rect 23085 13024 23149 13028
rect 33792 13084 33856 13088
rect 33792 13028 33796 13084
rect 33796 13028 33852 13084
rect 33852 13028 33856 13084
rect 33792 13024 33856 13028
rect 33872 13084 33936 13088
rect 33872 13028 33876 13084
rect 33876 13028 33932 13084
rect 33932 13028 33936 13084
rect 33872 13024 33936 13028
rect 33952 13084 34016 13088
rect 33952 13028 33956 13084
rect 33956 13028 34012 13084
rect 34012 13028 34016 13084
rect 33952 13024 34016 13028
rect 34032 13084 34096 13088
rect 34032 13028 34036 13084
rect 34036 13028 34092 13084
rect 34092 13028 34096 13084
rect 34032 13024 34096 13028
rect 44739 13084 44803 13088
rect 44739 13028 44743 13084
rect 44743 13028 44799 13084
rect 44799 13028 44803 13084
rect 44739 13024 44803 13028
rect 44819 13084 44883 13088
rect 44819 13028 44823 13084
rect 44823 13028 44879 13084
rect 44879 13028 44883 13084
rect 44819 13024 44883 13028
rect 44899 13084 44963 13088
rect 44899 13028 44903 13084
rect 44903 13028 44959 13084
rect 44959 13028 44963 13084
rect 44899 13024 44963 13028
rect 44979 13084 45043 13088
rect 44979 13028 44983 13084
rect 44983 13028 45039 13084
rect 45039 13028 45043 13084
rect 44979 13024 45043 13028
rect 6425 12540 6489 12544
rect 6425 12484 6429 12540
rect 6429 12484 6485 12540
rect 6485 12484 6489 12540
rect 6425 12480 6489 12484
rect 6505 12540 6569 12544
rect 6505 12484 6509 12540
rect 6509 12484 6565 12540
rect 6565 12484 6569 12540
rect 6505 12480 6569 12484
rect 6585 12540 6649 12544
rect 6585 12484 6589 12540
rect 6589 12484 6645 12540
rect 6645 12484 6649 12540
rect 6585 12480 6649 12484
rect 6665 12540 6729 12544
rect 6665 12484 6669 12540
rect 6669 12484 6725 12540
rect 6725 12484 6729 12540
rect 6665 12480 6729 12484
rect 17372 12540 17436 12544
rect 17372 12484 17376 12540
rect 17376 12484 17432 12540
rect 17432 12484 17436 12540
rect 17372 12480 17436 12484
rect 17452 12540 17516 12544
rect 17452 12484 17456 12540
rect 17456 12484 17512 12540
rect 17512 12484 17516 12540
rect 17452 12480 17516 12484
rect 17532 12540 17596 12544
rect 17532 12484 17536 12540
rect 17536 12484 17592 12540
rect 17592 12484 17596 12540
rect 17532 12480 17596 12484
rect 17612 12540 17676 12544
rect 17612 12484 17616 12540
rect 17616 12484 17672 12540
rect 17672 12484 17676 12540
rect 17612 12480 17676 12484
rect 28319 12540 28383 12544
rect 28319 12484 28323 12540
rect 28323 12484 28379 12540
rect 28379 12484 28383 12540
rect 28319 12480 28383 12484
rect 28399 12540 28463 12544
rect 28399 12484 28403 12540
rect 28403 12484 28459 12540
rect 28459 12484 28463 12540
rect 28399 12480 28463 12484
rect 28479 12540 28543 12544
rect 28479 12484 28483 12540
rect 28483 12484 28539 12540
rect 28539 12484 28543 12540
rect 28479 12480 28543 12484
rect 28559 12540 28623 12544
rect 28559 12484 28563 12540
rect 28563 12484 28619 12540
rect 28619 12484 28623 12540
rect 28559 12480 28623 12484
rect 39266 12540 39330 12544
rect 39266 12484 39270 12540
rect 39270 12484 39326 12540
rect 39326 12484 39330 12540
rect 39266 12480 39330 12484
rect 39346 12540 39410 12544
rect 39346 12484 39350 12540
rect 39350 12484 39406 12540
rect 39406 12484 39410 12540
rect 39346 12480 39410 12484
rect 39426 12540 39490 12544
rect 39426 12484 39430 12540
rect 39430 12484 39486 12540
rect 39486 12484 39490 12540
rect 39426 12480 39490 12484
rect 39506 12540 39570 12544
rect 39506 12484 39510 12540
rect 39510 12484 39566 12540
rect 39566 12484 39570 12540
rect 39506 12480 39570 12484
rect 11898 11996 11962 12000
rect 11898 11940 11902 11996
rect 11902 11940 11958 11996
rect 11958 11940 11962 11996
rect 11898 11936 11962 11940
rect 11978 11996 12042 12000
rect 11978 11940 11982 11996
rect 11982 11940 12038 11996
rect 12038 11940 12042 11996
rect 11978 11936 12042 11940
rect 12058 11996 12122 12000
rect 12058 11940 12062 11996
rect 12062 11940 12118 11996
rect 12118 11940 12122 11996
rect 12058 11936 12122 11940
rect 12138 11996 12202 12000
rect 12138 11940 12142 11996
rect 12142 11940 12198 11996
rect 12198 11940 12202 11996
rect 12138 11936 12202 11940
rect 22845 11996 22909 12000
rect 22845 11940 22849 11996
rect 22849 11940 22905 11996
rect 22905 11940 22909 11996
rect 22845 11936 22909 11940
rect 22925 11996 22989 12000
rect 22925 11940 22929 11996
rect 22929 11940 22985 11996
rect 22985 11940 22989 11996
rect 22925 11936 22989 11940
rect 23005 11996 23069 12000
rect 23005 11940 23009 11996
rect 23009 11940 23065 11996
rect 23065 11940 23069 11996
rect 23005 11936 23069 11940
rect 23085 11996 23149 12000
rect 23085 11940 23089 11996
rect 23089 11940 23145 11996
rect 23145 11940 23149 11996
rect 23085 11936 23149 11940
rect 33792 11996 33856 12000
rect 33792 11940 33796 11996
rect 33796 11940 33852 11996
rect 33852 11940 33856 11996
rect 33792 11936 33856 11940
rect 33872 11996 33936 12000
rect 33872 11940 33876 11996
rect 33876 11940 33932 11996
rect 33932 11940 33936 11996
rect 33872 11936 33936 11940
rect 33952 11996 34016 12000
rect 33952 11940 33956 11996
rect 33956 11940 34012 11996
rect 34012 11940 34016 11996
rect 33952 11936 34016 11940
rect 34032 11996 34096 12000
rect 34032 11940 34036 11996
rect 34036 11940 34092 11996
rect 34092 11940 34096 11996
rect 34032 11936 34096 11940
rect 44739 11996 44803 12000
rect 44739 11940 44743 11996
rect 44743 11940 44799 11996
rect 44799 11940 44803 11996
rect 44739 11936 44803 11940
rect 44819 11996 44883 12000
rect 44819 11940 44823 11996
rect 44823 11940 44879 11996
rect 44879 11940 44883 11996
rect 44819 11936 44883 11940
rect 44899 11996 44963 12000
rect 44899 11940 44903 11996
rect 44903 11940 44959 11996
rect 44959 11940 44963 11996
rect 44899 11936 44963 11940
rect 44979 11996 45043 12000
rect 44979 11940 44983 11996
rect 44983 11940 45039 11996
rect 45039 11940 45043 11996
rect 44979 11936 45043 11940
rect 6425 11452 6489 11456
rect 6425 11396 6429 11452
rect 6429 11396 6485 11452
rect 6485 11396 6489 11452
rect 6425 11392 6489 11396
rect 6505 11452 6569 11456
rect 6505 11396 6509 11452
rect 6509 11396 6565 11452
rect 6565 11396 6569 11452
rect 6505 11392 6569 11396
rect 6585 11452 6649 11456
rect 6585 11396 6589 11452
rect 6589 11396 6645 11452
rect 6645 11396 6649 11452
rect 6585 11392 6649 11396
rect 6665 11452 6729 11456
rect 6665 11396 6669 11452
rect 6669 11396 6725 11452
rect 6725 11396 6729 11452
rect 6665 11392 6729 11396
rect 17372 11452 17436 11456
rect 17372 11396 17376 11452
rect 17376 11396 17432 11452
rect 17432 11396 17436 11452
rect 17372 11392 17436 11396
rect 17452 11452 17516 11456
rect 17452 11396 17456 11452
rect 17456 11396 17512 11452
rect 17512 11396 17516 11452
rect 17452 11392 17516 11396
rect 17532 11452 17596 11456
rect 17532 11396 17536 11452
rect 17536 11396 17592 11452
rect 17592 11396 17596 11452
rect 17532 11392 17596 11396
rect 17612 11452 17676 11456
rect 17612 11396 17616 11452
rect 17616 11396 17672 11452
rect 17672 11396 17676 11452
rect 17612 11392 17676 11396
rect 28319 11452 28383 11456
rect 28319 11396 28323 11452
rect 28323 11396 28379 11452
rect 28379 11396 28383 11452
rect 28319 11392 28383 11396
rect 28399 11452 28463 11456
rect 28399 11396 28403 11452
rect 28403 11396 28459 11452
rect 28459 11396 28463 11452
rect 28399 11392 28463 11396
rect 28479 11452 28543 11456
rect 28479 11396 28483 11452
rect 28483 11396 28539 11452
rect 28539 11396 28543 11452
rect 28479 11392 28543 11396
rect 28559 11452 28623 11456
rect 28559 11396 28563 11452
rect 28563 11396 28619 11452
rect 28619 11396 28623 11452
rect 28559 11392 28623 11396
rect 39266 11452 39330 11456
rect 39266 11396 39270 11452
rect 39270 11396 39326 11452
rect 39326 11396 39330 11452
rect 39266 11392 39330 11396
rect 39346 11452 39410 11456
rect 39346 11396 39350 11452
rect 39350 11396 39406 11452
rect 39406 11396 39410 11452
rect 39346 11392 39410 11396
rect 39426 11452 39490 11456
rect 39426 11396 39430 11452
rect 39430 11396 39486 11452
rect 39486 11396 39490 11452
rect 39426 11392 39490 11396
rect 39506 11452 39570 11456
rect 39506 11396 39510 11452
rect 39510 11396 39566 11452
rect 39566 11396 39570 11452
rect 39506 11392 39570 11396
rect 11898 10908 11962 10912
rect 11898 10852 11902 10908
rect 11902 10852 11958 10908
rect 11958 10852 11962 10908
rect 11898 10848 11962 10852
rect 11978 10908 12042 10912
rect 11978 10852 11982 10908
rect 11982 10852 12038 10908
rect 12038 10852 12042 10908
rect 11978 10848 12042 10852
rect 12058 10908 12122 10912
rect 12058 10852 12062 10908
rect 12062 10852 12118 10908
rect 12118 10852 12122 10908
rect 12058 10848 12122 10852
rect 12138 10908 12202 10912
rect 12138 10852 12142 10908
rect 12142 10852 12198 10908
rect 12198 10852 12202 10908
rect 12138 10848 12202 10852
rect 22845 10908 22909 10912
rect 22845 10852 22849 10908
rect 22849 10852 22905 10908
rect 22905 10852 22909 10908
rect 22845 10848 22909 10852
rect 22925 10908 22989 10912
rect 22925 10852 22929 10908
rect 22929 10852 22985 10908
rect 22985 10852 22989 10908
rect 22925 10848 22989 10852
rect 23005 10908 23069 10912
rect 23005 10852 23009 10908
rect 23009 10852 23065 10908
rect 23065 10852 23069 10908
rect 23005 10848 23069 10852
rect 23085 10908 23149 10912
rect 23085 10852 23089 10908
rect 23089 10852 23145 10908
rect 23145 10852 23149 10908
rect 23085 10848 23149 10852
rect 33792 10908 33856 10912
rect 33792 10852 33796 10908
rect 33796 10852 33852 10908
rect 33852 10852 33856 10908
rect 33792 10848 33856 10852
rect 33872 10908 33936 10912
rect 33872 10852 33876 10908
rect 33876 10852 33932 10908
rect 33932 10852 33936 10908
rect 33872 10848 33936 10852
rect 33952 10908 34016 10912
rect 33952 10852 33956 10908
rect 33956 10852 34012 10908
rect 34012 10852 34016 10908
rect 33952 10848 34016 10852
rect 34032 10908 34096 10912
rect 34032 10852 34036 10908
rect 34036 10852 34092 10908
rect 34092 10852 34096 10908
rect 34032 10848 34096 10852
rect 44739 10908 44803 10912
rect 44739 10852 44743 10908
rect 44743 10852 44799 10908
rect 44799 10852 44803 10908
rect 44739 10848 44803 10852
rect 44819 10908 44883 10912
rect 44819 10852 44823 10908
rect 44823 10852 44879 10908
rect 44879 10852 44883 10908
rect 44819 10848 44883 10852
rect 44899 10908 44963 10912
rect 44899 10852 44903 10908
rect 44903 10852 44959 10908
rect 44959 10852 44963 10908
rect 44899 10848 44963 10852
rect 44979 10908 45043 10912
rect 44979 10852 44983 10908
rect 44983 10852 45039 10908
rect 45039 10852 45043 10908
rect 44979 10848 45043 10852
rect 6425 10364 6489 10368
rect 6425 10308 6429 10364
rect 6429 10308 6485 10364
rect 6485 10308 6489 10364
rect 6425 10304 6489 10308
rect 6505 10364 6569 10368
rect 6505 10308 6509 10364
rect 6509 10308 6565 10364
rect 6565 10308 6569 10364
rect 6505 10304 6569 10308
rect 6585 10364 6649 10368
rect 6585 10308 6589 10364
rect 6589 10308 6645 10364
rect 6645 10308 6649 10364
rect 6585 10304 6649 10308
rect 6665 10364 6729 10368
rect 6665 10308 6669 10364
rect 6669 10308 6725 10364
rect 6725 10308 6729 10364
rect 6665 10304 6729 10308
rect 17372 10364 17436 10368
rect 17372 10308 17376 10364
rect 17376 10308 17432 10364
rect 17432 10308 17436 10364
rect 17372 10304 17436 10308
rect 17452 10364 17516 10368
rect 17452 10308 17456 10364
rect 17456 10308 17512 10364
rect 17512 10308 17516 10364
rect 17452 10304 17516 10308
rect 17532 10364 17596 10368
rect 17532 10308 17536 10364
rect 17536 10308 17592 10364
rect 17592 10308 17596 10364
rect 17532 10304 17596 10308
rect 17612 10364 17676 10368
rect 17612 10308 17616 10364
rect 17616 10308 17672 10364
rect 17672 10308 17676 10364
rect 17612 10304 17676 10308
rect 28319 10364 28383 10368
rect 28319 10308 28323 10364
rect 28323 10308 28379 10364
rect 28379 10308 28383 10364
rect 28319 10304 28383 10308
rect 28399 10364 28463 10368
rect 28399 10308 28403 10364
rect 28403 10308 28459 10364
rect 28459 10308 28463 10364
rect 28399 10304 28463 10308
rect 28479 10364 28543 10368
rect 28479 10308 28483 10364
rect 28483 10308 28539 10364
rect 28539 10308 28543 10364
rect 28479 10304 28543 10308
rect 28559 10364 28623 10368
rect 28559 10308 28563 10364
rect 28563 10308 28619 10364
rect 28619 10308 28623 10364
rect 28559 10304 28623 10308
rect 39266 10364 39330 10368
rect 39266 10308 39270 10364
rect 39270 10308 39326 10364
rect 39326 10308 39330 10364
rect 39266 10304 39330 10308
rect 39346 10364 39410 10368
rect 39346 10308 39350 10364
rect 39350 10308 39406 10364
rect 39406 10308 39410 10364
rect 39346 10304 39410 10308
rect 39426 10364 39490 10368
rect 39426 10308 39430 10364
rect 39430 10308 39486 10364
rect 39486 10308 39490 10364
rect 39426 10304 39490 10308
rect 39506 10364 39570 10368
rect 39506 10308 39510 10364
rect 39510 10308 39566 10364
rect 39566 10308 39570 10364
rect 39506 10304 39570 10308
rect 11898 9820 11962 9824
rect 11898 9764 11902 9820
rect 11902 9764 11958 9820
rect 11958 9764 11962 9820
rect 11898 9760 11962 9764
rect 11978 9820 12042 9824
rect 11978 9764 11982 9820
rect 11982 9764 12038 9820
rect 12038 9764 12042 9820
rect 11978 9760 12042 9764
rect 12058 9820 12122 9824
rect 12058 9764 12062 9820
rect 12062 9764 12118 9820
rect 12118 9764 12122 9820
rect 12058 9760 12122 9764
rect 12138 9820 12202 9824
rect 12138 9764 12142 9820
rect 12142 9764 12198 9820
rect 12198 9764 12202 9820
rect 12138 9760 12202 9764
rect 22845 9820 22909 9824
rect 22845 9764 22849 9820
rect 22849 9764 22905 9820
rect 22905 9764 22909 9820
rect 22845 9760 22909 9764
rect 22925 9820 22989 9824
rect 22925 9764 22929 9820
rect 22929 9764 22985 9820
rect 22985 9764 22989 9820
rect 22925 9760 22989 9764
rect 23005 9820 23069 9824
rect 23005 9764 23009 9820
rect 23009 9764 23065 9820
rect 23065 9764 23069 9820
rect 23005 9760 23069 9764
rect 23085 9820 23149 9824
rect 23085 9764 23089 9820
rect 23089 9764 23145 9820
rect 23145 9764 23149 9820
rect 23085 9760 23149 9764
rect 33792 9820 33856 9824
rect 33792 9764 33796 9820
rect 33796 9764 33852 9820
rect 33852 9764 33856 9820
rect 33792 9760 33856 9764
rect 33872 9820 33936 9824
rect 33872 9764 33876 9820
rect 33876 9764 33932 9820
rect 33932 9764 33936 9820
rect 33872 9760 33936 9764
rect 33952 9820 34016 9824
rect 33952 9764 33956 9820
rect 33956 9764 34012 9820
rect 34012 9764 34016 9820
rect 33952 9760 34016 9764
rect 34032 9820 34096 9824
rect 34032 9764 34036 9820
rect 34036 9764 34092 9820
rect 34092 9764 34096 9820
rect 34032 9760 34096 9764
rect 44739 9820 44803 9824
rect 44739 9764 44743 9820
rect 44743 9764 44799 9820
rect 44799 9764 44803 9820
rect 44739 9760 44803 9764
rect 44819 9820 44883 9824
rect 44819 9764 44823 9820
rect 44823 9764 44879 9820
rect 44879 9764 44883 9820
rect 44819 9760 44883 9764
rect 44899 9820 44963 9824
rect 44899 9764 44903 9820
rect 44903 9764 44959 9820
rect 44959 9764 44963 9820
rect 44899 9760 44963 9764
rect 44979 9820 45043 9824
rect 44979 9764 44983 9820
rect 44983 9764 45039 9820
rect 45039 9764 45043 9820
rect 44979 9760 45043 9764
rect 6425 9276 6489 9280
rect 6425 9220 6429 9276
rect 6429 9220 6485 9276
rect 6485 9220 6489 9276
rect 6425 9216 6489 9220
rect 6505 9276 6569 9280
rect 6505 9220 6509 9276
rect 6509 9220 6565 9276
rect 6565 9220 6569 9276
rect 6505 9216 6569 9220
rect 6585 9276 6649 9280
rect 6585 9220 6589 9276
rect 6589 9220 6645 9276
rect 6645 9220 6649 9276
rect 6585 9216 6649 9220
rect 6665 9276 6729 9280
rect 6665 9220 6669 9276
rect 6669 9220 6725 9276
rect 6725 9220 6729 9276
rect 6665 9216 6729 9220
rect 17372 9276 17436 9280
rect 17372 9220 17376 9276
rect 17376 9220 17432 9276
rect 17432 9220 17436 9276
rect 17372 9216 17436 9220
rect 17452 9276 17516 9280
rect 17452 9220 17456 9276
rect 17456 9220 17512 9276
rect 17512 9220 17516 9276
rect 17452 9216 17516 9220
rect 17532 9276 17596 9280
rect 17532 9220 17536 9276
rect 17536 9220 17592 9276
rect 17592 9220 17596 9276
rect 17532 9216 17596 9220
rect 17612 9276 17676 9280
rect 17612 9220 17616 9276
rect 17616 9220 17672 9276
rect 17672 9220 17676 9276
rect 17612 9216 17676 9220
rect 28319 9276 28383 9280
rect 28319 9220 28323 9276
rect 28323 9220 28379 9276
rect 28379 9220 28383 9276
rect 28319 9216 28383 9220
rect 28399 9276 28463 9280
rect 28399 9220 28403 9276
rect 28403 9220 28459 9276
rect 28459 9220 28463 9276
rect 28399 9216 28463 9220
rect 28479 9276 28543 9280
rect 28479 9220 28483 9276
rect 28483 9220 28539 9276
rect 28539 9220 28543 9276
rect 28479 9216 28543 9220
rect 28559 9276 28623 9280
rect 28559 9220 28563 9276
rect 28563 9220 28619 9276
rect 28619 9220 28623 9276
rect 28559 9216 28623 9220
rect 39266 9276 39330 9280
rect 39266 9220 39270 9276
rect 39270 9220 39326 9276
rect 39326 9220 39330 9276
rect 39266 9216 39330 9220
rect 39346 9276 39410 9280
rect 39346 9220 39350 9276
rect 39350 9220 39406 9276
rect 39406 9220 39410 9276
rect 39346 9216 39410 9220
rect 39426 9276 39490 9280
rect 39426 9220 39430 9276
rect 39430 9220 39486 9276
rect 39486 9220 39490 9276
rect 39426 9216 39490 9220
rect 39506 9276 39570 9280
rect 39506 9220 39510 9276
rect 39510 9220 39566 9276
rect 39566 9220 39570 9276
rect 39506 9216 39570 9220
rect 11898 8732 11962 8736
rect 11898 8676 11902 8732
rect 11902 8676 11958 8732
rect 11958 8676 11962 8732
rect 11898 8672 11962 8676
rect 11978 8732 12042 8736
rect 11978 8676 11982 8732
rect 11982 8676 12038 8732
rect 12038 8676 12042 8732
rect 11978 8672 12042 8676
rect 12058 8732 12122 8736
rect 12058 8676 12062 8732
rect 12062 8676 12118 8732
rect 12118 8676 12122 8732
rect 12058 8672 12122 8676
rect 12138 8732 12202 8736
rect 12138 8676 12142 8732
rect 12142 8676 12198 8732
rect 12198 8676 12202 8732
rect 12138 8672 12202 8676
rect 22845 8732 22909 8736
rect 22845 8676 22849 8732
rect 22849 8676 22905 8732
rect 22905 8676 22909 8732
rect 22845 8672 22909 8676
rect 22925 8732 22989 8736
rect 22925 8676 22929 8732
rect 22929 8676 22985 8732
rect 22985 8676 22989 8732
rect 22925 8672 22989 8676
rect 23005 8732 23069 8736
rect 23005 8676 23009 8732
rect 23009 8676 23065 8732
rect 23065 8676 23069 8732
rect 23005 8672 23069 8676
rect 23085 8732 23149 8736
rect 23085 8676 23089 8732
rect 23089 8676 23145 8732
rect 23145 8676 23149 8732
rect 23085 8672 23149 8676
rect 33792 8732 33856 8736
rect 33792 8676 33796 8732
rect 33796 8676 33852 8732
rect 33852 8676 33856 8732
rect 33792 8672 33856 8676
rect 33872 8732 33936 8736
rect 33872 8676 33876 8732
rect 33876 8676 33932 8732
rect 33932 8676 33936 8732
rect 33872 8672 33936 8676
rect 33952 8732 34016 8736
rect 33952 8676 33956 8732
rect 33956 8676 34012 8732
rect 34012 8676 34016 8732
rect 33952 8672 34016 8676
rect 34032 8732 34096 8736
rect 34032 8676 34036 8732
rect 34036 8676 34092 8732
rect 34092 8676 34096 8732
rect 34032 8672 34096 8676
rect 44739 8732 44803 8736
rect 44739 8676 44743 8732
rect 44743 8676 44799 8732
rect 44799 8676 44803 8732
rect 44739 8672 44803 8676
rect 44819 8732 44883 8736
rect 44819 8676 44823 8732
rect 44823 8676 44879 8732
rect 44879 8676 44883 8732
rect 44819 8672 44883 8676
rect 44899 8732 44963 8736
rect 44899 8676 44903 8732
rect 44903 8676 44959 8732
rect 44959 8676 44963 8732
rect 44899 8672 44963 8676
rect 44979 8732 45043 8736
rect 44979 8676 44983 8732
rect 44983 8676 45039 8732
rect 45039 8676 45043 8732
rect 44979 8672 45043 8676
rect 6425 8188 6489 8192
rect 6425 8132 6429 8188
rect 6429 8132 6485 8188
rect 6485 8132 6489 8188
rect 6425 8128 6489 8132
rect 6505 8188 6569 8192
rect 6505 8132 6509 8188
rect 6509 8132 6565 8188
rect 6565 8132 6569 8188
rect 6505 8128 6569 8132
rect 6585 8188 6649 8192
rect 6585 8132 6589 8188
rect 6589 8132 6645 8188
rect 6645 8132 6649 8188
rect 6585 8128 6649 8132
rect 6665 8188 6729 8192
rect 6665 8132 6669 8188
rect 6669 8132 6725 8188
rect 6725 8132 6729 8188
rect 6665 8128 6729 8132
rect 17372 8188 17436 8192
rect 17372 8132 17376 8188
rect 17376 8132 17432 8188
rect 17432 8132 17436 8188
rect 17372 8128 17436 8132
rect 17452 8188 17516 8192
rect 17452 8132 17456 8188
rect 17456 8132 17512 8188
rect 17512 8132 17516 8188
rect 17452 8128 17516 8132
rect 17532 8188 17596 8192
rect 17532 8132 17536 8188
rect 17536 8132 17592 8188
rect 17592 8132 17596 8188
rect 17532 8128 17596 8132
rect 17612 8188 17676 8192
rect 17612 8132 17616 8188
rect 17616 8132 17672 8188
rect 17672 8132 17676 8188
rect 17612 8128 17676 8132
rect 28319 8188 28383 8192
rect 28319 8132 28323 8188
rect 28323 8132 28379 8188
rect 28379 8132 28383 8188
rect 28319 8128 28383 8132
rect 28399 8188 28463 8192
rect 28399 8132 28403 8188
rect 28403 8132 28459 8188
rect 28459 8132 28463 8188
rect 28399 8128 28463 8132
rect 28479 8188 28543 8192
rect 28479 8132 28483 8188
rect 28483 8132 28539 8188
rect 28539 8132 28543 8188
rect 28479 8128 28543 8132
rect 28559 8188 28623 8192
rect 28559 8132 28563 8188
rect 28563 8132 28619 8188
rect 28619 8132 28623 8188
rect 28559 8128 28623 8132
rect 39266 8188 39330 8192
rect 39266 8132 39270 8188
rect 39270 8132 39326 8188
rect 39326 8132 39330 8188
rect 39266 8128 39330 8132
rect 39346 8188 39410 8192
rect 39346 8132 39350 8188
rect 39350 8132 39406 8188
rect 39406 8132 39410 8188
rect 39346 8128 39410 8132
rect 39426 8188 39490 8192
rect 39426 8132 39430 8188
rect 39430 8132 39486 8188
rect 39486 8132 39490 8188
rect 39426 8128 39490 8132
rect 39506 8188 39570 8192
rect 39506 8132 39510 8188
rect 39510 8132 39566 8188
rect 39566 8132 39570 8188
rect 39506 8128 39570 8132
rect 11898 7644 11962 7648
rect 11898 7588 11902 7644
rect 11902 7588 11958 7644
rect 11958 7588 11962 7644
rect 11898 7584 11962 7588
rect 11978 7644 12042 7648
rect 11978 7588 11982 7644
rect 11982 7588 12038 7644
rect 12038 7588 12042 7644
rect 11978 7584 12042 7588
rect 12058 7644 12122 7648
rect 12058 7588 12062 7644
rect 12062 7588 12118 7644
rect 12118 7588 12122 7644
rect 12058 7584 12122 7588
rect 12138 7644 12202 7648
rect 12138 7588 12142 7644
rect 12142 7588 12198 7644
rect 12198 7588 12202 7644
rect 12138 7584 12202 7588
rect 22845 7644 22909 7648
rect 22845 7588 22849 7644
rect 22849 7588 22905 7644
rect 22905 7588 22909 7644
rect 22845 7584 22909 7588
rect 22925 7644 22989 7648
rect 22925 7588 22929 7644
rect 22929 7588 22985 7644
rect 22985 7588 22989 7644
rect 22925 7584 22989 7588
rect 23005 7644 23069 7648
rect 23005 7588 23009 7644
rect 23009 7588 23065 7644
rect 23065 7588 23069 7644
rect 23005 7584 23069 7588
rect 23085 7644 23149 7648
rect 23085 7588 23089 7644
rect 23089 7588 23145 7644
rect 23145 7588 23149 7644
rect 23085 7584 23149 7588
rect 33792 7644 33856 7648
rect 33792 7588 33796 7644
rect 33796 7588 33852 7644
rect 33852 7588 33856 7644
rect 33792 7584 33856 7588
rect 33872 7644 33936 7648
rect 33872 7588 33876 7644
rect 33876 7588 33932 7644
rect 33932 7588 33936 7644
rect 33872 7584 33936 7588
rect 33952 7644 34016 7648
rect 33952 7588 33956 7644
rect 33956 7588 34012 7644
rect 34012 7588 34016 7644
rect 33952 7584 34016 7588
rect 34032 7644 34096 7648
rect 34032 7588 34036 7644
rect 34036 7588 34092 7644
rect 34092 7588 34096 7644
rect 34032 7584 34096 7588
rect 44739 7644 44803 7648
rect 44739 7588 44743 7644
rect 44743 7588 44799 7644
rect 44799 7588 44803 7644
rect 44739 7584 44803 7588
rect 44819 7644 44883 7648
rect 44819 7588 44823 7644
rect 44823 7588 44879 7644
rect 44879 7588 44883 7644
rect 44819 7584 44883 7588
rect 44899 7644 44963 7648
rect 44899 7588 44903 7644
rect 44903 7588 44959 7644
rect 44959 7588 44963 7644
rect 44899 7584 44963 7588
rect 44979 7644 45043 7648
rect 44979 7588 44983 7644
rect 44983 7588 45039 7644
rect 45039 7588 45043 7644
rect 44979 7584 45043 7588
rect 6425 7100 6489 7104
rect 6425 7044 6429 7100
rect 6429 7044 6485 7100
rect 6485 7044 6489 7100
rect 6425 7040 6489 7044
rect 6505 7100 6569 7104
rect 6505 7044 6509 7100
rect 6509 7044 6565 7100
rect 6565 7044 6569 7100
rect 6505 7040 6569 7044
rect 6585 7100 6649 7104
rect 6585 7044 6589 7100
rect 6589 7044 6645 7100
rect 6645 7044 6649 7100
rect 6585 7040 6649 7044
rect 6665 7100 6729 7104
rect 6665 7044 6669 7100
rect 6669 7044 6725 7100
rect 6725 7044 6729 7100
rect 6665 7040 6729 7044
rect 17372 7100 17436 7104
rect 17372 7044 17376 7100
rect 17376 7044 17432 7100
rect 17432 7044 17436 7100
rect 17372 7040 17436 7044
rect 17452 7100 17516 7104
rect 17452 7044 17456 7100
rect 17456 7044 17512 7100
rect 17512 7044 17516 7100
rect 17452 7040 17516 7044
rect 17532 7100 17596 7104
rect 17532 7044 17536 7100
rect 17536 7044 17592 7100
rect 17592 7044 17596 7100
rect 17532 7040 17596 7044
rect 17612 7100 17676 7104
rect 17612 7044 17616 7100
rect 17616 7044 17672 7100
rect 17672 7044 17676 7100
rect 17612 7040 17676 7044
rect 28319 7100 28383 7104
rect 28319 7044 28323 7100
rect 28323 7044 28379 7100
rect 28379 7044 28383 7100
rect 28319 7040 28383 7044
rect 28399 7100 28463 7104
rect 28399 7044 28403 7100
rect 28403 7044 28459 7100
rect 28459 7044 28463 7100
rect 28399 7040 28463 7044
rect 28479 7100 28543 7104
rect 28479 7044 28483 7100
rect 28483 7044 28539 7100
rect 28539 7044 28543 7100
rect 28479 7040 28543 7044
rect 28559 7100 28623 7104
rect 28559 7044 28563 7100
rect 28563 7044 28619 7100
rect 28619 7044 28623 7100
rect 28559 7040 28623 7044
rect 39266 7100 39330 7104
rect 39266 7044 39270 7100
rect 39270 7044 39326 7100
rect 39326 7044 39330 7100
rect 39266 7040 39330 7044
rect 39346 7100 39410 7104
rect 39346 7044 39350 7100
rect 39350 7044 39406 7100
rect 39406 7044 39410 7100
rect 39346 7040 39410 7044
rect 39426 7100 39490 7104
rect 39426 7044 39430 7100
rect 39430 7044 39486 7100
rect 39486 7044 39490 7100
rect 39426 7040 39490 7044
rect 39506 7100 39570 7104
rect 39506 7044 39510 7100
rect 39510 7044 39566 7100
rect 39566 7044 39570 7100
rect 39506 7040 39570 7044
rect 11898 6556 11962 6560
rect 11898 6500 11902 6556
rect 11902 6500 11958 6556
rect 11958 6500 11962 6556
rect 11898 6496 11962 6500
rect 11978 6556 12042 6560
rect 11978 6500 11982 6556
rect 11982 6500 12038 6556
rect 12038 6500 12042 6556
rect 11978 6496 12042 6500
rect 12058 6556 12122 6560
rect 12058 6500 12062 6556
rect 12062 6500 12118 6556
rect 12118 6500 12122 6556
rect 12058 6496 12122 6500
rect 12138 6556 12202 6560
rect 12138 6500 12142 6556
rect 12142 6500 12198 6556
rect 12198 6500 12202 6556
rect 12138 6496 12202 6500
rect 22845 6556 22909 6560
rect 22845 6500 22849 6556
rect 22849 6500 22905 6556
rect 22905 6500 22909 6556
rect 22845 6496 22909 6500
rect 22925 6556 22989 6560
rect 22925 6500 22929 6556
rect 22929 6500 22985 6556
rect 22985 6500 22989 6556
rect 22925 6496 22989 6500
rect 23005 6556 23069 6560
rect 23005 6500 23009 6556
rect 23009 6500 23065 6556
rect 23065 6500 23069 6556
rect 23005 6496 23069 6500
rect 23085 6556 23149 6560
rect 23085 6500 23089 6556
rect 23089 6500 23145 6556
rect 23145 6500 23149 6556
rect 23085 6496 23149 6500
rect 33792 6556 33856 6560
rect 33792 6500 33796 6556
rect 33796 6500 33852 6556
rect 33852 6500 33856 6556
rect 33792 6496 33856 6500
rect 33872 6556 33936 6560
rect 33872 6500 33876 6556
rect 33876 6500 33932 6556
rect 33932 6500 33936 6556
rect 33872 6496 33936 6500
rect 33952 6556 34016 6560
rect 33952 6500 33956 6556
rect 33956 6500 34012 6556
rect 34012 6500 34016 6556
rect 33952 6496 34016 6500
rect 34032 6556 34096 6560
rect 34032 6500 34036 6556
rect 34036 6500 34092 6556
rect 34092 6500 34096 6556
rect 34032 6496 34096 6500
rect 44739 6556 44803 6560
rect 44739 6500 44743 6556
rect 44743 6500 44799 6556
rect 44799 6500 44803 6556
rect 44739 6496 44803 6500
rect 44819 6556 44883 6560
rect 44819 6500 44823 6556
rect 44823 6500 44879 6556
rect 44879 6500 44883 6556
rect 44819 6496 44883 6500
rect 44899 6556 44963 6560
rect 44899 6500 44903 6556
rect 44903 6500 44959 6556
rect 44959 6500 44963 6556
rect 44899 6496 44963 6500
rect 44979 6556 45043 6560
rect 44979 6500 44983 6556
rect 44983 6500 45039 6556
rect 45039 6500 45043 6556
rect 44979 6496 45043 6500
rect 6425 6012 6489 6016
rect 6425 5956 6429 6012
rect 6429 5956 6485 6012
rect 6485 5956 6489 6012
rect 6425 5952 6489 5956
rect 6505 6012 6569 6016
rect 6505 5956 6509 6012
rect 6509 5956 6565 6012
rect 6565 5956 6569 6012
rect 6505 5952 6569 5956
rect 6585 6012 6649 6016
rect 6585 5956 6589 6012
rect 6589 5956 6645 6012
rect 6645 5956 6649 6012
rect 6585 5952 6649 5956
rect 6665 6012 6729 6016
rect 6665 5956 6669 6012
rect 6669 5956 6725 6012
rect 6725 5956 6729 6012
rect 6665 5952 6729 5956
rect 17372 6012 17436 6016
rect 17372 5956 17376 6012
rect 17376 5956 17432 6012
rect 17432 5956 17436 6012
rect 17372 5952 17436 5956
rect 17452 6012 17516 6016
rect 17452 5956 17456 6012
rect 17456 5956 17512 6012
rect 17512 5956 17516 6012
rect 17452 5952 17516 5956
rect 17532 6012 17596 6016
rect 17532 5956 17536 6012
rect 17536 5956 17592 6012
rect 17592 5956 17596 6012
rect 17532 5952 17596 5956
rect 17612 6012 17676 6016
rect 17612 5956 17616 6012
rect 17616 5956 17672 6012
rect 17672 5956 17676 6012
rect 17612 5952 17676 5956
rect 28319 6012 28383 6016
rect 28319 5956 28323 6012
rect 28323 5956 28379 6012
rect 28379 5956 28383 6012
rect 28319 5952 28383 5956
rect 28399 6012 28463 6016
rect 28399 5956 28403 6012
rect 28403 5956 28459 6012
rect 28459 5956 28463 6012
rect 28399 5952 28463 5956
rect 28479 6012 28543 6016
rect 28479 5956 28483 6012
rect 28483 5956 28539 6012
rect 28539 5956 28543 6012
rect 28479 5952 28543 5956
rect 28559 6012 28623 6016
rect 28559 5956 28563 6012
rect 28563 5956 28619 6012
rect 28619 5956 28623 6012
rect 28559 5952 28623 5956
rect 39266 6012 39330 6016
rect 39266 5956 39270 6012
rect 39270 5956 39326 6012
rect 39326 5956 39330 6012
rect 39266 5952 39330 5956
rect 39346 6012 39410 6016
rect 39346 5956 39350 6012
rect 39350 5956 39406 6012
rect 39406 5956 39410 6012
rect 39346 5952 39410 5956
rect 39426 6012 39490 6016
rect 39426 5956 39430 6012
rect 39430 5956 39486 6012
rect 39486 5956 39490 6012
rect 39426 5952 39490 5956
rect 39506 6012 39570 6016
rect 39506 5956 39510 6012
rect 39510 5956 39566 6012
rect 39566 5956 39570 6012
rect 39506 5952 39570 5956
rect 11898 5468 11962 5472
rect 11898 5412 11902 5468
rect 11902 5412 11958 5468
rect 11958 5412 11962 5468
rect 11898 5408 11962 5412
rect 11978 5468 12042 5472
rect 11978 5412 11982 5468
rect 11982 5412 12038 5468
rect 12038 5412 12042 5468
rect 11978 5408 12042 5412
rect 12058 5468 12122 5472
rect 12058 5412 12062 5468
rect 12062 5412 12118 5468
rect 12118 5412 12122 5468
rect 12058 5408 12122 5412
rect 12138 5468 12202 5472
rect 12138 5412 12142 5468
rect 12142 5412 12198 5468
rect 12198 5412 12202 5468
rect 12138 5408 12202 5412
rect 22845 5468 22909 5472
rect 22845 5412 22849 5468
rect 22849 5412 22905 5468
rect 22905 5412 22909 5468
rect 22845 5408 22909 5412
rect 22925 5468 22989 5472
rect 22925 5412 22929 5468
rect 22929 5412 22985 5468
rect 22985 5412 22989 5468
rect 22925 5408 22989 5412
rect 23005 5468 23069 5472
rect 23005 5412 23009 5468
rect 23009 5412 23065 5468
rect 23065 5412 23069 5468
rect 23005 5408 23069 5412
rect 23085 5468 23149 5472
rect 23085 5412 23089 5468
rect 23089 5412 23145 5468
rect 23145 5412 23149 5468
rect 23085 5408 23149 5412
rect 33792 5468 33856 5472
rect 33792 5412 33796 5468
rect 33796 5412 33852 5468
rect 33852 5412 33856 5468
rect 33792 5408 33856 5412
rect 33872 5468 33936 5472
rect 33872 5412 33876 5468
rect 33876 5412 33932 5468
rect 33932 5412 33936 5468
rect 33872 5408 33936 5412
rect 33952 5468 34016 5472
rect 33952 5412 33956 5468
rect 33956 5412 34012 5468
rect 34012 5412 34016 5468
rect 33952 5408 34016 5412
rect 34032 5468 34096 5472
rect 34032 5412 34036 5468
rect 34036 5412 34092 5468
rect 34092 5412 34096 5468
rect 34032 5408 34096 5412
rect 44739 5468 44803 5472
rect 44739 5412 44743 5468
rect 44743 5412 44799 5468
rect 44799 5412 44803 5468
rect 44739 5408 44803 5412
rect 44819 5468 44883 5472
rect 44819 5412 44823 5468
rect 44823 5412 44879 5468
rect 44879 5412 44883 5468
rect 44819 5408 44883 5412
rect 44899 5468 44963 5472
rect 44899 5412 44903 5468
rect 44903 5412 44959 5468
rect 44959 5412 44963 5468
rect 44899 5408 44963 5412
rect 44979 5468 45043 5472
rect 44979 5412 44983 5468
rect 44983 5412 45039 5468
rect 45039 5412 45043 5468
rect 44979 5408 45043 5412
rect 6425 4924 6489 4928
rect 6425 4868 6429 4924
rect 6429 4868 6485 4924
rect 6485 4868 6489 4924
rect 6425 4864 6489 4868
rect 6505 4924 6569 4928
rect 6505 4868 6509 4924
rect 6509 4868 6565 4924
rect 6565 4868 6569 4924
rect 6505 4864 6569 4868
rect 6585 4924 6649 4928
rect 6585 4868 6589 4924
rect 6589 4868 6645 4924
rect 6645 4868 6649 4924
rect 6585 4864 6649 4868
rect 6665 4924 6729 4928
rect 6665 4868 6669 4924
rect 6669 4868 6725 4924
rect 6725 4868 6729 4924
rect 6665 4864 6729 4868
rect 17372 4924 17436 4928
rect 17372 4868 17376 4924
rect 17376 4868 17432 4924
rect 17432 4868 17436 4924
rect 17372 4864 17436 4868
rect 17452 4924 17516 4928
rect 17452 4868 17456 4924
rect 17456 4868 17512 4924
rect 17512 4868 17516 4924
rect 17452 4864 17516 4868
rect 17532 4924 17596 4928
rect 17532 4868 17536 4924
rect 17536 4868 17592 4924
rect 17592 4868 17596 4924
rect 17532 4864 17596 4868
rect 17612 4924 17676 4928
rect 17612 4868 17616 4924
rect 17616 4868 17672 4924
rect 17672 4868 17676 4924
rect 17612 4864 17676 4868
rect 28319 4924 28383 4928
rect 28319 4868 28323 4924
rect 28323 4868 28379 4924
rect 28379 4868 28383 4924
rect 28319 4864 28383 4868
rect 28399 4924 28463 4928
rect 28399 4868 28403 4924
rect 28403 4868 28459 4924
rect 28459 4868 28463 4924
rect 28399 4864 28463 4868
rect 28479 4924 28543 4928
rect 28479 4868 28483 4924
rect 28483 4868 28539 4924
rect 28539 4868 28543 4924
rect 28479 4864 28543 4868
rect 28559 4924 28623 4928
rect 28559 4868 28563 4924
rect 28563 4868 28619 4924
rect 28619 4868 28623 4924
rect 28559 4864 28623 4868
rect 39266 4924 39330 4928
rect 39266 4868 39270 4924
rect 39270 4868 39326 4924
rect 39326 4868 39330 4924
rect 39266 4864 39330 4868
rect 39346 4924 39410 4928
rect 39346 4868 39350 4924
rect 39350 4868 39406 4924
rect 39406 4868 39410 4924
rect 39346 4864 39410 4868
rect 39426 4924 39490 4928
rect 39426 4868 39430 4924
rect 39430 4868 39486 4924
rect 39486 4868 39490 4924
rect 39426 4864 39490 4868
rect 39506 4924 39570 4928
rect 39506 4868 39510 4924
rect 39510 4868 39566 4924
rect 39566 4868 39570 4924
rect 39506 4864 39570 4868
rect 11898 4380 11962 4384
rect 11898 4324 11902 4380
rect 11902 4324 11958 4380
rect 11958 4324 11962 4380
rect 11898 4320 11962 4324
rect 11978 4380 12042 4384
rect 11978 4324 11982 4380
rect 11982 4324 12038 4380
rect 12038 4324 12042 4380
rect 11978 4320 12042 4324
rect 12058 4380 12122 4384
rect 12058 4324 12062 4380
rect 12062 4324 12118 4380
rect 12118 4324 12122 4380
rect 12058 4320 12122 4324
rect 12138 4380 12202 4384
rect 12138 4324 12142 4380
rect 12142 4324 12198 4380
rect 12198 4324 12202 4380
rect 12138 4320 12202 4324
rect 22845 4380 22909 4384
rect 22845 4324 22849 4380
rect 22849 4324 22905 4380
rect 22905 4324 22909 4380
rect 22845 4320 22909 4324
rect 22925 4380 22989 4384
rect 22925 4324 22929 4380
rect 22929 4324 22985 4380
rect 22985 4324 22989 4380
rect 22925 4320 22989 4324
rect 23005 4380 23069 4384
rect 23005 4324 23009 4380
rect 23009 4324 23065 4380
rect 23065 4324 23069 4380
rect 23005 4320 23069 4324
rect 23085 4380 23149 4384
rect 23085 4324 23089 4380
rect 23089 4324 23145 4380
rect 23145 4324 23149 4380
rect 23085 4320 23149 4324
rect 33792 4380 33856 4384
rect 33792 4324 33796 4380
rect 33796 4324 33852 4380
rect 33852 4324 33856 4380
rect 33792 4320 33856 4324
rect 33872 4380 33936 4384
rect 33872 4324 33876 4380
rect 33876 4324 33932 4380
rect 33932 4324 33936 4380
rect 33872 4320 33936 4324
rect 33952 4380 34016 4384
rect 33952 4324 33956 4380
rect 33956 4324 34012 4380
rect 34012 4324 34016 4380
rect 33952 4320 34016 4324
rect 34032 4380 34096 4384
rect 34032 4324 34036 4380
rect 34036 4324 34092 4380
rect 34092 4324 34096 4380
rect 34032 4320 34096 4324
rect 44739 4380 44803 4384
rect 44739 4324 44743 4380
rect 44743 4324 44799 4380
rect 44799 4324 44803 4380
rect 44739 4320 44803 4324
rect 44819 4380 44883 4384
rect 44819 4324 44823 4380
rect 44823 4324 44879 4380
rect 44879 4324 44883 4380
rect 44819 4320 44883 4324
rect 44899 4380 44963 4384
rect 44899 4324 44903 4380
rect 44903 4324 44959 4380
rect 44959 4324 44963 4380
rect 44899 4320 44963 4324
rect 44979 4380 45043 4384
rect 44979 4324 44983 4380
rect 44983 4324 45039 4380
rect 45039 4324 45043 4380
rect 44979 4320 45043 4324
rect 6425 3836 6489 3840
rect 6425 3780 6429 3836
rect 6429 3780 6485 3836
rect 6485 3780 6489 3836
rect 6425 3776 6489 3780
rect 6505 3836 6569 3840
rect 6505 3780 6509 3836
rect 6509 3780 6565 3836
rect 6565 3780 6569 3836
rect 6505 3776 6569 3780
rect 6585 3836 6649 3840
rect 6585 3780 6589 3836
rect 6589 3780 6645 3836
rect 6645 3780 6649 3836
rect 6585 3776 6649 3780
rect 6665 3836 6729 3840
rect 6665 3780 6669 3836
rect 6669 3780 6725 3836
rect 6725 3780 6729 3836
rect 6665 3776 6729 3780
rect 17372 3836 17436 3840
rect 17372 3780 17376 3836
rect 17376 3780 17432 3836
rect 17432 3780 17436 3836
rect 17372 3776 17436 3780
rect 17452 3836 17516 3840
rect 17452 3780 17456 3836
rect 17456 3780 17512 3836
rect 17512 3780 17516 3836
rect 17452 3776 17516 3780
rect 17532 3836 17596 3840
rect 17532 3780 17536 3836
rect 17536 3780 17592 3836
rect 17592 3780 17596 3836
rect 17532 3776 17596 3780
rect 17612 3836 17676 3840
rect 17612 3780 17616 3836
rect 17616 3780 17672 3836
rect 17672 3780 17676 3836
rect 17612 3776 17676 3780
rect 28319 3836 28383 3840
rect 28319 3780 28323 3836
rect 28323 3780 28379 3836
rect 28379 3780 28383 3836
rect 28319 3776 28383 3780
rect 28399 3836 28463 3840
rect 28399 3780 28403 3836
rect 28403 3780 28459 3836
rect 28459 3780 28463 3836
rect 28399 3776 28463 3780
rect 28479 3836 28543 3840
rect 28479 3780 28483 3836
rect 28483 3780 28539 3836
rect 28539 3780 28543 3836
rect 28479 3776 28543 3780
rect 28559 3836 28623 3840
rect 28559 3780 28563 3836
rect 28563 3780 28619 3836
rect 28619 3780 28623 3836
rect 28559 3776 28623 3780
rect 39266 3836 39330 3840
rect 39266 3780 39270 3836
rect 39270 3780 39326 3836
rect 39326 3780 39330 3836
rect 39266 3776 39330 3780
rect 39346 3836 39410 3840
rect 39346 3780 39350 3836
rect 39350 3780 39406 3836
rect 39406 3780 39410 3836
rect 39346 3776 39410 3780
rect 39426 3836 39490 3840
rect 39426 3780 39430 3836
rect 39430 3780 39486 3836
rect 39486 3780 39490 3836
rect 39426 3776 39490 3780
rect 39506 3836 39570 3840
rect 39506 3780 39510 3836
rect 39510 3780 39566 3836
rect 39566 3780 39570 3836
rect 39506 3776 39570 3780
rect 11898 3292 11962 3296
rect 11898 3236 11902 3292
rect 11902 3236 11958 3292
rect 11958 3236 11962 3292
rect 11898 3232 11962 3236
rect 11978 3292 12042 3296
rect 11978 3236 11982 3292
rect 11982 3236 12038 3292
rect 12038 3236 12042 3292
rect 11978 3232 12042 3236
rect 12058 3292 12122 3296
rect 12058 3236 12062 3292
rect 12062 3236 12118 3292
rect 12118 3236 12122 3292
rect 12058 3232 12122 3236
rect 12138 3292 12202 3296
rect 12138 3236 12142 3292
rect 12142 3236 12198 3292
rect 12198 3236 12202 3292
rect 12138 3232 12202 3236
rect 22845 3292 22909 3296
rect 22845 3236 22849 3292
rect 22849 3236 22905 3292
rect 22905 3236 22909 3292
rect 22845 3232 22909 3236
rect 22925 3292 22989 3296
rect 22925 3236 22929 3292
rect 22929 3236 22985 3292
rect 22985 3236 22989 3292
rect 22925 3232 22989 3236
rect 23005 3292 23069 3296
rect 23005 3236 23009 3292
rect 23009 3236 23065 3292
rect 23065 3236 23069 3292
rect 23005 3232 23069 3236
rect 23085 3292 23149 3296
rect 23085 3236 23089 3292
rect 23089 3236 23145 3292
rect 23145 3236 23149 3292
rect 23085 3232 23149 3236
rect 33792 3292 33856 3296
rect 33792 3236 33796 3292
rect 33796 3236 33852 3292
rect 33852 3236 33856 3292
rect 33792 3232 33856 3236
rect 33872 3292 33936 3296
rect 33872 3236 33876 3292
rect 33876 3236 33932 3292
rect 33932 3236 33936 3292
rect 33872 3232 33936 3236
rect 33952 3292 34016 3296
rect 33952 3236 33956 3292
rect 33956 3236 34012 3292
rect 34012 3236 34016 3292
rect 33952 3232 34016 3236
rect 34032 3292 34096 3296
rect 34032 3236 34036 3292
rect 34036 3236 34092 3292
rect 34092 3236 34096 3292
rect 34032 3232 34096 3236
rect 44739 3292 44803 3296
rect 44739 3236 44743 3292
rect 44743 3236 44799 3292
rect 44799 3236 44803 3292
rect 44739 3232 44803 3236
rect 44819 3292 44883 3296
rect 44819 3236 44823 3292
rect 44823 3236 44879 3292
rect 44879 3236 44883 3292
rect 44819 3232 44883 3236
rect 44899 3292 44963 3296
rect 44899 3236 44903 3292
rect 44903 3236 44959 3292
rect 44959 3236 44963 3292
rect 44899 3232 44963 3236
rect 44979 3292 45043 3296
rect 44979 3236 44983 3292
rect 44983 3236 45039 3292
rect 45039 3236 45043 3292
rect 44979 3232 45043 3236
rect 6425 2748 6489 2752
rect 6425 2692 6429 2748
rect 6429 2692 6485 2748
rect 6485 2692 6489 2748
rect 6425 2688 6489 2692
rect 6505 2748 6569 2752
rect 6505 2692 6509 2748
rect 6509 2692 6565 2748
rect 6565 2692 6569 2748
rect 6505 2688 6569 2692
rect 6585 2748 6649 2752
rect 6585 2692 6589 2748
rect 6589 2692 6645 2748
rect 6645 2692 6649 2748
rect 6585 2688 6649 2692
rect 6665 2748 6729 2752
rect 6665 2692 6669 2748
rect 6669 2692 6725 2748
rect 6725 2692 6729 2748
rect 6665 2688 6729 2692
rect 17372 2748 17436 2752
rect 17372 2692 17376 2748
rect 17376 2692 17432 2748
rect 17432 2692 17436 2748
rect 17372 2688 17436 2692
rect 17452 2748 17516 2752
rect 17452 2692 17456 2748
rect 17456 2692 17512 2748
rect 17512 2692 17516 2748
rect 17452 2688 17516 2692
rect 17532 2748 17596 2752
rect 17532 2692 17536 2748
rect 17536 2692 17592 2748
rect 17592 2692 17596 2748
rect 17532 2688 17596 2692
rect 17612 2748 17676 2752
rect 17612 2692 17616 2748
rect 17616 2692 17672 2748
rect 17672 2692 17676 2748
rect 17612 2688 17676 2692
rect 28319 2748 28383 2752
rect 28319 2692 28323 2748
rect 28323 2692 28379 2748
rect 28379 2692 28383 2748
rect 28319 2688 28383 2692
rect 28399 2748 28463 2752
rect 28399 2692 28403 2748
rect 28403 2692 28459 2748
rect 28459 2692 28463 2748
rect 28399 2688 28463 2692
rect 28479 2748 28543 2752
rect 28479 2692 28483 2748
rect 28483 2692 28539 2748
rect 28539 2692 28543 2748
rect 28479 2688 28543 2692
rect 28559 2748 28623 2752
rect 28559 2692 28563 2748
rect 28563 2692 28619 2748
rect 28619 2692 28623 2748
rect 28559 2688 28623 2692
rect 39266 2748 39330 2752
rect 39266 2692 39270 2748
rect 39270 2692 39326 2748
rect 39326 2692 39330 2748
rect 39266 2688 39330 2692
rect 39346 2748 39410 2752
rect 39346 2692 39350 2748
rect 39350 2692 39406 2748
rect 39406 2692 39410 2748
rect 39346 2688 39410 2692
rect 39426 2748 39490 2752
rect 39426 2692 39430 2748
rect 39430 2692 39486 2748
rect 39486 2692 39490 2748
rect 39426 2688 39490 2692
rect 39506 2748 39570 2752
rect 39506 2692 39510 2748
rect 39510 2692 39566 2748
rect 39566 2692 39570 2748
rect 39506 2688 39570 2692
rect 11898 2204 11962 2208
rect 11898 2148 11902 2204
rect 11902 2148 11958 2204
rect 11958 2148 11962 2204
rect 11898 2144 11962 2148
rect 11978 2204 12042 2208
rect 11978 2148 11982 2204
rect 11982 2148 12038 2204
rect 12038 2148 12042 2204
rect 11978 2144 12042 2148
rect 12058 2204 12122 2208
rect 12058 2148 12062 2204
rect 12062 2148 12118 2204
rect 12118 2148 12122 2204
rect 12058 2144 12122 2148
rect 12138 2204 12202 2208
rect 12138 2148 12142 2204
rect 12142 2148 12198 2204
rect 12198 2148 12202 2204
rect 12138 2144 12202 2148
rect 22845 2204 22909 2208
rect 22845 2148 22849 2204
rect 22849 2148 22905 2204
rect 22905 2148 22909 2204
rect 22845 2144 22909 2148
rect 22925 2204 22989 2208
rect 22925 2148 22929 2204
rect 22929 2148 22985 2204
rect 22985 2148 22989 2204
rect 22925 2144 22989 2148
rect 23005 2204 23069 2208
rect 23005 2148 23009 2204
rect 23009 2148 23065 2204
rect 23065 2148 23069 2204
rect 23005 2144 23069 2148
rect 23085 2204 23149 2208
rect 23085 2148 23089 2204
rect 23089 2148 23145 2204
rect 23145 2148 23149 2204
rect 23085 2144 23149 2148
rect 33792 2204 33856 2208
rect 33792 2148 33796 2204
rect 33796 2148 33852 2204
rect 33852 2148 33856 2204
rect 33792 2144 33856 2148
rect 33872 2204 33936 2208
rect 33872 2148 33876 2204
rect 33876 2148 33932 2204
rect 33932 2148 33936 2204
rect 33872 2144 33936 2148
rect 33952 2204 34016 2208
rect 33952 2148 33956 2204
rect 33956 2148 34012 2204
rect 34012 2148 34016 2204
rect 33952 2144 34016 2148
rect 34032 2204 34096 2208
rect 34032 2148 34036 2204
rect 34036 2148 34092 2204
rect 34092 2148 34096 2204
rect 34032 2144 34096 2148
rect 44739 2204 44803 2208
rect 44739 2148 44743 2204
rect 44743 2148 44799 2204
rect 44799 2148 44803 2204
rect 44739 2144 44803 2148
rect 44819 2204 44883 2208
rect 44819 2148 44823 2204
rect 44823 2148 44879 2204
rect 44879 2148 44883 2204
rect 44819 2144 44883 2148
rect 44899 2204 44963 2208
rect 44899 2148 44903 2204
rect 44903 2148 44959 2204
rect 44959 2148 44963 2204
rect 44899 2144 44963 2148
rect 44979 2204 45043 2208
rect 44979 2148 44983 2204
rect 44983 2148 45039 2204
rect 45039 2148 45043 2204
rect 44979 2144 45043 2148
<< metal4 >>
rect 6417 16896 6737 17456
rect 6417 16832 6425 16896
rect 6489 16832 6505 16896
rect 6569 16832 6585 16896
rect 6649 16832 6665 16896
rect 6729 16832 6737 16896
rect 6417 15808 6737 16832
rect 6417 15744 6425 15808
rect 6489 15744 6505 15808
rect 6569 15744 6585 15808
rect 6649 15744 6665 15808
rect 6729 15744 6737 15808
rect 6417 14720 6737 15744
rect 6417 14656 6425 14720
rect 6489 14656 6505 14720
rect 6569 14656 6585 14720
rect 6649 14656 6665 14720
rect 6729 14656 6737 14720
rect 6417 13632 6737 14656
rect 6417 13568 6425 13632
rect 6489 13568 6505 13632
rect 6569 13568 6585 13632
rect 6649 13568 6665 13632
rect 6729 13568 6737 13632
rect 6417 12544 6737 13568
rect 6417 12480 6425 12544
rect 6489 12480 6505 12544
rect 6569 12480 6585 12544
rect 6649 12480 6665 12544
rect 6729 12480 6737 12544
rect 6417 11456 6737 12480
rect 6417 11392 6425 11456
rect 6489 11392 6505 11456
rect 6569 11392 6585 11456
rect 6649 11392 6665 11456
rect 6729 11392 6737 11456
rect 6417 10368 6737 11392
rect 6417 10304 6425 10368
rect 6489 10304 6505 10368
rect 6569 10304 6585 10368
rect 6649 10304 6665 10368
rect 6729 10304 6737 10368
rect 6417 9280 6737 10304
rect 6417 9216 6425 9280
rect 6489 9216 6505 9280
rect 6569 9216 6585 9280
rect 6649 9216 6665 9280
rect 6729 9216 6737 9280
rect 6417 8192 6737 9216
rect 6417 8128 6425 8192
rect 6489 8128 6505 8192
rect 6569 8128 6585 8192
rect 6649 8128 6665 8192
rect 6729 8128 6737 8192
rect 6417 7104 6737 8128
rect 6417 7040 6425 7104
rect 6489 7040 6505 7104
rect 6569 7040 6585 7104
rect 6649 7040 6665 7104
rect 6729 7040 6737 7104
rect 6417 6016 6737 7040
rect 6417 5952 6425 6016
rect 6489 5952 6505 6016
rect 6569 5952 6585 6016
rect 6649 5952 6665 6016
rect 6729 5952 6737 6016
rect 6417 4928 6737 5952
rect 6417 4864 6425 4928
rect 6489 4864 6505 4928
rect 6569 4864 6585 4928
rect 6649 4864 6665 4928
rect 6729 4864 6737 4928
rect 6417 3840 6737 4864
rect 6417 3776 6425 3840
rect 6489 3776 6505 3840
rect 6569 3776 6585 3840
rect 6649 3776 6665 3840
rect 6729 3776 6737 3840
rect 6417 2752 6737 3776
rect 6417 2688 6425 2752
rect 6489 2688 6505 2752
rect 6569 2688 6585 2752
rect 6649 2688 6665 2752
rect 6729 2688 6737 2752
rect 6417 2128 6737 2688
rect 11890 17440 12210 17456
rect 11890 17376 11898 17440
rect 11962 17376 11978 17440
rect 12042 17376 12058 17440
rect 12122 17376 12138 17440
rect 12202 17376 12210 17440
rect 11890 16352 12210 17376
rect 11890 16288 11898 16352
rect 11962 16288 11978 16352
rect 12042 16288 12058 16352
rect 12122 16288 12138 16352
rect 12202 16288 12210 16352
rect 11890 15264 12210 16288
rect 11890 15200 11898 15264
rect 11962 15200 11978 15264
rect 12042 15200 12058 15264
rect 12122 15200 12138 15264
rect 12202 15200 12210 15264
rect 11890 14176 12210 15200
rect 11890 14112 11898 14176
rect 11962 14112 11978 14176
rect 12042 14112 12058 14176
rect 12122 14112 12138 14176
rect 12202 14112 12210 14176
rect 11890 13088 12210 14112
rect 11890 13024 11898 13088
rect 11962 13024 11978 13088
rect 12042 13024 12058 13088
rect 12122 13024 12138 13088
rect 12202 13024 12210 13088
rect 11890 12000 12210 13024
rect 11890 11936 11898 12000
rect 11962 11936 11978 12000
rect 12042 11936 12058 12000
rect 12122 11936 12138 12000
rect 12202 11936 12210 12000
rect 11890 10912 12210 11936
rect 11890 10848 11898 10912
rect 11962 10848 11978 10912
rect 12042 10848 12058 10912
rect 12122 10848 12138 10912
rect 12202 10848 12210 10912
rect 11890 9824 12210 10848
rect 11890 9760 11898 9824
rect 11962 9760 11978 9824
rect 12042 9760 12058 9824
rect 12122 9760 12138 9824
rect 12202 9760 12210 9824
rect 11890 8736 12210 9760
rect 11890 8672 11898 8736
rect 11962 8672 11978 8736
rect 12042 8672 12058 8736
rect 12122 8672 12138 8736
rect 12202 8672 12210 8736
rect 11890 7648 12210 8672
rect 11890 7584 11898 7648
rect 11962 7584 11978 7648
rect 12042 7584 12058 7648
rect 12122 7584 12138 7648
rect 12202 7584 12210 7648
rect 11890 6560 12210 7584
rect 11890 6496 11898 6560
rect 11962 6496 11978 6560
rect 12042 6496 12058 6560
rect 12122 6496 12138 6560
rect 12202 6496 12210 6560
rect 11890 5472 12210 6496
rect 11890 5408 11898 5472
rect 11962 5408 11978 5472
rect 12042 5408 12058 5472
rect 12122 5408 12138 5472
rect 12202 5408 12210 5472
rect 11890 4384 12210 5408
rect 11890 4320 11898 4384
rect 11962 4320 11978 4384
rect 12042 4320 12058 4384
rect 12122 4320 12138 4384
rect 12202 4320 12210 4384
rect 11890 3296 12210 4320
rect 11890 3232 11898 3296
rect 11962 3232 11978 3296
rect 12042 3232 12058 3296
rect 12122 3232 12138 3296
rect 12202 3232 12210 3296
rect 11890 2208 12210 3232
rect 11890 2144 11898 2208
rect 11962 2144 11978 2208
rect 12042 2144 12058 2208
rect 12122 2144 12138 2208
rect 12202 2144 12210 2208
rect 11890 2128 12210 2144
rect 17364 16896 17684 17456
rect 17364 16832 17372 16896
rect 17436 16832 17452 16896
rect 17516 16832 17532 16896
rect 17596 16832 17612 16896
rect 17676 16832 17684 16896
rect 17364 15808 17684 16832
rect 17364 15744 17372 15808
rect 17436 15744 17452 15808
rect 17516 15744 17532 15808
rect 17596 15744 17612 15808
rect 17676 15744 17684 15808
rect 17364 14720 17684 15744
rect 17364 14656 17372 14720
rect 17436 14656 17452 14720
rect 17516 14656 17532 14720
rect 17596 14656 17612 14720
rect 17676 14656 17684 14720
rect 17364 13632 17684 14656
rect 17364 13568 17372 13632
rect 17436 13568 17452 13632
rect 17516 13568 17532 13632
rect 17596 13568 17612 13632
rect 17676 13568 17684 13632
rect 17364 12544 17684 13568
rect 17364 12480 17372 12544
rect 17436 12480 17452 12544
rect 17516 12480 17532 12544
rect 17596 12480 17612 12544
rect 17676 12480 17684 12544
rect 17364 11456 17684 12480
rect 17364 11392 17372 11456
rect 17436 11392 17452 11456
rect 17516 11392 17532 11456
rect 17596 11392 17612 11456
rect 17676 11392 17684 11456
rect 17364 10368 17684 11392
rect 17364 10304 17372 10368
rect 17436 10304 17452 10368
rect 17516 10304 17532 10368
rect 17596 10304 17612 10368
rect 17676 10304 17684 10368
rect 17364 9280 17684 10304
rect 17364 9216 17372 9280
rect 17436 9216 17452 9280
rect 17516 9216 17532 9280
rect 17596 9216 17612 9280
rect 17676 9216 17684 9280
rect 17364 8192 17684 9216
rect 17364 8128 17372 8192
rect 17436 8128 17452 8192
rect 17516 8128 17532 8192
rect 17596 8128 17612 8192
rect 17676 8128 17684 8192
rect 17364 7104 17684 8128
rect 17364 7040 17372 7104
rect 17436 7040 17452 7104
rect 17516 7040 17532 7104
rect 17596 7040 17612 7104
rect 17676 7040 17684 7104
rect 17364 6016 17684 7040
rect 17364 5952 17372 6016
rect 17436 5952 17452 6016
rect 17516 5952 17532 6016
rect 17596 5952 17612 6016
rect 17676 5952 17684 6016
rect 17364 4928 17684 5952
rect 17364 4864 17372 4928
rect 17436 4864 17452 4928
rect 17516 4864 17532 4928
rect 17596 4864 17612 4928
rect 17676 4864 17684 4928
rect 17364 3840 17684 4864
rect 17364 3776 17372 3840
rect 17436 3776 17452 3840
rect 17516 3776 17532 3840
rect 17596 3776 17612 3840
rect 17676 3776 17684 3840
rect 17364 2752 17684 3776
rect 17364 2688 17372 2752
rect 17436 2688 17452 2752
rect 17516 2688 17532 2752
rect 17596 2688 17612 2752
rect 17676 2688 17684 2752
rect 17364 2128 17684 2688
rect 22837 17440 23157 17456
rect 22837 17376 22845 17440
rect 22909 17376 22925 17440
rect 22989 17376 23005 17440
rect 23069 17376 23085 17440
rect 23149 17376 23157 17440
rect 22837 16352 23157 17376
rect 22837 16288 22845 16352
rect 22909 16288 22925 16352
rect 22989 16288 23005 16352
rect 23069 16288 23085 16352
rect 23149 16288 23157 16352
rect 22837 15264 23157 16288
rect 22837 15200 22845 15264
rect 22909 15200 22925 15264
rect 22989 15200 23005 15264
rect 23069 15200 23085 15264
rect 23149 15200 23157 15264
rect 22837 14176 23157 15200
rect 22837 14112 22845 14176
rect 22909 14112 22925 14176
rect 22989 14112 23005 14176
rect 23069 14112 23085 14176
rect 23149 14112 23157 14176
rect 22837 13088 23157 14112
rect 22837 13024 22845 13088
rect 22909 13024 22925 13088
rect 22989 13024 23005 13088
rect 23069 13024 23085 13088
rect 23149 13024 23157 13088
rect 22837 12000 23157 13024
rect 22837 11936 22845 12000
rect 22909 11936 22925 12000
rect 22989 11936 23005 12000
rect 23069 11936 23085 12000
rect 23149 11936 23157 12000
rect 22837 10912 23157 11936
rect 22837 10848 22845 10912
rect 22909 10848 22925 10912
rect 22989 10848 23005 10912
rect 23069 10848 23085 10912
rect 23149 10848 23157 10912
rect 22837 9824 23157 10848
rect 22837 9760 22845 9824
rect 22909 9760 22925 9824
rect 22989 9760 23005 9824
rect 23069 9760 23085 9824
rect 23149 9760 23157 9824
rect 22837 8736 23157 9760
rect 22837 8672 22845 8736
rect 22909 8672 22925 8736
rect 22989 8672 23005 8736
rect 23069 8672 23085 8736
rect 23149 8672 23157 8736
rect 22837 7648 23157 8672
rect 22837 7584 22845 7648
rect 22909 7584 22925 7648
rect 22989 7584 23005 7648
rect 23069 7584 23085 7648
rect 23149 7584 23157 7648
rect 22837 6560 23157 7584
rect 22837 6496 22845 6560
rect 22909 6496 22925 6560
rect 22989 6496 23005 6560
rect 23069 6496 23085 6560
rect 23149 6496 23157 6560
rect 22837 5472 23157 6496
rect 22837 5408 22845 5472
rect 22909 5408 22925 5472
rect 22989 5408 23005 5472
rect 23069 5408 23085 5472
rect 23149 5408 23157 5472
rect 22837 4384 23157 5408
rect 22837 4320 22845 4384
rect 22909 4320 22925 4384
rect 22989 4320 23005 4384
rect 23069 4320 23085 4384
rect 23149 4320 23157 4384
rect 22837 3296 23157 4320
rect 22837 3232 22845 3296
rect 22909 3232 22925 3296
rect 22989 3232 23005 3296
rect 23069 3232 23085 3296
rect 23149 3232 23157 3296
rect 22837 2208 23157 3232
rect 22837 2144 22845 2208
rect 22909 2144 22925 2208
rect 22989 2144 23005 2208
rect 23069 2144 23085 2208
rect 23149 2144 23157 2208
rect 22837 2128 23157 2144
rect 28311 16896 28631 17456
rect 28311 16832 28319 16896
rect 28383 16832 28399 16896
rect 28463 16832 28479 16896
rect 28543 16832 28559 16896
rect 28623 16832 28631 16896
rect 28311 15808 28631 16832
rect 28311 15744 28319 15808
rect 28383 15744 28399 15808
rect 28463 15744 28479 15808
rect 28543 15744 28559 15808
rect 28623 15744 28631 15808
rect 28311 14720 28631 15744
rect 28311 14656 28319 14720
rect 28383 14656 28399 14720
rect 28463 14656 28479 14720
rect 28543 14656 28559 14720
rect 28623 14656 28631 14720
rect 28311 13632 28631 14656
rect 28311 13568 28319 13632
rect 28383 13568 28399 13632
rect 28463 13568 28479 13632
rect 28543 13568 28559 13632
rect 28623 13568 28631 13632
rect 28311 12544 28631 13568
rect 28311 12480 28319 12544
rect 28383 12480 28399 12544
rect 28463 12480 28479 12544
rect 28543 12480 28559 12544
rect 28623 12480 28631 12544
rect 28311 11456 28631 12480
rect 28311 11392 28319 11456
rect 28383 11392 28399 11456
rect 28463 11392 28479 11456
rect 28543 11392 28559 11456
rect 28623 11392 28631 11456
rect 28311 10368 28631 11392
rect 28311 10304 28319 10368
rect 28383 10304 28399 10368
rect 28463 10304 28479 10368
rect 28543 10304 28559 10368
rect 28623 10304 28631 10368
rect 28311 9280 28631 10304
rect 28311 9216 28319 9280
rect 28383 9216 28399 9280
rect 28463 9216 28479 9280
rect 28543 9216 28559 9280
rect 28623 9216 28631 9280
rect 28311 8192 28631 9216
rect 28311 8128 28319 8192
rect 28383 8128 28399 8192
rect 28463 8128 28479 8192
rect 28543 8128 28559 8192
rect 28623 8128 28631 8192
rect 28311 7104 28631 8128
rect 28311 7040 28319 7104
rect 28383 7040 28399 7104
rect 28463 7040 28479 7104
rect 28543 7040 28559 7104
rect 28623 7040 28631 7104
rect 28311 6016 28631 7040
rect 28311 5952 28319 6016
rect 28383 5952 28399 6016
rect 28463 5952 28479 6016
rect 28543 5952 28559 6016
rect 28623 5952 28631 6016
rect 28311 4928 28631 5952
rect 28311 4864 28319 4928
rect 28383 4864 28399 4928
rect 28463 4864 28479 4928
rect 28543 4864 28559 4928
rect 28623 4864 28631 4928
rect 28311 3840 28631 4864
rect 28311 3776 28319 3840
rect 28383 3776 28399 3840
rect 28463 3776 28479 3840
rect 28543 3776 28559 3840
rect 28623 3776 28631 3840
rect 28311 2752 28631 3776
rect 28311 2688 28319 2752
rect 28383 2688 28399 2752
rect 28463 2688 28479 2752
rect 28543 2688 28559 2752
rect 28623 2688 28631 2752
rect 28311 2128 28631 2688
rect 33784 17440 34104 17456
rect 33784 17376 33792 17440
rect 33856 17376 33872 17440
rect 33936 17376 33952 17440
rect 34016 17376 34032 17440
rect 34096 17376 34104 17440
rect 33784 16352 34104 17376
rect 33784 16288 33792 16352
rect 33856 16288 33872 16352
rect 33936 16288 33952 16352
rect 34016 16288 34032 16352
rect 34096 16288 34104 16352
rect 33784 15264 34104 16288
rect 33784 15200 33792 15264
rect 33856 15200 33872 15264
rect 33936 15200 33952 15264
rect 34016 15200 34032 15264
rect 34096 15200 34104 15264
rect 33784 14176 34104 15200
rect 33784 14112 33792 14176
rect 33856 14112 33872 14176
rect 33936 14112 33952 14176
rect 34016 14112 34032 14176
rect 34096 14112 34104 14176
rect 33784 13088 34104 14112
rect 33784 13024 33792 13088
rect 33856 13024 33872 13088
rect 33936 13024 33952 13088
rect 34016 13024 34032 13088
rect 34096 13024 34104 13088
rect 33784 12000 34104 13024
rect 33784 11936 33792 12000
rect 33856 11936 33872 12000
rect 33936 11936 33952 12000
rect 34016 11936 34032 12000
rect 34096 11936 34104 12000
rect 33784 10912 34104 11936
rect 33784 10848 33792 10912
rect 33856 10848 33872 10912
rect 33936 10848 33952 10912
rect 34016 10848 34032 10912
rect 34096 10848 34104 10912
rect 33784 9824 34104 10848
rect 33784 9760 33792 9824
rect 33856 9760 33872 9824
rect 33936 9760 33952 9824
rect 34016 9760 34032 9824
rect 34096 9760 34104 9824
rect 33784 8736 34104 9760
rect 33784 8672 33792 8736
rect 33856 8672 33872 8736
rect 33936 8672 33952 8736
rect 34016 8672 34032 8736
rect 34096 8672 34104 8736
rect 33784 7648 34104 8672
rect 33784 7584 33792 7648
rect 33856 7584 33872 7648
rect 33936 7584 33952 7648
rect 34016 7584 34032 7648
rect 34096 7584 34104 7648
rect 33784 6560 34104 7584
rect 33784 6496 33792 6560
rect 33856 6496 33872 6560
rect 33936 6496 33952 6560
rect 34016 6496 34032 6560
rect 34096 6496 34104 6560
rect 33784 5472 34104 6496
rect 33784 5408 33792 5472
rect 33856 5408 33872 5472
rect 33936 5408 33952 5472
rect 34016 5408 34032 5472
rect 34096 5408 34104 5472
rect 33784 4384 34104 5408
rect 33784 4320 33792 4384
rect 33856 4320 33872 4384
rect 33936 4320 33952 4384
rect 34016 4320 34032 4384
rect 34096 4320 34104 4384
rect 33784 3296 34104 4320
rect 33784 3232 33792 3296
rect 33856 3232 33872 3296
rect 33936 3232 33952 3296
rect 34016 3232 34032 3296
rect 34096 3232 34104 3296
rect 33784 2208 34104 3232
rect 33784 2144 33792 2208
rect 33856 2144 33872 2208
rect 33936 2144 33952 2208
rect 34016 2144 34032 2208
rect 34096 2144 34104 2208
rect 33784 2128 34104 2144
rect 39258 16896 39578 17456
rect 39258 16832 39266 16896
rect 39330 16832 39346 16896
rect 39410 16832 39426 16896
rect 39490 16832 39506 16896
rect 39570 16832 39578 16896
rect 39258 15808 39578 16832
rect 39258 15744 39266 15808
rect 39330 15744 39346 15808
rect 39410 15744 39426 15808
rect 39490 15744 39506 15808
rect 39570 15744 39578 15808
rect 39258 14720 39578 15744
rect 39258 14656 39266 14720
rect 39330 14656 39346 14720
rect 39410 14656 39426 14720
rect 39490 14656 39506 14720
rect 39570 14656 39578 14720
rect 39258 13632 39578 14656
rect 39258 13568 39266 13632
rect 39330 13568 39346 13632
rect 39410 13568 39426 13632
rect 39490 13568 39506 13632
rect 39570 13568 39578 13632
rect 39258 12544 39578 13568
rect 39258 12480 39266 12544
rect 39330 12480 39346 12544
rect 39410 12480 39426 12544
rect 39490 12480 39506 12544
rect 39570 12480 39578 12544
rect 39258 11456 39578 12480
rect 39258 11392 39266 11456
rect 39330 11392 39346 11456
rect 39410 11392 39426 11456
rect 39490 11392 39506 11456
rect 39570 11392 39578 11456
rect 39258 10368 39578 11392
rect 39258 10304 39266 10368
rect 39330 10304 39346 10368
rect 39410 10304 39426 10368
rect 39490 10304 39506 10368
rect 39570 10304 39578 10368
rect 39258 9280 39578 10304
rect 39258 9216 39266 9280
rect 39330 9216 39346 9280
rect 39410 9216 39426 9280
rect 39490 9216 39506 9280
rect 39570 9216 39578 9280
rect 39258 8192 39578 9216
rect 39258 8128 39266 8192
rect 39330 8128 39346 8192
rect 39410 8128 39426 8192
rect 39490 8128 39506 8192
rect 39570 8128 39578 8192
rect 39258 7104 39578 8128
rect 39258 7040 39266 7104
rect 39330 7040 39346 7104
rect 39410 7040 39426 7104
rect 39490 7040 39506 7104
rect 39570 7040 39578 7104
rect 39258 6016 39578 7040
rect 39258 5952 39266 6016
rect 39330 5952 39346 6016
rect 39410 5952 39426 6016
rect 39490 5952 39506 6016
rect 39570 5952 39578 6016
rect 39258 4928 39578 5952
rect 39258 4864 39266 4928
rect 39330 4864 39346 4928
rect 39410 4864 39426 4928
rect 39490 4864 39506 4928
rect 39570 4864 39578 4928
rect 39258 3840 39578 4864
rect 39258 3776 39266 3840
rect 39330 3776 39346 3840
rect 39410 3776 39426 3840
rect 39490 3776 39506 3840
rect 39570 3776 39578 3840
rect 39258 2752 39578 3776
rect 39258 2688 39266 2752
rect 39330 2688 39346 2752
rect 39410 2688 39426 2752
rect 39490 2688 39506 2752
rect 39570 2688 39578 2752
rect 39258 2128 39578 2688
rect 44731 17440 45051 17456
rect 44731 17376 44739 17440
rect 44803 17376 44819 17440
rect 44883 17376 44899 17440
rect 44963 17376 44979 17440
rect 45043 17376 45051 17440
rect 44731 16352 45051 17376
rect 44731 16288 44739 16352
rect 44803 16288 44819 16352
rect 44883 16288 44899 16352
rect 44963 16288 44979 16352
rect 45043 16288 45051 16352
rect 44731 15264 45051 16288
rect 44731 15200 44739 15264
rect 44803 15200 44819 15264
rect 44883 15200 44899 15264
rect 44963 15200 44979 15264
rect 45043 15200 45051 15264
rect 44731 14176 45051 15200
rect 44731 14112 44739 14176
rect 44803 14112 44819 14176
rect 44883 14112 44899 14176
rect 44963 14112 44979 14176
rect 45043 14112 45051 14176
rect 44731 13088 45051 14112
rect 44731 13024 44739 13088
rect 44803 13024 44819 13088
rect 44883 13024 44899 13088
rect 44963 13024 44979 13088
rect 45043 13024 45051 13088
rect 44731 12000 45051 13024
rect 44731 11936 44739 12000
rect 44803 11936 44819 12000
rect 44883 11936 44899 12000
rect 44963 11936 44979 12000
rect 45043 11936 45051 12000
rect 44731 10912 45051 11936
rect 44731 10848 44739 10912
rect 44803 10848 44819 10912
rect 44883 10848 44899 10912
rect 44963 10848 44979 10912
rect 45043 10848 45051 10912
rect 44731 9824 45051 10848
rect 44731 9760 44739 9824
rect 44803 9760 44819 9824
rect 44883 9760 44899 9824
rect 44963 9760 44979 9824
rect 45043 9760 45051 9824
rect 44731 8736 45051 9760
rect 44731 8672 44739 8736
rect 44803 8672 44819 8736
rect 44883 8672 44899 8736
rect 44963 8672 44979 8736
rect 45043 8672 45051 8736
rect 44731 7648 45051 8672
rect 44731 7584 44739 7648
rect 44803 7584 44819 7648
rect 44883 7584 44899 7648
rect 44963 7584 44979 7648
rect 45043 7584 45051 7648
rect 44731 6560 45051 7584
rect 44731 6496 44739 6560
rect 44803 6496 44819 6560
rect 44883 6496 44899 6560
rect 44963 6496 44979 6560
rect 45043 6496 45051 6560
rect 44731 5472 45051 6496
rect 44731 5408 44739 5472
rect 44803 5408 44819 5472
rect 44883 5408 44899 5472
rect 44963 5408 44979 5472
rect 45043 5408 45051 5472
rect 44731 4384 45051 5408
rect 44731 4320 44739 4384
rect 44803 4320 44819 4384
rect 44883 4320 44899 4384
rect 44963 4320 44979 4384
rect 45043 4320 45051 4384
rect 44731 3296 45051 4320
rect 44731 3232 44739 3296
rect 44803 3232 44819 3296
rect 44883 3232 44899 3296
rect 44963 3232 44979 3296
rect 45043 3232 45051 3296
rect 44731 2208 45051 3232
rect 44731 2144 44739 2208
rect 44803 2144 44819 2208
rect 44883 2144 44899 2208
rect 44963 2144 44979 2208
rect 45043 2144 45051 2208
rect 44731 2128 45051 2144
use sky130_fd_sc_hd__diode_2  ANTENNA_1 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 32844 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1676037725
transform -1 0 8004 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 1380 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 1840 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 2484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29
timestamp 1676037725
transform 1 0 3772 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34
timestamp 1676037725
transform 1 0 4232 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41
timestamp 1676037725
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57
timestamp 1676037725
transform 1 0 6348 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_69
timestamp 1676037725
transform 1 0 7452 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_76 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 8096 0 1 2176
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85
timestamp 1676037725
transform 1 0 8924 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97
timestamp 1676037725
transform 1 0 10028 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_109
timestamp 1676037725
transform 1 0 11132 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_113
timestamp 1676037725
transform 1 0 11500 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_118
timestamp 1676037725
transform 1 0 11960 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_126
timestamp 1676037725
transform 1 0 12696 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_131
timestamp 1676037725
transform 1 0 13156 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_138
timestamp 1676037725
transform 1 0 13800 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_141 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 14076 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_147
timestamp 1676037725
transform 1 0 14628 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_151
timestamp 1676037725
transform 1 0 14996 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_158
timestamp 1676037725
transform 1 0 15640 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_166
timestamp 1676037725
transform 1 0 16376 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_169
timestamp 1676037725
transform 1 0 16652 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_174
timestamp 1676037725
transform 1 0 17112 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_188
timestamp 1676037725
transform 1 0 18400 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_197
timestamp 1676037725
transform 1 0 19228 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_202
timestamp 1676037725
transform 1 0 19688 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_210
timestamp 1676037725
transform 1 0 20424 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_216
timestamp 1676037725
transform 1 0 20976 0 1 2176
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_225
timestamp 1676037725
transform 1 0 21804 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_237
timestamp 1676037725
transform 1 0 22908 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_249
timestamp 1676037725
transform 1 0 24012 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_253
timestamp 1676037725
transform 1 0 24380 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_258
timestamp 1676037725
transform 1 0 24840 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_266
timestamp 1676037725
transform 1 0 25576 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_272
timestamp 1676037725
transform 1 0 26128 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_281
timestamp 1676037725
transform 1 0 26956 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_289
timestamp 1676037725
transform 1 0 27692 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_301
timestamp 1676037725
transform 1 0 28796 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_307
timestamp 1676037725
transform 1 0 29348 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_309
timestamp 1676037725
transform 1 0 29532 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_314
timestamp 1676037725
transform 1 0 29992 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_321
timestamp 1676037725
transform 1 0 30636 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_333
timestamp 1676037725
transform 1 0 31740 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_337
timestamp 1676037725
transform 1 0 32108 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_343
timestamp 1676037725
transform 1 0 32660 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_355
timestamp 1676037725
transform 1 0 33764 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_363
timestamp 1676037725
transform 1 0 34500 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_365
timestamp 1676037725
transform 1 0 34684 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_377
timestamp 1676037725
transform 1 0 35788 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_389
timestamp 1676037725
transform 1 0 36892 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_393
timestamp 1676037725
transform 1 0 37260 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_398
timestamp 1676037725
transform 1 0 37720 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_406
timestamp 1676037725
transform 1 0 38456 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_412
timestamp 1676037725
transform 1 0 39008 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_421
timestamp 1676037725
transform 1 0 39836 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_426
timestamp 1676037725
transform 1 0 40296 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_438
timestamp 1676037725
transform 1 0 41400 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_446
timestamp 1676037725
transform 1 0 42136 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_449
timestamp 1676037725
transform 1 0 42412 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_455
timestamp 1676037725
transform 1 0 42964 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_463
timestamp 1676037725
transform 1 0 43700 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_468
timestamp 1676037725
transform 1 0 44160 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_472
timestamp 1676037725
transform 1 0 44528 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_3
timestamp 1676037725
transform 1 0 1380 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_8
timestamp 1676037725
transform 1 0 1840 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_20
timestamp 1676037725
transform 1 0 2944 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_32
timestamp 1676037725
transform 1 0 4048 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_44
timestamp 1676037725
transform 1 0 5152 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_57
timestamp 1676037725
transform 1 0 6348 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_65
timestamp 1676037725
transform 1 0 7084 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_82
timestamp 1676037725
transform 1 0 8648 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_94
timestamp 1676037725
transform 1 0 9752 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_106
timestamp 1676037725
transform 1 0 10856 0 -1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_1_113
timestamp 1676037725
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_125
timestamp 1676037725
transform 1 0 12604 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_133
timestamp 1676037725
transform 1 0 13340 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_140
timestamp 1676037725
transform 1 0 13984 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_144
timestamp 1676037725
transform 1 0 14352 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_166
timestamp 1676037725
transform 1 0 16376 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_169
timestamp 1676037725
transform 1 0 16652 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_175
timestamp 1676037725
transform 1 0 17204 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_179
timestamp 1676037725
transform 1 0 17572 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_204
timestamp 1676037725
transform 1 0 19872 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_211
timestamp 1676037725
transform 1 0 20516 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_223
timestamp 1676037725
transform 1 0 21620 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_225
timestamp 1676037725
transform 1 0 21804 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_253
timestamp 1676037725
transform 1 0 24380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_265
timestamp 1676037725
transform 1 0 25484 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_1_277
timestamp 1676037725
transform 1 0 26588 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_1_281
timestamp 1676037725
transform 1 0 26956 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_293
timestamp 1676037725
transform 1 0 28060 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_305
timestamp 1676037725
transform 1 0 29164 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_317
timestamp 1676037725
transform 1 0 30268 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_329
timestamp 1676037725
transform 1 0 31372 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_335
timestamp 1676037725
transform 1 0 31924 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_337
timestamp 1676037725
transform 1 0 32108 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_349
timestamp 1676037725
transform 1 0 33212 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_357
timestamp 1676037725
transform 1 0 33948 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_1_376
timestamp 1676037725
transform 1 0 35696 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_388
timestamp 1676037725
transform 1 0 36800 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_393
timestamp 1676037725
transform 1 0 37260 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_405
timestamp 1676037725
transform 1 0 38364 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_417
timestamp 1676037725
transform 1 0 39468 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_429
timestamp 1676037725
transform 1 0 40572 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_441
timestamp 1676037725
transform 1 0 41676 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_447
timestamp 1676037725
transform 1 0 42228 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_449
timestamp 1676037725
transform 1 0 42412 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_461
timestamp 1676037725
transform 1 0 43516 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_467
timestamp 1676037725
transform 1 0 44068 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_471
timestamp 1676037725
transform 1 0 44436 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_3
timestamp 1676037725
transform 1 0 1380 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_8
timestamp 1676037725
transform 1 0 1840 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_20
timestamp 1676037725
transform 1 0 2944 0 1 3264
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_2_29
timestamp 1676037725
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_41
timestamp 1676037725
transform 1 0 4876 0 1 3264
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_2_65
timestamp 1676037725
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_77
timestamp 1676037725
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 1676037725
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_85
timestamp 1676037725
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_97
timestamp 1676037725
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_109
timestamp 1676037725
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_121
timestamp 1676037725
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_2_133
timestamp 1676037725
transform 1 0 13340 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_138
timestamp 1676037725
transform 1 0 13800 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_141
timestamp 1676037725
transform 1 0 14076 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_145
timestamp 1676037725
transform 1 0 14444 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_149
timestamp 1676037725
transform 1 0 14812 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_156
timestamp 1676037725
transform 1 0 15456 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_181
timestamp 1676037725
transform 1 0 17756 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_188
timestamp 1676037725
transform 1 0 18400 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_197
timestamp 1676037725
transform 1 0 19228 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_2_202
timestamp 1676037725
transform 1 0 19688 0 1 3264
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_2_213
timestamp 1676037725
transform 1 0 20700 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_225
timestamp 1676037725
transform 1 0 21804 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_237
timestamp 1676037725
transform 1 0 22908 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_245
timestamp 1676037725
transform 1 0 23644 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_250
timestamp 1676037725
transform 1 0 24104 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_2_253
timestamp 1676037725
transform 1 0 24380 0 1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_2_260
timestamp 1676037725
transform 1 0 25024 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_272
timestamp 1676037725
transform 1 0 26128 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_278
timestamp 1676037725
transform 1 0 26680 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_282
timestamp 1676037725
transform 1 0 27048 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_294
timestamp 1676037725
transform 1 0 28152 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_2_306
timestamp 1676037725
transform 1 0 29256 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_309
timestamp 1676037725
transform 1 0 29532 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_318
timestamp 1676037725
transform 1 0 30360 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_330
timestamp 1676037725
transform 1 0 31464 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_342
timestamp 1676037725
transform 1 0 32568 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_354
timestamp 1676037725
transform 1 0 33672 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_362
timestamp 1676037725
transform 1 0 34408 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_365
timestamp 1676037725
transform 1 0 34684 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_377
timestamp 1676037725
transform 1 0 35788 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_389
timestamp 1676037725
transform 1 0 36892 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_401
timestamp 1676037725
transform 1 0 37996 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_413
timestamp 1676037725
transform 1 0 39100 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_419
timestamp 1676037725
transform 1 0 39652 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_421
timestamp 1676037725
transform 1 0 39836 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_433
timestamp 1676037725
transform 1 0 40940 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_445
timestamp 1676037725
transform 1 0 42044 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_457
timestamp 1676037725
transform 1 0 43148 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_2_465
timestamp 1676037725
transform 1 0 43884 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_471
timestamp 1676037725
transform 1 0 44436 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3
timestamp 1676037725
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_15
timestamp 1676037725
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_27
timestamp 1676037725
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_39
timestamp 1676037725
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_51
timestamp 1676037725
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 1676037725
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_57
timestamp 1676037725
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_69
timestamp 1676037725
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_81
timestamp 1676037725
transform 1 0 8556 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_87
timestamp 1676037725
transform 1 0 9108 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_92
timestamp 1676037725
transform 1 0 9568 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_104
timestamp 1676037725
transform 1 0 10672 0 -1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_3_113
timestamp 1676037725
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_3_125
timestamp 1676037725
transform 1 0 12604 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_129
timestamp 1676037725
transform 1 0 12972 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_144
timestamp 1676037725
transform 1 0 14352 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_156
timestamp 1676037725
transform 1 0 15456 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_162
timestamp 1676037725
transform 1 0 16008 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_166
timestamp 1676037725
transform 1 0 16376 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_169
timestamp 1676037725
transform 1 0 16652 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_176
timestamp 1676037725
transform 1 0 17296 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_183
timestamp 1676037725
transform 1 0 17940 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_187
timestamp 1676037725
transform 1 0 18308 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_192
timestamp 1676037725
transform 1 0 18768 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_199
timestamp 1676037725
transform 1 0 19412 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_3_210
timestamp 1676037725
transform 1 0 20424 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_218
timestamp 1676037725
transform 1 0 21160 0 -1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_3_225
timestamp 1676037725
transform 1 0 21804 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_237
timestamp 1676037725
transform 1 0 22908 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_3_265
timestamp 1676037725
transform 1 0 25484 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_272
timestamp 1676037725
transform 1 0 26128 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_281
timestamp 1676037725
transform 1 0 26956 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_3_287
timestamp 1676037725
transform 1 0 27508 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_295
timestamp 1676037725
transform 1 0 28244 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_299
timestamp 1676037725
transform 1 0 28612 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_3_330
timestamp 1676037725
transform 1 0 31464 0 -1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_3_337
timestamp 1676037725
transform 1 0 32108 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_349
timestamp 1676037725
transform 1 0 33212 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_361
timestamp 1676037725
transform 1 0 34316 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_373
timestamp 1676037725
transform 1 0 35420 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_385
timestamp 1676037725
transform 1 0 36524 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_391
timestamp 1676037725
transform 1 0 37076 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_393
timestamp 1676037725
transform 1 0 37260 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_405
timestamp 1676037725
transform 1 0 38364 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_417
timestamp 1676037725
transform 1 0 39468 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_429
timestamp 1676037725
transform 1 0 40572 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_441
timestamp 1676037725
transform 1 0 41676 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_447
timestamp 1676037725
transform 1 0 42228 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_449
timestamp 1676037725
transform 1 0 42412 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_461
timestamp 1676037725
transform 1 0 43516 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3
timestamp 1676037725
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_15
timestamp 1676037725
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1676037725
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_29
timestamp 1676037725
transform 1 0 3772 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_37
timestamp 1676037725
transform 1 0 4508 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_43
timestamp 1676037725
transform 1 0 5060 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_55
timestamp 1676037725
transform 1 0 6164 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_67
timestamp 1676037725
transform 1 0 7268 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_79
timestamp 1676037725
transform 1 0 8372 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 1676037725
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_85
timestamp 1676037725
transform 1 0 8924 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_4_97
timestamp 1676037725
transform 1 0 10028 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_4_104
timestamp 1676037725
transform 1 0 10672 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_136
timestamp 1676037725
transform 1 0 13616 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_141
timestamp 1676037725
transform 1 0 14076 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_147
timestamp 1676037725
transform 1 0 14628 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_4_154
timestamp 1676037725
transform 1 0 15272 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_166
timestamp 1676037725
transform 1 0 16376 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_194
timestamp 1676037725
transform 1 0 18952 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_197
timestamp 1676037725
transform 1 0 19228 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_219
timestamp 1676037725
transform 1 0 21252 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_4_226
timestamp 1676037725
transform 1 0 21896 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_238
timestamp 1676037725
transform 1 0 23000 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_4_250
timestamp 1676037725
transform 1 0 24104 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_253
timestamp 1676037725
transform 1 0 24380 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_261
timestamp 1676037725
transform 1 0 25116 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_265
timestamp 1676037725
transform 1 0 25484 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_286
timestamp 1676037725
transform 1 0 27416 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_298
timestamp 1676037725
transform 1 0 28520 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_306
timestamp 1676037725
transform 1 0 29256 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_309
timestamp 1676037725
transform 1 0 29532 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_314
timestamp 1676037725
transform 1 0 29992 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_4_321
timestamp 1676037725
transform 1 0 30636 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_333
timestamp 1676037725
transform 1 0 31740 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_345
timestamp 1676037725
transform 1 0 32844 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_357
timestamp 1676037725
transform 1 0 33948 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_363
timestamp 1676037725
transform 1 0 34500 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_365
timestamp 1676037725
transform 1 0 34684 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_370
timestamp 1676037725
transform 1 0 35144 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_382
timestamp 1676037725
transform 1 0 36248 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_4_392
timestamp 1676037725
transform 1 0 37168 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_398
timestamp 1676037725
transform 1 0 37720 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_406
timestamp 1676037725
transform 1 0 38456 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_4_418
timestamp 1676037725
transform 1 0 39560 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_421
timestamp 1676037725
transform 1 0 39836 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_433
timestamp 1676037725
transform 1 0 40940 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_445
timestamp 1676037725
transform 1 0 42044 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_457
timestamp 1676037725
transform 1 0 43148 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_469
timestamp 1676037725
transform 1 0 44252 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_3
timestamp 1676037725
transform 1 0 1380 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_15
timestamp 1676037725
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_27
timestamp 1676037725
transform 1 0 3588 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_40
timestamp 1676037725
transform 1 0 4784 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_49
timestamp 1676037725
transform 1 0 5612 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1676037725
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_5_57
timestamp 1676037725
transform 1 0 6348 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_5_83
timestamp 1676037725
transform 1 0 8740 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_107
timestamp 1676037725
transform 1 0 10948 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1676037725
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_5_113
timestamp 1676037725
transform 1 0 11500 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_119
timestamp 1676037725
transform 1 0 12052 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_123
timestamp 1676037725
transform 1 0 12420 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_131
timestamp 1676037725
transform 1 0 13156 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_155
timestamp 1676037725
transform 1 0 15364 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_163
timestamp 1676037725
transform 1 0 16100 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 1676037725
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_5_169
timestamp 1676037725
transform 1 0 16652 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_177
timestamp 1676037725
transform 1 0 17388 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_188
timestamp 1676037725
transform 1 0 18400 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_197
timestamp 1676037725
transform 1 0 19228 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_5_208
timestamp 1676037725
transform 1 0 20240 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_215
timestamp 1676037725
transform 1 0 20884 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_222
timestamp 1676037725
transform 1 0 21528 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_5_225
timestamp 1676037725
transform 1 0 21804 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_233
timestamp 1676037725
transform 1 0 22540 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_237
timestamp 1676037725
transform 1 0 22908 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_244
timestamp 1676037725
transform 1 0 23552 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_255
timestamp 1676037725
transform 1 0 24564 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_264
timestamp 1676037725
transform 1 0 25392 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_271
timestamp 1676037725
transform 1 0 26036 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_278
timestamp 1676037725
transform 1 0 26680 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_281
timestamp 1676037725
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_313
timestamp 1676037725
transform 1 0 29900 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_325
timestamp 1676037725
transform 1 0 31004 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_5_333
timestamp 1676037725
transform 1 0 31740 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_5_337
timestamp 1676037725
transform 1 0 32108 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_345
timestamp 1676037725
transform 1 0 32844 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_349
timestamp 1676037725
transform 1 0 33212 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_369
timestamp 1676037725
transform 1 0 35052 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_5_389
timestamp 1676037725
transform 1 0 36892 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_393
timestamp 1676037725
transform 1 0 37260 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_5_398
timestamp 1676037725
transform 1 0 37720 0 -1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_5_412
timestamp 1676037725
transform 1 0 39008 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_424
timestamp 1676037725
transform 1 0 40112 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_5_436
timestamp 1676037725
transform 1 0 41216 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_443
timestamp 1676037725
transform 1 0 41860 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_447
timestamp 1676037725
transform 1 0 42228 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_449
timestamp 1676037725
transform 1 0 42412 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_469
timestamp 1676037725
transform 1 0 44252 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_3
timestamp 1676037725
transform 1 0 1380 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_6_8
timestamp 1676037725
transform 1 0 1840 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_16
timestamp 1676037725
transform 1 0 2576 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_6_21
timestamp 1676037725
transform 1 0 3036 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1676037725
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_29
timestamp 1676037725
transform 1 0 3772 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_47
timestamp 1676037725
transform 1 0 5428 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_6_57
timestamp 1676037725
transform 1 0 6348 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_6_65
timestamp 1676037725
transform 1 0 7084 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_71
timestamp 1676037725
transform 1 0 7636 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_75
timestamp 1676037725
transform 1 0 8004 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_82
timestamp 1676037725
transform 1 0 8648 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_85
timestamp 1676037725
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_97
timestamp 1676037725
transform 1 0 10028 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_121
timestamp 1676037725
transform 1 0 12236 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_6_128
timestamp 1676037725
transform 1 0 12880 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_6_138
timestamp 1676037725
transform 1 0 13800 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_141
timestamp 1676037725
transform 1 0 14076 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_159
timestamp 1676037725
transform 1 0 15732 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_6_166
timestamp 1676037725
transform 1 0 16376 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_6_178
timestamp 1676037725
transform 1 0 17480 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_183
timestamp 1676037725
transform 1 0 17940 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_194
timestamp 1676037725
transform 1 0 18952 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_197
timestamp 1676037725
transform 1 0 19228 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_206
timestamp 1676037725
transform 1 0 20056 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_216
timestamp 1676037725
transform 1 0 20976 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_6_223
timestamp 1676037725
transform 1 0 21620 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_6_234
timestamp 1676037725
transform 1 0 22632 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_241
timestamp 1676037725
transform 1 0 23276 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_250
timestamp 1676037725
transform 1 0 24104 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_253
timestamp 1676037725
transform 1 0 24380 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_6_261
timestamp 1676037725
transform 1 0 25116 0 1 5440
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_6_273
timestamp 1676037725
transform 1 0 26220 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_6_285
timestamp 1676037725
transform 1 0 27324 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_6_290
timestamp 1676037725
transform 1 0 27784 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_298
timestamp 1676037725
transform 1 0 28520 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_303
timestamp 1676037725
transform 1 0 28980 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_307
timestamp 1676037725
transform 1 0 29348 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_309
timestamp 1676037725
transform 1 0 29532 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_315
timestamp 1676037725
transform 1 0 30084 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_323
timestamp 1676037725
transform 1 0 30820 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_6_347
timestamp 1676037725
transform 1 0 33028 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_355
timestamp 1676037725
transform 1 0 33764 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_362
timestamp 1676037725
transform 1 0 34408 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_365
timestamp 1676037725
transform 1 0 34684 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_383
timestamp 1676037725
transform 1 0 36340 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_6_392
timestamp 1676037725
transform 1 0 37168 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_400
timestamp 1676037725
transform 1 0 37904 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_409
timestamp 1676037725
transform 1 0 38732 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_6_417
timestamp 1676037725
transform 1 0 39468 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_6_421
timestamp 1676037725
transform 1 0 39836 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_429
timestamp 1676037725
transform 1 0 40572 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_447
timestamp 1676037725
transform 1 0 42228 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_459
timestamp 1676037725
transform 1 0 43332 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_6_471
timestamp 1676037725
transform 1 0 44436 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_7_3
timestamp 1676037725
transform 1 0 1380 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_9
timestamp 1676037725
transform 1 0 1932 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_26
timestamp 1676037725
transform 1 0 3496 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_30
timestamp 1676037725
transform 1 0 3864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_47
timestamp 1676037725
transform 1 0 5428 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_54
timestamp 1676037725
transform 1 0 6072 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_57
timestamp 1676037725
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_69
timestamp 1676037725
transform 1 0 7452 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_77
timestamp 1676037725
transform 1 0 8188 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_81
timestamp 1676037725
transform 1 0 8556 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_91
timestamp 1676037725
transform 1 0 9476 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_101
timestamp 1676037725
transform 1 0 10396 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_108
timestamp 1676037725
transform 1 0 11040 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_7_113
timestamp 1676037725
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_125
timestamp 1676037725
transform 1 0 12604 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_149
timestamp 1676037725
transform 1 0 14812 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_7_160
timestamp 1676037725
transform 1 0 15824 0 -1 6528
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_7_169
timestamp 1676037725
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_189
timestamp 1676037725
transform 1 0 18492 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_201
timestamp 1676037725
transform 1 0 19596 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_215
timestamp 1676037725
transform 1 0 20884 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_223
timestamp 1676037725
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_225
timestamp 1676037725
transform 1 0 21804 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_237
timestamp 1676037725
transform 1 0 22908 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_242
timestamp 1676037725
transform 1 0 23368 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_251
timestamp 1676037725
transform 1 0 24196 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_275
timestamp 1676037725
transform 1 0 26404 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_279
timestamp 1676037725
transform 1 0 26772 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_281
timestamp 1676037725
transform 1 0 26956 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_7_286
timestamp 1676037725
transform 1 0 27416 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_7_294
timestamp 1676037725
transform 1 0 28152 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_7_300
timestamp 1676037725
transform 1 0 28704 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_307
timestamp 1676037725
transform 1 0 29348 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_315
timestamp 1676037725
transform 1 0 30084 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_322
timestamp 1676037725
transform 1 0 30728 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_7_329
timestamp 1676037725
transform 1 0 31372 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_335
timestamp 1676037725
transform 1 0 31924 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_337
timestamp 1676037725
transform 1 0 32108 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_352
timestamp 1676037725
transform 1 0 33488 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_363
timestamp 1676037725
transform 1 0 34500 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_7_378
timestamp 1676037725
transform 1 0 35880 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_388
timestamp 1676037725
transform 1 0 36800 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_393
timestamp 1676037725
transform 1 0 37260 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_7_398
timestamp 1676037725
transform 1 0 37720 0 -1 6528
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_7_415
timestamp 1676037725
transform 1 0 39284 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_427
timestamp 1676037725
transform 1 0 40388 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_433
timestamp 1676037725
transform 1 0 40940 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_7_441
timestamp 1676037725
transform 1 0 41676 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_447
timestamp 1676037725
transform 1 0 42228 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_449
timestamp 1676037725
transform 1 0 42412 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_454
timestamp 1676037725
transform 1 0 42872 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_466
timestamp 1676037725
transform 1 0 43976 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_472
timestamp 1676037725
transform 1 0 44528 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_8_3
timestamp 1676037725
transform 1 0 1380 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_9
timestamp 1676037725
transform 1 0 1932 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_26
timestamp 1676037725
transform 1 0 3496 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_29
timestamp 1676037725
transform 1 0 3772 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_8_47
timestamp 1676037725
transform 1 0 5428 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_55
timestamp 1676037725
transform 1 0 6164 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_60
timestamp 1676037725
transform 1 0 6624 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_72
timestamp 1676037725
transform 1 0 7728 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_8_82
timestamp 1676037725
transform 1 0 8648 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_85
timestamp 1676037725
transform 1 0 8924 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_8_107
timestamp 1676037725
transform 1 0 10948 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_8_118
timestamp 1676037725
transform 1 0 11960 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_125
timestamp 1676037725
transform 1 0 12604 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_138
timestamp 1676037725
transform 1 0 13800 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_141
timestamp 1676037725
transform 1 0 14076 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_8_146
timestamp 1676037725
transform 1 0 14536 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_8_170
timestamp 1676037725
transform 1 0 16744 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_183
timestamp 1676037725
transform 1 0 17940 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_194
timestamp 1676037725
transform 1 0 18952 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_8_197
timestamp 1676037725
transform 1 0 19228 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_205
timestamp 1676037725
transform 1 0 19964 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_216
timestamp 1676037725
transform 1 0 20976 0 1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_8_228
timestamp 1676037725
transform 1 0 22080 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_240
timestamp 1676037725
transform 1 0 23184 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_250
timestamp 1676037725
transform 1 0 24104 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_253
timestamp 1676037725
transform 1 0 24380 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_8_262
timestamp 1676037725
transform 1 0 25208 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_8_271
timestamp 1676037725
transform 1 0 26036 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_8_280
timestamp 1676037725
transform 1 0 26864 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_300
timestamp 1676037725
transform 1 0 28704 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_309
timestamp 1676037725
transform 1 0 29532 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_327
timestamp 1676037725
transform 1 0 31188 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_339
timestamp 1676037725
transform 1 0 32292 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_346
timestamp 1676037725
transform 1 0 32936 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_8_354
timestamp 1676037725
transform 1 0 33672 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_362
timestamp 1676037725
transform 1 0 34408 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_8_365
timestamp 1676037725
transform 1 0 34684 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_371
timestamp 1676037725
transform 1 0 35236 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_379
timestamp 1676037725
transform 1 0 35972 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_390
timestamp 1676037725
transform 1 0 36984 0 1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_8_397
timestamp 1676037725
transform 1 0 37628 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_409
timestamp 1676037725
transform 1 0 38732 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_8_418
timestamp 1676037725
transform 1 0 39560 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_421
timestamp 1676037725
transform 1 0 39836 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_8_431
timestamp 1676037725
transform 1 0 40756 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_8_453
timestamp 1676037725
transform 1 0 42780 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_464
timestamp 1676037725
transform 1 0 43792 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_472
timestamp 1676037725
transform 1 0 44528 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_9_3
timestamp 1676037725
transform 1 0 1380 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_9_12
timestamp 1676037725
transform 1 0 2208 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_36
timestamp 1676037725
transform 1 0 4416 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_49
timestamp 1676037725
transform 1 0 5612 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 1676037725
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_57
timestamp 1676037725
transform 1 0 6348 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_9_68
timestamp 1676037725
transform 1 0 7360 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_88
timestamp 1676037725
transform 1 0 9200 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_92
timestamp 1676037725
transform 1 0 9568 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_97
timestamp 1676037725
transform 1 0 10028 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_105
timestamp 1676037725
transform 1 0 10764 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_110
timestamp 1676037725
transform 1 0 11224 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_113
timestamp 1676037725
transform 1 0 11500 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_118
timestamp 1676037725
transform 1 0 11960 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_125
timestamp 1676037725
transform 1 0 12604 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_131
timestamp 1676037725
transform 1 0 13156 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_148
timestamp 1676037725
transform 1 0 14720 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_161
timestamp 1676037725
transform 1 0 15916 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_167
timestamp 1676037725
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_9_169
timestamp 1676037725
transform 1 0 16652 0 -1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_9_178
timestamp 1676037725
transform 1 0 17480 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_190
timestamp 1676037725
transform 1 0 18584 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_202
timestamp 1676037725
transform 1 0 19688 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_220
timestamp 1676037725
transform 1 0 21344 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_9_225
timestamp 1676037725
transform 1 0 21804 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_237
timestamp 1676037725
transform 1 0 22908 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_255
timestamp 1676037725
transform 1 0 24564 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_267
timestamp 1676037725
transform 1 0 25668 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_276
timestamp 1676037725
transform 1 0 26496 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_281
timestamp 1676037725
transform 1 0 26956 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_306
timestamp 1676037725
transform 1 0 29256 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_313
timestamp 1676037725
transform 1 0 29900 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_320
timestamp 1676037725
transform 1 0 30544 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_324
timestamp 1676037725
transform 1 0 30912 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_9_333
timestamp 1676037725
transform 1 0 31740 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_337
timestamp 1676037725
transform 1 0 32108 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_347
timestamp 1676037725
transform 1 0 33028 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_356
timestamp 1676037725
transform 1 0 33856 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_360
timestamp 1676037725
transform 1 0 34224 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_364
timestamp 1676037725
transform 1 0 34592 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_374
timestamp 1676037725
transform 1 0 35512 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_378
timestamp 1676037725
transform 1 0 35880 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_387
timestamp 1676037725
transform 1 0 36708 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_391
timestamp 1676037725
transform 1 0 37076 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_393
timestamp 1676037725
transform 1 0 37260 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_398
timestamp 1676037725
transform 1 0 37720 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_402
timestamp 1676037725
transform 1 0 38088 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_9_408
timestamp 1676037725
transform 1 0 38640 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_9_422
timestamp 1676037725
transform 1 0 39928 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_434
timestamp 1676037725
transform 1 0 41032 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_441
timestamp 1676037725
transform 1 0 41676 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_447
timestamp 1676037725
transform 1 0 42228 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_449
timestamp 1676037725
transform 1 0 42412 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_454
timestamp 1676037725
transform 1 0 42872 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_466
timestamp 1676037725
transform 1 0 43976 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_472
timestamp 1676037725
transform 1 0 44528 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_3
timestamp 1676037725
transform 1 0 1380 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_10_8
timestamp 1676037725
transform 1 0 1840 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_16
timestamp 1676037725
transform 1 0 2576 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_26
timestamp 1676037725
transform 1 0 3496 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_29
timestamp 1676037725
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_41
timestamp 1676037725
transform 1 0 4876 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_10_65
timestamp 1676037725
transform 1 0 7084 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_82
timestamp 1676037725
transform 1 0 8648 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_10_85
timestamp 1676037725
transform 1 0 8924 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_10_96
timestamp 1676037725
transform 1 0 9936 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_10_119
timestamp 1676037725
transform 1 0 12052 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_10_132
timestamp 1676037725
transform 1 0 13248 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_10_141
timestamp 1676037725
transform 1 0 14076 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_10_165
timestamp 1676037725
transform 1 0 16284 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_10_172
timestamp 1676037725
transform 1 0 16928 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_180
timestamp 1676037725
transform 1 0 17664 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_10_190
timestamp 1676037725
transform 1 0 18584 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_10_197
timestamp 1676037725
transform 1 0 19228 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_203
timestamp 1676037725
transform 1 0 19780 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_220
timestamp 1676037725
transform 1 0 21344 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_10_227
timestamp 1676037725
transform 1 0 21988 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_10_236
timestamp 1676037725
transform 1 0 22816 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_240
timestamp 1676037725
transform 1 0 23184 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_244
timestamp 1676037725
transform 1 0 23552 0 1 7616
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_10_253
timestamp 1676037725
transform 1 0 24380 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_265
timestamp 1676037725
transform 1 0 25484 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_269
timestamp 1676037725
transform 1 0 25852 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_294
timestamp 1676037725
transform 1 0 28152 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_298
timestamp 1676037725
transform 1 0 28520 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_303
timestamp 1676037725
transform 1 0 28980 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_307
timestamp 1676037725
transform 1 0 29348 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_309
timestamp 1676037725
transform 1 0 29532 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_10_333
timestamp 1676037725
transform 1 0 31740 0 1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_10_342
timestamp 1676037725
transform 1 0 32568 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_354
timestamp 1676037725
transform 1 0 33672 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_362
timestamp 1676037725
transform 1 0 34408 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_365
timestamp 1676037725
transform 1 0 34684 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_369
timestamp 1676037725
transform 1 0 35052 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_386
timestamp 1676037725
transform 1 0 36616 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_395
timestamp 1676037725
transform 1 0 37444 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_10_402
timestamp 1676037725
transform 1 0 38088 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_418
timestamp 1676037725
transform 1 0 39560 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_10_421
timestamp 1676037725
transform 1 0 39836 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_427
timestamp 1676037725
transform 1 0 40388 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_444
timestamp 1676037725
transform 1 0 41952 0 1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_10_451
timestamp 1676037725
transform 1 0 42596 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_463
timestamp 1676037725
transform 1 0 43700 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_467
timestamp 1676037725
transform 1 0 44068 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_471
timestamp 1676037725
transform 1 0 44436 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_3
timestamp 1676037725
transform 1 0 1380 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_11_27
timestamp 1676037725
transform 1 0 3588 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_47
timestamp 1676037725
transform 1 0 5428 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 1676037725
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_57
timestamp 1676037725
transform 1 0 6348 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_75
timestamp 1676037725
transform 1 0 8004 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_95
timestamp 1676037725
transform 1 0 9844 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_99
timestamp 1676037725
transform 1 0 10212 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_103
timestamp 1676037725
transform 1 0 10580 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_110
timestamp 1676037725
transform 1 0 11224 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_113
timestamp 1676037725
transform 1 0 11500 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_135
timestamp 1676037725
transform 1 0 13524 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_147
timestamp 1676037725
transform 1 0 14628 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_151
timestamp 1676037725
transform 1 0 14996 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_11_161
timestamp 1676037725
transform 1 0 15916 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_167
timestamp 1676037725
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_11_169
timestamp 1676037725
transform 1 0 16652 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_11_191
timestamp 1676037725
transform 1 0 18676 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_11_208
timestamp 1676037725
transform 1 0 20240 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_11_221
timestamp 1676037725
transform 1 0 21436 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_225
timestamp 1676037725
transform 1 0 21804 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_11_246
timestamp 1676037725
transform 1 0 23736 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_258
timestamp 1676037725
transform 1 0 24840 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_11_266
timestamp 1676037725
transform 1 0 25576 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_11_278
timestamp 1676037725
transform 1 0 26680 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_281
timestamp 1676037725
transform 1 0 26956 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_295
timestamp 1676037725
transform 1 0 28244 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_11_319
timestamp 1676037725
transform 1 0 30452 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_11_330
timestamp 1676037725
transform 1 0 31464 0 -1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_11_337
timestamp 1676037725
transform 1 0 32108 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_349
timestamp 1676037725
transform 1 0 33212 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_11_361
timestamp 1676037725
transform 1 0 34316 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_369
timestamp 1676037725
transform 1 0 35052 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_378
timestamp 1676037725
transform 1 0 35880 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_387
timestamp 1676037725
transform 1 0 36708 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_391
timestamp 1676037725
transform 1 0 37076 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_393
timestamp 1676037725
transform 1 0 37260 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_405
timestamp 1676037725
transform 1 0 38364 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_11_410
timestamp 1676037725
transform 1 0 38824 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_11_424
timestamp 1676037725
transform 1 0 40112 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_436
timestamp 1676037725
transform 1 0 41216 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_11_445
timestamp 1676037725
transform 1 0 42044 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_449
timestamp 1676037725
transform 1 0 42412 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_458
timestamp 1676037725
transform 1 0 43240 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_466
timestamp 1676037725
transform 1 0 43976 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_471
timestamp 1676037725
transform 1 0 44436 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3
timestamp 1676037725
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_15
timestamp 1676037725
transform 1 0 2484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 1676037725
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_29
timestamp 1676037725
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_41
timestamp 1676037725
transform 1 0 4876 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_65
timestamp 1676037725
transform 1 0 7084 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_78
timestamp 1676037725
transform 1 0 8280 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_12_85
timestamp 1676037725
transform 1 0 8924 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_93
timestamp 1676037725
transform 1 0 9660 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_97
timestamp 1676037725
transform 1 0 10028 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_121
timestamp 1676037725
transform 1 0 12236 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_134
timestamp 1676037725
transform 1 0 13432 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_12_141
timestamp 1676037725
transform 1 0 14076 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_146
timestamp 1676037725
transform 1 0 14536 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_158
timestamp 1676037725
transform 1 0 15640 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_12_180
timestamp 1676037725
transform 1 0 17664 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_12_187
timestamp 1676037725
transform 1 0 18308 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_195
timestamp 1676037725
transform 1 0 19044 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_12_197
timestamp 1676037725
transform 1 0 19228 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_12_203
timestamp 1676037725
transform 1 0 19780 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_210
timestamp 1676037725
transform 1 0 20424 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_234
timestamp 1676037725
transform 1 0 22632 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_12_244
timestamp 1676037725
transform 1 0 23552 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_253
timestamp 1676037725
transform 1 0 24380 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_275
timestamp 1676037725
transform 1 0 26404 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_285
timestamp 1676037725
transform 1 0 27324 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_289
timestamp 1676037725
transform 1 0 27692 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_306
timestamp 1676037725
transform 1 0 29256 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_12_309
timestamp 1676037725
transform 1 0 29532 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_315
timestamp 1676037725
transform 1 0 30084 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_325
timestamp 1676037725
transform 1 0 31004 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_329
timestamp 1676037725
transform 1 0 31372 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_337
timestamp 1676037725
transform 1 0 32108 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_349
timestamp 1676037725
transform 1 0 33212 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_12_362
timestamp 1676037725
transform 1 0 34408 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_365
timestamp 1676037725
transform 1 0 34684 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_369
timestamp 1676037725
transform 1 0 35052 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_378
timestamp 1676037725
transform 1 0 35880 0 1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_12_386
timestamp 1676037725
transform 1 0 36616 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_398
timestamp 1676037725
transform 1 0 37720 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_406
timestamp 1676037725
transform 1 0 38456 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_410
timestamp 1676037725
transform 1 0 38824 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_418
timestamp 1676037725
transform 1 0 39560 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_421
timestamp 1676037725
transform 1 0 39836 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_426
timestamp 1676037725
transform 1 0 40296 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_446
timestamp 1676037725
transform 1 0 42136 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_466
timestamp 1676037725
transform 1 0 43976 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_472
timestamp 1676037725
transform 1 0 44528 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3
timestamp 1676037725
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_31
timestamp 1676037725
transform 1 0 3956 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_43
timestamp 1676037725
transform 1 0 5060 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_54
timestamp 1676037725
transform 1 0 6072 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_57
timestamp 1676037725
transform 1 0 6348 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_13_75
timestamp 1676037725
transform 1 0 8004 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_87
timestamp 1676037725
transform 1 0 9108 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_99
timestamp 1676037725
transform 1 0 10212 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_110
timestamp 1676037725
transform 1 0 11224 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_113
timestamp 1676037725
transform 1 0 11500 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_135
timestamp 1676037725
transform 1 0 13524 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_142
timestamp 1676037725
transform 1 0 14168 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_166
timestamp 1676037725
transform 1 0 16376 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_169
timestamp 1676037725
transform 1 0 16652 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_13_187
timestamp 1676037725
transform 1 0 18308 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_13_195
timestamp 1676037725
transform 1 0 19044 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_201
timestamp 1676037725
transform 1 0 19596 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_209
timestamp 1676037725
transform 1 0 20332 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_222
timestamp 1676037725
transform 1 0 21528 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_225
timestamp 1676037725
transform 1 0 21804 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_249
timestamp 1676037725
transform 1 0 24012 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_13_257
timestamp 1676037725
transform 1 0 24748 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_263
timestamp 1676037725
transform 1 0 25300 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_278
timestamp 1676037725
transform 1 0 26680 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_281
timestamp 1676037725
transform 1 0 26956 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_286
timestamp 1676037725
transform 1 0 27416 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_293
timestamp 1676037725
transform 1 0 28060 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_302
timestamp 1676037725
transform 1 0 28888 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_322
timestamp 1676037725
transform 1 0 30728 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_329
timestamp 1676037725
transform 1 0 31372 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_335
timestamp 1676037725
transform 1 0 31924 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_13_337
timestamp 1676037725
transform 1 0 32108 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_343
timestamp 1676037725
transform 1 0 32660 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_347
timestamp 1676037725
transform 1 0 33028 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_13_352
timestamp 1676037725
transform 1 0 33488 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_13_364
timestamp 1676037725
transform 1 0 34592 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_368
timestamp 1676037725
transform 1 0 34960 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_380
timestamp 1676037725
transform 1 0 36064 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_390
timestamp 1676037725
transform 1 0 36984 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_393
timestamp 1676037725
transform 1 0 37260 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_13_398
timestamp 1676037725
transform 1 0 37720 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_410
timestamp 1676037725
transform 1 0 38824 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_13_420
timestamp 1676037725
transform 1 0 39744 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_432
timestamp 1676037725
transform 1 0 40848 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_13_445
timestamp 1676037725
transform 1 0 42044 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_449
timestamp 1676037725
transform 1 0 42412 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_13_454
timestamp 1676037725
transform 1 0 42872 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_466
timestamp 1676037725
transform 1 0 43976 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_472
timestamp 1676037725
transform 1 0 44528 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_3
timestamp 1676037725
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_15
timestamp 1676037725
transform 1 0 2484 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_22
timestamp 1676037725
transform 1 0 3128 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_14_29
timestamp 1676037725
transform 1 0 3772 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_40
timestamp 1676037725
transform 1 0 4784 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_52
timestamp 1676037725
transform 1 0 5888 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_58
timestamp 1676037725
transform 1 0 6440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_75
timestamp 1676037725
transform 1 0 8004 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1676037725
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_85
timestamp 1676037725
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_14_97
timestamp 1676037725
transform 1 0 10028 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_14_121
timestamp 1676037725
transform 1 0 12236 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_14_132
timestamp 1676037725
transform 1 0 13248 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_141
timestamp 1676037725
transform 1 0 14076 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_146
timestamp 1676037725
transform 1 0 14536 0 1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_14_153
timestamp 1676037725
transform 1 0 15180 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_165
timestamp 1676037725
transform 1 0 16284 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_170
timestamp 1676037725
transform 1 0 16744 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_183
timestamp 1676037725
transform 1 0 17940 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_192
timestamp 1676037725
transform 1 0 18768 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_197
timestamp 1676037725
transform 1 0 19228 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_207
timestamp 1676037725
transform 1 0 20148 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_232
timestamp 1676037725
transform 1 0 22448 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_245
timestamp 1676037725
transform 1 0 23644 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_251
timestamp 1676037725
transform 1 0 24196 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_253
timestamp 1676037725
transform 1 0 24380 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_265
timestamp 1676037725
transform 1 0 25484 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_271
timestamp 1676037725
transform 1 0 26036 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_275
timestamp 1676037725
transform 1 0 26404 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_282
timestamp 1676037725
transform 1 0 27048 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_286
timestamp 1676037725
transform 1 0 27416 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_291
timestamp 1676037725
transform 1 0 27876 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_298
timestamp 1676037725
transform 1 0 28520 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_306
timestamp 1676037725
transform 1 0 29256 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_309
timestamp 1676037725
transform 1 0 29532 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_314
timestamp 1676037725
transform 1 0 29992 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_318
timestamp 1676037725
transform 1 0 30360 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_322
timestamp 1676037725
transform 1 0 30728 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_334
timestamp 1676037725
transform 1 0 31832 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_342
timestamp 1676037725
transform 1 0 32568 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_350
timestamp 1676037725
transform 1 0 33304 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_355
timestamp 1676037725
transform 1 0 33764 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_362
timestamp 1676037725
transform 1 0 34408 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_365
timestamp 1676037725
transform 1 0 34684 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_387
timestamp 1676037725
transform 1 0 36708 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_398
timestamp 1676037725
transform 1 0 37720 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_406
timestamp 1676037725
transform 1 0 38456 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_412
timestamp 1676037725
transform 1 0 39008 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_418
timestamp 1676037725
transform 1 0 39560 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_421
timestamp 1676037725
transform 1 0 39836 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_429
timestamp 1676037725
transform 1 0 40572 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_449
timestamp 1676037725
transform 1 0 42412 0 1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_14_457
timestamp 1676037725
transform 1 0 43148 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_469
timestamp 1676037725
transform 1 0 44252 0 1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_3
timestamp 1676037725
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_15_15
timestamp 1676037725
transform 1 0 2484 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_20
timestamp 1676037725
transform 1 0 2944 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_15_40
timestamp 1676037725
transform 1 0 4784 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_15_51
timestamp 1676037725
transform 1 0 5796 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_55
timestamp 1676037725
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_57
timestamp 1676037725
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_69
timestamp 1676037725
transform 1 0 7452 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_15_93
timestamp 1676037725
transform 1 0 9660 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_110
timestamp 1676037725
transform 1 0 11224 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_113
timestamp 1676037725
transform 1 0 11500 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_125
timestamp 1676037725
transform 1 0 12604 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_15_149
timestamp 1676037725
transform 1 0 14812 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_15_158
timestamp 1676037725
transform 1 0 15640 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_166
timestamp 1676037725
transform 1 0 16376 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_169
timestamp 1676037725
transform 1 0 16652 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_15_191
timestamp 1676037725
transform 1 0 18676 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_15_203
timestamp 1676037725
transform 1 0 19780 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_209
timestamp 1676037725
transform 1 0 20332 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_222
timestamp 1676037725
transform 1 0 21528 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_225
timestamp 1676037725
transform 1 0 21804 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_229
timestamp 1676037725
transform 1 0 22172 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_246
timestamp 1676037725
transform 1 0 23736 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_258
timestamp 1676037725
transform 1 0 24840 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_15_270
timestamp 1676037725
transform 1 0 25944 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_278
timestamp 1676037725
transform 1 0 26680 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_281
timestamp 1676037725
transform 1 0 26956 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_306
timestamp 1676037725
transform 1 0 29256 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_15_330
timestamp 1676037725
transform 1 0 31464 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_15_337
timestamp 1676037725
transform 1 0 32108 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_361
timestamp 1676037725
transform 1 0 34316 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_15_385
timestamp 1676037725
transform 1 0 36524 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_391
timestamp 1676037725
transform 1 0 37076 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_393
timestamp 1676037725
transform 1 0 37260 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_15_398
timestamp 1676037725
transform 1 0 37720 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_410
timestamp 1676037725
transform 1 0 38824 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_417
timestamp 1676037725
transform 1 0 39468 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_426
timestamp 1676037725
transform 1 0 40296 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_446
timestamp 1676037725
transform 1 0 42136 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_449
timestamp 1676037725
transform 1 0 42412 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_15_454
timestamp 1676037725
transform 1 0 42872 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_466
timestamp 1676037725
transform 1 0 43976 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_472
timestamp 1676037725
transform 1 0 44528 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_16_3
timestamp 1676037725
transform 1 0 1380 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_9
timestamp 1676037725
transform 1 0 1932 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_26
timestamp 1676037725
transform 1 0 3496 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_29
timestamp 1676037725
transform 1 0 3772 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_40
timestamp 1676037725
transform 1 0 4784 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_48
timestamp 1676037725
transform 1 0 5520 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_68
timestamp 1676037725
transform 1 0 7360 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_75
timestamp 1676037725
transform 1 0 8004 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1676037725
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_85
timestamp 1676037725
transform 1 0 8924 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_93
timestamp 1676037725
transform 1 0 9660 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_97
timestamp 1676037725
transform 1 0 10028 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_16_114
timestamp 1676037725
transform 1 0 11592 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_127
timestamp 1676037725
transform 1 0 12788 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_133
timestamp 1676037725
transform 1 0 13340 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_16_137
timestamp 1676037725
transform 1 0 13708 0 1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_16_141
timestamp 1676037725
transform 1 0 14076 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_153
timestamp 1676037725
transform 1 0 15180 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_16_165
timestamp 1676037725
transform 1 0 16284 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_172
timestamp 1676037725
transform 1 0 16928 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_16_181
timestamp 1676037725
transform 1 0 17756 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_16_193
timestamp 1676037725
transform 1 0 18860 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_16_197
timestamp 1676037725
transform 1 0 19228 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_205
timestamp 1676037725
transform 1 0 19964 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_209
timestamp 1676037725
transform 1 0 20332 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_233
timestamp 1676037725
transform 1 0 22540 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_239
timestamp 1676037725
transform 1 0 23092 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_244
timestamp 1676037725
transform 1 0 23552 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_16_253
timestamp 1676037725
transform 1 0 24380 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_16_281
timestamp 1676037725
transform 1 0 26956 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_290
timestamp 1676037725
transform 1 0 27784 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_296
timestamp 1676037725
transform 1 0 28336 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_16_305
timestamp 1676037725
transform 1 0 29164 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_16_309
timestamp 1676037725
transform 1 0 29532 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_16_320
timestamp 1676037725
transform 1 0 30544 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_344
timestamp 1676037725
transform 1 0 32752 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_351
timestamp 1676037725
transform 1 0 33396 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_358
timestamp 1676037725
transform 1 0 34040 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_16_365
timestamp 1676037725
transform 1 0 34684 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_373
timestamp 1676037725
transform 1 0 35420 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_382
timestamp 1676037725
transform 1 0 36248 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_390
timestamp 1676037725
transform 1 0 36984 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_399
timestamp 1676037725
transform 1 0 37812 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_406
timestamp 1676037725
transform 1 0 38456 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_413
timestamp 1676037725
transform 1 0 39100 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_419
timestamp 1676037725
transform 1 0 39652 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_421
timestamp 1676037725
transform 1 0 39836 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_16_428
timestamp 1676037725
transform 1 0 40480 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_436
timestamp 1676037725
transform 1 0 41216 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_447
timestamp 1676037725
transform 1 0 42228 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_459
timestamp 1676037725
transform 1 0 43332 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_467
timestamp 1676037725
transform 1 0 44068 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_471
timestamp 1676037725
transform 1 0 44436 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_17_3
timestamp 1676037725
transform 1 0 1380 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_17_25
timestamp 1676037725
transform 1 0 3404 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_45
timestamp 1676037725
transform 1 0 5244 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_54
timestamp 1676037725
transform 1 0 6072 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_57
timestamp 1676037725
transform 1 0 6348 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_68
timestamp 1676037725
transform 1 0 7360 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_80
timestamp 1676037725
transform 1 0 8464 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_92
timestamp 1676037725
transform 1 0 9568 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_17_100
timestamp 1676037725
transform 1 0 10304 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_110
timestamp 1676037725
transform 1 0 11224 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_113
timestamp 1676037725
transform 1 0 11500 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_117
timestamp 1676037725
transform 1 0 11868 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_127
timestamp 1676037725
transform 1 0 12788 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_17_140
timestamp 1676037725
transform 1 0 13984 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_152
timestamp 1676037725
transform 1 0 15088 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_164
timestamp 1676037725
transform 1 0 16192 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_169
timestamp 1676037725
transform 1 0 16652 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_180
timestamp 1676037725
transform 1 0 17664 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_187
timestamp 1676037725
transform 1 0 18308 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_17_194
timestamp 1676037725
transform 1 0 18952 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_206
timestamp 1676037725
transform 1 0 20056 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_212
timestamp 1676037725
transform 1 0 20608 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_222
timestamp 1676037725
transform 1 0 21528 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_225
timestamp 1676037725
transform 1 0 21804 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_236
timestamp 1676037725
transform 1 0 22816 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_248
timestamp 1676037725
transform 1 0 23920 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_260
timestamp 1676037725
transform 1 0 25024 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_17_272
timestamp 1676037725
transform 1 0 26128 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_278
timestamp 1676037725
transform 1 0 26680 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_281
timestamp 1676037725
transform 1 0 26956 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_285
timestamp 1676037725
transform 1 0 27324 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_291
timestamp 1676037725
transform 1 0 27876 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_17_299
timestamp 1676037725
transform 1 0 28612 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_17_306
timestamp 1676037725
transform 1 0 29256 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_17_317
timestamp 1676037725
transform 1 0 30268 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_17_328
timestamp 1676037725
transform 1 0 31280 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_337
timestamp 1676037725
transform 1 0 32108 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_344
timestamp 1676037725
transform 1 0 32752 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_356
timestamp 1676037725
transform 1 0 33856 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_368
timestamp 1676037725
transform 1 0 34960 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_374
timestamp 1676037725
transform 1 0 35512 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_378
timestamp 1676037725
transform 1 0 35880 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_387
timestamp 1676037725
transform 1 0 36708 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_391
timestamp 1676037725
transform 1 0 37076 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_393
timestamp 1676037725
transform 1 0 37260 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_17_398
timestamp 1676037725
transform 1 0 37720 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_404
timestamp 1676037725
transform 1 0 38272 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_421
timestamp 1676037725
transform 1 0 39836 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_429
timestamp 1676037725
transform 1 0 40572 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_446
timestamp 1676037725
transform 1 0 42136 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_449
timestamp 1676037725
transform 1 0 42412 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_461
timestamp 1676037725
transform 1 0 43516 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_3
timestamp 1676037725
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_15
timestamp 1676037725
transform 1 0 2484 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_26
timestamp 1676037725
transform 1 0 3496 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_29
timestamp 1676037725
transform 1 0 3772 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_34
timestamp 1676037725
transform 1 0 4232 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_44
timestamp 1676037725
transform 1 0 5152 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_64
timestamp 1676037725
transform 1 0 6992 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_70
timestamp 1676037725
transform 1 0 7544 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_74
timestamp 1676037725
transform 1 0 7912 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_82
timestamp 1676037725
transform 1 0 8648 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_18_85
timestamp 1676037725
transform 1 0 8924 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_91
timestamp 1676037725
transform 1 0 9476 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_99
timestamp 1676037725
transform 1 0 10212 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_111
timestamp 1676037725
transform 1 0 11316 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_123
timestamp 1676037725
transform 1 0 12420 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_138
timestamp 1676037725
transform 1 0 13800 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_141
timestamp 1676037725
transform 1 0 14076 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_151
timestamp 1676037725
transform 1 0 14996 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_163
timestamp 1676037725
transform 1 0 16100 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_167
timestamp 1676037725
transform 1 0 16468 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_18_175
timestamp 1676037725
transform 1 0 17204 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_181
timestamp 1676037725
transform 1 0 17756 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_185
timestamp 1676037725
transform 1 0 18124 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_18_193
timestamp 1676037725
transform 1 0 18860 0 1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_18_197
timestamp 1676037725
transform 1 0 19228 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_209
timestamp 1676037725
transform 1 0 20332 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_213
timestamp 1676037725
transform 1 0 20700 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_217
timestamp 1676037725
transform 1 0 21068 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_225
timestamp 1676037725
transform 1 0 21804 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_232
timestamp 1676037725
transform 1 0 22448 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_240
timestamp 1676037725
transform 1 0 23184 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_250
timestamp 1676037725
transform 1 0 24104 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_253
timestamp 1676037725
transform 1 0 24380 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_258
timestamp 1676037725
transform 1 0 24840 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_265
timestamp 1676037725
transform 1 0 25484 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_271
timestamp 1676037725
transform 1 0 26036 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_292
timestamp 1676037725
transform 1 0 27968 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_302
timestamp 1676037725
transform 1 0 28888 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_18_309
timestamp 1676037725
transform 1 0 29532 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_18_323
timestamp 1676037725
transform 1 0 30820 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_347
timestamp 1676037725
transform 1 0 33028 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_355
timestamp 1676037725
transform 1 0 33764 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_362
timestamp 1676037725
transform 1 0 34408 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_365
timestamp 1676037725
transform 1 0 34684 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_387
timestamp 1676037725
transform 1 0 36708 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_391
timestamp 1676037725
transform 1 0 37076 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_412
timestamp 1676037725
transform 1 0 39008 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_421
timestamp 1676037725
transform 1 0 39836 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_426
timestamp 1676037725
transform 1 0 40296 0 1 11968
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_18_450
timestamp 1676037725
transform 1 0 42504 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_462
timestamp 1676037725
transform 1 0 43608 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_18_470
timestamp 1676037725
transform 1 0 44344 0 1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_19_3
timestamp 1676037725
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_15
timestamp 1676037725
transform 1 0 2484 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_21
timestamp 1676037725
transform 1 0 3036 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_27
timestamp 1676037725
transform 1 0 3588 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_19_38
timestamp 1676037725
transform 1 0 4600 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_45
timestamp 1676037725
transform 1 0 5244 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_54
timestamp 1676037725
transform 1 0 6072 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_57
timestamp 1676037725
transform 1 0 6348 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_64
timestamp 1676037725
transform 1 0 6992 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_19_71
timestamp 1676037725
transform 1 0 7636 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_83
timestamp 1676037725
transform 1 0 8740 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_89
timestamp 1676037725
transform 1 0 9292 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_93
timestamp 1676037725
transform 1 0 9660 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_19_105
timestamp 1676037725
transform 1 0 10764 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_110
timestamp 1676037725
transform 1 0 11224 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_113
timestamp 1676037725
transform 1 0 11500 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_125
timestamp 1676037725
transform 1 0 12604 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_145
timestamp 1676037725
transform 1 0 14444 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_19_152
timestamp 1676037725
transform 1 0 15088 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_164
timestamp 1676037725
transform 1 0 16192 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_169
timestamp 1676037725
transform 1 0 16652 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_177
timestamp 1676037725
transform 1 0 17388 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_194
timestamp 1676037725
transform 1 0 18952 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_214
timestamp 1676037725
transform 1 0 20792 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_222
timestamp 1676037725
transform 1 0 21528 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_225
timestamp 1676037725
transform 1 0 21804 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_19_236
timestamp 1676037725
transform 1 0 22816 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_19_260
timestamp 1676037725
transform 1 0 25024 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_19_272
timestamp 1676037725
transform 1 0 26128 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_278
timestamp 1676037725
transform 1 0 26680 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_281
timestamp 1676037725
transform 1 0 26956 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_19_286
timestamp 1676037725
transform 1 0 27416 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_19_312
timestamp 1676037725
transform 1 0 29808 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_319
timestamp 1676037725
transform 1 0 30452 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_323
timestamp 1676037725
transform 1 0 30820 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_19_333
timestamp 1676037725
transform 1 0 31740 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_337
timestamp 1676037725
transform 1 0 32108 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_344
timestamp 1676037725
transform 1 0 32752 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_19_351
timestamp 1676037725
transform 1 0 33396 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_363
timestamp 1676037725
transform 1 0 34500 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_19_375
timestamp 1676037725
transform 1 0 35604 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_382
timestamp 1676037725
transform 1 0 36248 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_19_389
timestamp 1676037725
transform 1 0 36892 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_393
timestamp 1676037725
transform 1 0 37260 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_19_398
timestamp 1676037725
transform 1 0 37720 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_404
timestamp 1676037725
transform 1 0 38272 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_428
timestamp 1676037725
transform 1 0 40480 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_19_435
timestamp 1676037725
transform 1 0 41124 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_19_447
timestamp 1676037725
transform 1 0 42228 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_449
timestamp 1676037725
transform 1 0 42412 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_461
timestamp 1676037725
transform 1 0 43516 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_467
timestamp 1676037725
transform 1 0 44068 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_471
timestamp 1676037725
transform 1 0 44436 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_3
timestamp 1676037725
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_15
timestamp 1676037725
transform 1 0 2484 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_26
timestamp 1676037725
transform 1 0 3496 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_29
timestamp 1676037725
transform 1 0 3772 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_47
timestamp 1676037725
transform 1 0 5428 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_56
timestamp 1676037725
transform 1 0 6256 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_67
timestamp 1676037725
transform 1 0 7268 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_76
timestamp 1676037725
transform 1 0 8096 0 1 13056
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_20_85
timestamp 1676037725
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_97
timestamp 1676037725
transform 1 0 10028 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_109
timestamp 1676037725
transform 1 0 11132 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_113
timestamp 1676037725
transform 1 0 11500 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_120
timestamp 1676037725
transform 1 0 12144 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_130
timestamp 1676037725
transform 1 0 13064 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_134
timestamp 1676037725
transform 1 0 13432 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_138
timestamp 1676037725
transform 1 0 13800 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_141
timestamp 1676037725
transform 1 0 14076 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_148
timestamp 1676037725
transform 1 0 14720 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_20_157
timestamp 1676037725
transform 1 0 15548 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_169
timestamp 1676037725
transform 1 0 16652 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_177
timestamp 1676037725
transform 1 0 17388 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_194
timestamp 1676037725
transform 1 0 18952 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_197
timestamp 1676037725
transform 1 0 19228 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_208
timestamp 1676037725
transform 1 0 20240 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_20_220
timestamp 1676037725
transform 1 0 21344 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_20_232
timestamp 1676037725
transform 1 0 22448 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_240
timestamp 1676037725
transform 1 0 23184 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_250
timestamp 1676037725
transform 1 0 24104 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_253
timestamp 1676037725
transform 1 0 24380 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_20_273
timestamp 1676037725
transform 1 0 26220 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_285
timestamp 1676037725
transform 1 0 27324 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_295
timestamp 1676037725
transform 1 0 28244 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_302
timestamp 1676037725
transform 1 0 28888 0 1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_20_309
timestamp 1676037725
transform 1 0 29532 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_321
timestamp 1676037725
transform 1 0 30636 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_338
timestamp 1676037725
transform 1 0 32200 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_20_345
timestamp 1676037725
transform 1 0 32844 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_357
timestamp 1676037725
transform 1 0 33948 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_363
timestamp 1676037725
transform 1 0 34500 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_365
timestamp 1676037725
transform 1 0 34684 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_377
timestamp 1676037725
transform 1 0 35788 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_20_399
timestamp 1676037725
transform 1 0 37812 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_20_406
timestamp 1676037725
transform 1 0 38456 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_20_418
timestamp 1676037725
transform 1 0 39560 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_421
timestamp 1676037725
transform 1 0 39836 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_433
timestamp 1676037725
transform 1 0 40940 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_445
timestamp 1676037725
transform 1 0 42044 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_457
timestamp 1676037725
transform 1 0 43148 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_469
timestamp 1676037725
transform 1 0 44252 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_3
timestamp 1676037725
transform 1 0 1380 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_8
timestamp 1676037725
transform 1 0 1840 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_16
timestamp 1676037725
transform 1 0 2576 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_21_35
timestamp 1676037725
transform 1 0 4324 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_41
timestamp 1676037725
transform 1 0 4876 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_46
timestamp 1676037725
transform 1 0 5336 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_54
timestamp 1676037725
transform 1 0 6072 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_57
timestamp 1676037725
transform 1 0 6348 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_75
timestamp 1676037725
transform 1 0 8004 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_21_84
timestamp 1676037725
transform 1 0 8832 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_96
timestamp 1676037725
transform 1 0 9936 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_104
timestamp 1676037725
transform 1 0 10672 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_110
timestamp 1676037725
transform 1 0 11224 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_113
timestamp 1676037725
transform 1 0 11500 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_122
timestamp 1676037725
transform 1 0 12328 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_131
timestamp 1676037725
transform 1 0 13156 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_151
timestamp 1676037725
transform 1 0 14996 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_21_158
timestamp 1676037725
transform 1 0 15640 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_166
timestamp 1676037725
transform 1 0 16376 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_169
timestamp 1676037725
transform 1 0 16652 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_21_181
timestamp 1676037725
transform 1 0 17756 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_185
timestamp 1676037725
transform 1 0 18124 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_205
timestamp 1676037725
transform 1 0 19964 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_21_218
timestamp 1676037725
transform 1 0 21160 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_21_225
timestamp 1676037725
transform 1 0 21804 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_243
timestamp 1676037725
transform 1 0 23460 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_21_256
timestamp 1676037725
transform 1 0 24656 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_268
timestamp 1676037725
transform 1 0 25760 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_281
timestamp 1676037725
transform 1 0 26956 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_293
timestamp 1676037725
transform 1 0 28060 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_305
timestamp 1676037725
transform 1 0 29164 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_311
timestamp 1676037725
transform 1 0 29716 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_317
timestamp 1676037725
transform 1 0 30268 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_325
timestamp 1676037725
transform 1 0 31004 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_331
timestamp 1676037725
transform 1 0 31556 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_335
timestamp 1676037725
transform 1 0 31924 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_337
timestamp 1676037725
transform 1 0 32108 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_345
timestamp 1676037725
transform 1 0 32844 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_363
timestamp 1676037725
transform 1 0 34500 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_21_374
timestamp 1676037725
transform 1 0 35512 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_387
timestamp 1676037725
transform 1 0 36708 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_391
timestamp 1676037725
transform 1 0 37076 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_393
timestamp 1676037725
transform 1 0 37260 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_404
timestamp 1676037725
transform 1 0 38272 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_408
timestamp 1676037725
transform 1 0 38640 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_425
timestamp 1676037725
transform 1 0 40204 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_446
timestamp 1676037725
transform 1 0 42136 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_449
timestamp 1676037725
transform 1 0 42412 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_461
timestamp 1676037725
transform 1 0 43516 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_3
timestamp 1676037725
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_15
timestamp 1676037725
transform 1 0 2484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 1676037725
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_29
timestamp 1676037725
transform 1 0 3772 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_37
timestamp 1676037725
transform 1 0 4508 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_22_42
timestamp 1676037725
transform 1 0 4968 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_48
timestamp 1676037725
transform 1 0 5520 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_52
timestamp 1676037725
transform 1 0 5888 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_61
timestamp 1676037725
transform 1 0 6716 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_22_81
timestamp 1676037725
transform 1 0 8556 0 1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_22_85
timestamp 1676037725
transform 1 0 8924 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_97
timestamp 1676037725
transform 1 0 10028 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_105
timestamp 1676037725
transform 1 0 10764 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_109
timestamp 1676037725
transform 1 0 11132 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_129
timestamp 1676037725
transform 1 0 12972 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_136
timestamp 1676037725
transform 1 0 13616 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_141
timestamp 1676037725
transform 1 0 14076 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_22_146
timestamp 1676037725
transform 1 0 14536 0 1 14144
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_22_163
timestamp 1676037725
transform 1 0 16100 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_22_175
timestamp 1676037725
transform 1 0 17204 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_181
timestamp 1676037725
transform 1 0 17756 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_194
timestamp 1676037725
transform 1 0 18952 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_197
timestamp 1676037725
transform 1 0 19228 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_208
timestamp 1676037725
transform 1 0 20240 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_220
timestamp 1676037725
transform 1 0 21344 0 1 14144
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_22_229
timestamp 1676037725
transform 1 0 22172 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_22_250
timestamp 1676037725
transform 1 0 24104 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_22_253
timestamp 1676037725
transform 1 0 24380 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_259
timestamp 1676037725
transform 1 0 24932 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_269
timestamp 1676037725
transform 1 0 25852 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_282
timestamp 1676037725
transform 1 0 27048 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_306
timestamp 1676037725
transform 1 0 29256 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_309
timestamp 1676037725
transform 1 0 29532 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_22_316
timestamp 1676037725
transform 1 0 30176 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_324
timestamp 1676037725
transform 1 0 30912 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_341
timestamp 1676037725
transform 1 0 32476 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_22_362
timestamp 1676037725
transform 1 0 34408 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_365
timestamp 1676037725
transform 1 0 34684 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_383
timestamp 1676037725
transform 1 0 36340 0 1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_22_396
timestamp 1676037725
transform 1 0 37536 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_408
timestamp 1676037725
transform 1 0 38640 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_414
timestamp 1676037725
transform 1 0 39192 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_418
timestamp 1676037725
transform 1 0 39560 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_421
timestamp 1676037725
transform 1 0 39836 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_439
timestamp 1676037725
transform 1 0 41492 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_22_451
timestamp 1676037725
transform 1 0 42596 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_469
timestamp 1676037725
transform 1 0 44252 0 1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_23_3
timestamp 1676037725
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_15
timestamp 1676037725
transform 1 0 2484 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_27
timestamp 1676037725
transform 1 0 3588 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_39
timestamp 1676037725
transform 1 0 4692 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_51
timestamp 1676037725
transform 1 0 5796 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_55
timestamp 1676037725
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_57
timestamp 1676037725
transform 1 0 6348 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_62
timestamp 1676037725
transform 1 0 6808 0 -1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_23_69
timestamp 1676037725
transform 1 0 7452 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_81
timestamp 1676037725
transform 1 0 8556 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_93
timestamp 1676037725
transform 1 0 9660 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_105
timestamp 1676037725
transform 1 0 10764 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_111
timestamp 1676037725
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_113
timestamp 1676037725
transform 1 0 11500 0 -1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_23_133
timestamp 1676037725
transform 1 0 13340 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_145
timestamp 1676037725
transform 1 0 14444 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_149
timestamp 1676037725
transform 1 0 14812 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_166
timestamp 1676037725
transform 1 0 16376 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_169
timestamp 1676037725
transform 1 0 16652 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_173
timestamp 1676037725
transform 1 0 17020 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_190
timestamp 1676037725
transform 1 0 18584 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_210
timestamp 1676037725
transform 1 0 20424 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_23_217
timestamp 1676037725
transform 1 0 21068 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_223
timestamp 1676037725
transform 1 0 21620 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_225
timestamp 1676037725
transform 1 0 21804 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_23_237
timestamp 1676037725
transform 1 0 22908 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_254
timestamp 1676037725
transform 1 0 24472 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_23_274
timestamp 1676037725
transform 1 0 26312 0 -1 15232
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_23_281
timestamp 1676037725
transform 1 0 26956 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_293
timestamp 1676037725
transform 1 0 28060 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_297
timestamp 1676037725
transform 1 0 28428 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_23_314
timestamp 1676037725
transform 1 0 29992 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_23_323
timestamp 1676037725
transform 1 0 30820 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_23_330
timestamp 1676037725
transform 1 0 31464 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_23_337
timestamp 1676037725
transform 1 0 32108 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_23_348
timestamp 1676037725
transform 1 0 33120 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_356
timestamp 1676037725
transform 1 0 33856 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_360
timestamp 1676037725
transform 1 0 34224 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_380
timestamp 1676037725
transform 1 0 36064 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_387
timestamp 1676037725
transform 1 0 36708 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_391
timestamp 1676037725
transform 1 0 37076 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_393
timestamp 1676037725
transform 1 0 37260 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_405
timestamp 1676037725
transform 1 0 38364 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_417
timestamp 1676037725
transform 1 0 39468 0 -1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_23_426
timestamp 1676037725
transform 1 0 40296 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_438
timestamp 1676037725
transform 1 0 41400 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_446
timestamp 1676037725
transform 1 0 42136 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_23_449
timestamp 1676037725
transform 1 0 42412 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_461
timestamp 1676037725
transform 1 0 43516 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_3
timestamp 1676037725
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_15
timestamp 1676037725
transform 1 0 2484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1676037725
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_29
timestamp 1676037725
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_41
timestamp 1676037725
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_53
timestamp 1676037725
transform 1 0 5980 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_65
timestamp 1676037725
transform 1 0 7084 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_77
timestamp 1676037725
transform 1 0 8188 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_83
timestamp 1676037725
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_85
timestamp 1676037725
transform 1 0 8924 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_97
timestamp 1676037725
transform 1 0 10028 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_114
timestamp 1676037725
transform 1 0 11592 0 1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_24_126
timestamp 1676037725
transform 1 0 12696 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_24_138
timestamp 1676037725
transform 1 0 13800 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_141
timestamp 1676037725
transform 1 0 14076 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_153
timestamp 1676037725
transform 1 0 15180 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_165
timestamp 1676037725
transform 1 0 16284 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_24_177
timestamp 1676037725
transform 1 0 17388 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_184
timestamp 1676037725
transform 1 0 18032 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_24_197
timestamp 1676037725
transform 1 0 19228 0 1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_24_209
timestamp 1676037725
transform 1 0 20332 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_221
timestamp 1676037725
transform 1 0 21436 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_233
timestamp 1676037725
transform 1 0 22540 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_245
timestamp 1676037725
transform 1 0 23644 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_251
timestamp 1676037725
transform 1 0 24196 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_24_253
timestamp 1676037725
transform 1 0 24380 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_259
timestamp 1676037725
transform 1 0 24932 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_263
timestamp 1676037725
transform 1 0 25300 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_275
timestamp 1676037725
transform 1 0 26404 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_287
timestamp 1676037725
transform 1 0 27508 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_299
timestamp 1676037725
transform 1 0 28612 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_307
timestamp 1676037725
transform 1 0 29348 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_309
timestamp 1676037725
transform 1 0 29532 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_321
timestamp 1676037725
transform 1 0 30636 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_333
timestamp 1676037725
transform 1 0 31740 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_345
timestamp 1676037725
transform 1 0 32844 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_357
timestamp 1676037725
transform 1 0 33948 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_363
timestamp 1676037725
transform 1 0 34500 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_365
timestamp 1676037725
transform 1 0 34684 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_24_373
timestamp 1676037725
transform 1 0 35420 0 1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_24_385
timestamp 1676037725
transform 1 0 36524 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_397
timestamp 1676037725
transform 1 0 37628 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_409
timestamp 1676037725
transform 1 0 38732 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_24_417
timestamp 1676037725
transform 1 0 39468 0 1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_24_421
timestamp 1676037725
transform 1 0 39836 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_433
timestamp 1676037725
transform 1 0 40940 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_445
timestamp 1676037725
transform 1 0 42044 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_24_469
timestamp 1676037725
transform 1 0 44252 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_3
timestamp 1676037725
transform 1 0 1380 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_8
timestamp 1676037725
transform 1 0 1840 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_20
timestamp 1676037725
transform 1 0 2944 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_32
timestamp 1676037725
transform 1 0 4048 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_44
timestamp 1676037725
transform 1 0 5152 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_57
timestamp 1676037725
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_69
timestamp 1676037725
transform 1 0 7452 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_81
timestamp 1676037725
transform 1 0 8556 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_93
timestamp 1676037725
transform 1 0 9660 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_105
timestamp 1676037725
transform 1 0 10764 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_111
timestamp 1676037725
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_113
timestamp 1676037725
transform 1 0 11500 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_125
timestamp 1676037725
transform 1 0 12604 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_137
timestamp 1676037725
transform 1 0 13708 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_149
timestamp 1676037725
transform 1 0 14812 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_161
timestamp 1676037725
transform 1 0 15916 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_167
timestamp 1676037725
transform 1 0 16468 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_169
timestamp 1676037725
transform 1 0 16652 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_181
timestamp 1676037725
transform 1 0 17756 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_193
timestamp 1676037725
transform 1 0 18860 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_205
timestamp 1676037725
transform 1 0 19964 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_217
timestamp 1676037725
transform 1 0 21068 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_223
timestamp 1676037725
transform 1 0 21620 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_225
timestamp 1676037725
transform 1 0 21804 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_237
timestamp 1676037725
transform 1 0 22908 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_249
timestamp 1676037725
transform 1 0 24012 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_261
timestamp 1676037725
transform 1 0 25116 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_273
timestamp 1676037725
transform 1 0 26220 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_279
timestamp 1676037725
transform 1 0 26772 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_281
timestamp 1676037725
transform 1 0 26956 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_293
timestamp 1676037725
transform 1 0 28060 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_305
timestamp 1676037725
transform 1 0 29164 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_317
timestamp 1676037725
transform 1 0 30268 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_329
timestamp 1676037725
transform 1 0 31372 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_335
timestamp 1676037725
transform 1 0 31924 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_337
timestamp 1676037725
transform 1 0 32108 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_349
timestamp 1676037725
transform 1 0 33212 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_361
timestamp 1676037725
transform 1 0 34316 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_25_373
timestamp 1676037725
transform 1 0 35420 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_25_384
timestamp 1676037725
transform 1 0 36432 0 -1 16320
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_25_393
timestamp 1676037725
transform 1 0 37260 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_405
timestamp 1676037725
transform 1 0 38364 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_417
timestamp 1676037725
transform 1 0 39468 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_429
timestamp 1676037725
transform 1 0 40572 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_441
timestamp 1676037725
transform 1 0 41676 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_447
timestamp 1676037725
transform 1 0 42228 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_449
timestamp 1676037725
transform 1 0 42412 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_461
timestamp 1676037725
transform 1 0 43516 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_467
timestamp 1676037725
transform 1 0 44068 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_471
timestamp 1676037725
transform 1 0 44436 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_3
timestamp 1676037725
transform 1 0 1380 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_9
timestamp 1676037725
transform 1 0 1932 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_21
timestamp 1676037725
transform 1 0 3036 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 1676037725
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_29
timestamp 1676037725
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_41
timestamp 1676037725
transform 1 0 4876 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_53
timestamp 1676037725
transform 1 0 5980 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_61
timestamp 1676037725
transform 1 0 6716 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_79
timestamp 1676037725
transform 1 0 8372 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_83
timestamp 1676037725
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_85
timestamp 1676037725
transform 1 0 8924 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_97
timestamp 1676037725
transform 1 0 10028 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_109
timestamp 1676037725
transform 1 0 11132 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_121
timestamp 1676037725
transform 1 0 12236 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_133
timestamp 1676037725
transform 1 0 13340 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_139
timestamp 1676037725
transform 1 0 13892 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_141
timestamp 1676037725
transform 1 0 14076 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_153
timestamp 1676037725
transform 1 0 15180 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_165
timestamp 1676037725
transform 1 0 16284 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_177
timestamp 1676037725
transform 1 0 17388 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_189
timestamp 1676037725
transform 1 0 18492 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_195
timestamp 1676037725
transform 1 0 19044 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_197
timestamp 1676037725
transform 1 0 19228 0 1 16320
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_26_221
timestamp 1676037725
transform 1 0 21436 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_233
timestamp 1676037725
transform 1 0 22540 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_245
timestamp 1676037725
transform 1 0 23644 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_251
timestamp 1676037725
transform 1 0 24196 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_253
timestamp 1676037725
transform 1 0 24380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_265
timestamp 1676037725
transform 1 0 25484 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_277
timestamp 1676037725
transform 1 0 26588 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_289
timestamp 1676037725
transform 1 0 27692 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_301
timestamp 1676037725
transform 1 0 28796 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_307
timestamp 1676037725
transform 1 0 29348 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_309
timestamp 1676037725
transform 1 0 29532 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_321
timestamp 1676037725
transform 1 0 30636 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_333
timestamp 1676037725
transform 1 0 31740 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_345
timestamp 1676037725
transform 1 0 32844 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_357
timestamp 1676037725
transform 1 0 33948 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_363
timestamp 1676037725
transform 1 0 34500 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_365
timestamp 1676037725
transform 1 0 34684 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_377
timestamp 1676037725
transform 1 0 35788 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_389
timestamp 1676037725
transform 1 0 36892 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_401
timestamp 1676037725
transform 1 0 37996 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_413
timestamp 1676037725
transform 1 0 39100 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_419
timestamp 1676037725
transform 1 0 39652 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_421
timestamp 1676037725
transform 1 0 39836 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_433
timestamp 1676037725
transform 1 0 40940 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_445
timestamp 1676037725
transform 1 0 42044 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_457
timestamp 1676037725
transform 1 0 43148 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_26_465
timestamp 1676037725
transform 1 0 43884 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_471
timestamp 1676037725
transform 1 0 44436 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_3
timestamp 1676037725
transform 1 0 1380 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_9
timestamp 1676037725
transform 1 0 1932 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_17
timestamp 1676037725
transform 1 0 2668 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_21
timestamp 1676037725
transform 1 0 3036 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_26
timestamp 1676037725
transform 1 0 3496 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_27_29
timestamp 1676037725
transform 1 0 3772 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_37
timestamp 1676037725
transform 1 0 4508 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_48
timestamp 1676037725
transform 1 0 5520 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_57
timestamp 1676037725
transform 1 0 6348 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_27_62
timestamp 1676037725
transform 1 0 6808 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_70
timestamp 1676037725
transform 1 0 7544 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_27_76
timestamp 1676037725
transform 1 0 8096 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_27_85
timestamp 1676037725
transform 1 0 8924 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_93
timestamp 1676037725
transform 1 0 9660 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_97
timestamp 1676037725
transform 1 0 10028 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_27_109
timestamp 1676037725
transform 1 0 11132 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_113
timestamp 1676037725
transform 1 0 11500 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_27_119
timestamp 1676037725
transform 1 0 12052 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_127
timestamp 1676037725
transform 1 0 12788 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_27_132
timestamp 1676037725
transform 1 0 13248 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_141
timestamp 1676037725
transform 1 0 14076 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_27_146
timestamp 1676037725
transform 1 0 14536 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_158
timestamp 1676037725
transform 1 0 15640 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_166
timestamp 1676037725
transform 1 0 16376 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_169
timestamp 1676037725
transform 1 0 16652 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_27_175
timestamp 1676037725
transform 1 0 17204 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_187
timestamp 1676037725
transform 1 0 18308 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_195
timestamp 1676037725
transform 1 0 19044 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_197
timestamp 1676037725
transform 1 0 19228 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_27_202
timestamp 1676037725
transform 1 0 19688 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_214
timestamp 1676037725
transform 1 0 20792 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_222
timestamp 1676037725
transform 1 0 21528 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_27_225
timestamp 1676037725
transform 1 0 21804 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_233
timestamp 1676037725
transform 1 0 22540 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_237
timestamp 1676037725
transform 1 0 22908 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_27_249
timestamp 1676037725
transform 1 0 24012 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_253
timestamp 1676037725
transform 1 0 24380 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_27_258
timestamp 1676037725
transform 1 0 24840 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_266
timestamp 1676037725
transform 1 0 25576 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_27_272
timestamp 1676037725
transform 1 0 26128 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_27_281
timestamp 1676037725
transform 1 0 26956 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_289
timestamp 1676037725
transform 1 0 27692 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_293
timestamp 1676037725
transform 1 0 28060 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_27_305
timestamp 1676037725
transform 1 0 29164 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_309
timestamp 1676037725
transform 1 0 29532 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_27_314
timestamp 1676037725
transform 1 0 29992 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_322
timestamp 1676037725
transform 1 0 30728 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_27_328
timestamp 1676037725
transform 1 0 31280 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_337
timestamp 1676037725
transform 1 0 32108 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_27_349
timestamp 1676037725
transform 1 0 33212 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_27_361
timestamp 1676037725
transform 1 0 34316 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_365
timestamp 1676037725
transform 1 0 34684 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_370
timestamp 1676037725
transform 1 0 35144 0 -1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_27_377
timestamp 1676037725
transform 1 0 35788 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_27_389
timestamp 1676037725
transform 1 0 36892 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_393
timestamp 1676037725
transform 1 0 37260 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_27_398
timestamp 1676037725
transform 1 0 37720 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_406
timestamp 1676037725
transform 1 0 38456 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_27_413
timestamp 1676037725
transform 1 0 39100 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_419
timestamp 1676037725
transform 1 0 39652 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_421
timestamp 1676037725
transform 1 0 39836 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_433
timestamp 1676037725
transform 1 0 40940 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_27_445
timestamp 1676037725
transform 1 0 42044 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_449
timestamp 1676037725
transform 1 0 42412 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_454
timestamp 1676037725
transform 1 0 42872 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_461
timestamp 1676037725
transform 1 0 43516 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_468
timestamp 1676037725
transform 1 0 44160 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_472
timestamp 1676037725
transform 1 0 44528 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1676037725
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1676037725
transform -1 0 44896 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1676037725
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1676037725
transform -1 0 44896 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1676037725
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1676037725
transform -1 0 44896 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1676037725
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1676037725
transform -1 0 44896 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1676037725
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1676037725
transform -1 0 44896 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1676037725
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1676037725
transform -1 0 44896 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1676037725
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1676037725
transform -1 0 44896 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1676037725
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1676037725
transform -1 0 44896 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1676037725
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1676037725
transform -1 0 44896 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1676037725
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1676037725
transform -1 0 44896 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1676037725
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1676037725
transform -1 0 44896 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1676037725
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1676037725
transform -1 0 44896 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1676037725
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1676037725
transform -1 0 44896 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1676037725
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1676037725
transform -1 0 44896 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1676037725
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1676037725
transform -1 0 44896 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1676037725
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1676037725
transform -1 0 44896 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1676037725
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1676037725
transform -1 0 44896 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1676037725
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1676037725
transform -1 0 44896 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1676037725
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1676037725
transform -1 0 44896 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1676037725
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1676037725
transform -1 0 44896 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1676037725
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1676037725
transform -1 0 44896 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1676037725
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1676037725
transform -1 0 44896 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1676037725
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1676037725
transform -1 0 44896 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1676037725
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1676037725
transform -1 0 44896 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1676037725
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1676037725
transform -1 0 44896 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1676037725
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1676037725
transform -1 0 44896 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1676037725
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1676037725
transform -1 0 44896 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1676037725
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1676037725
transform -1 0 44896 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_56 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_57
timestamp 1676037725
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_58
timestamp 1676037725
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_59
timestamp 1676037725
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_60
timestamp 1676037725
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_61
timestamp 1676037725
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_62
timestamp 1676037725
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_63
timestamp 1676037725
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_64
timestamp 1676037725
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_65
timestamp 1676037725
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_66
timestamp 1676037725
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_67
timestamp 1676037725
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_68
timestamp 1676037725
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_69
timestamp 1676037725
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_70
timestamp 1676037725
transform 1 0 39744 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_71
timestamp 1676037725
transform 1 0 42320 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_72
timestamp 1676037725
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_73
timestamp 1676037725
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_74
timestamp 1676037725
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_75
timestamp 1676037725
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_76
timestamp 1676037725
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_77
timestamp 1676037725
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_78
timestamp 1676037725
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_79
timestamp 1676037725
transform 1 0 42320 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_80
timestamp 1676037725
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_81
timestamp 1676037725
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_82
timestamp 1676037725
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_83
timestamp 1676037725
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_84
timestamp 1676037725
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_85
timestamp 1676037725
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_86
timestamp 1676037725
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_87
timestamp 1676037725
transform 1 0 39744 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_88
timestamp 1676037725
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_89
timestamp 1676037725
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_90
timestamp 1676037725
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_91
timestamp 1676037725
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_92
timestamp 1676037725
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_93
timestamp 1676037725
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94
timestamp 1676037725
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1676037725
transform 1 0 42320 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 1676037725
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 1676037725
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 1676037725
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 1676037725
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 1676037725
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_101
timestamp 1676037725
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102
timestamp 1676037725
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 1676037725
transform 1 0 39744 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 1676037725
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 1676037725
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 1676037725
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 1676037725
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 1676037725
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1676037725
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1676037725
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1676037725
transform 1 0 42320 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1676037725
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1676037725
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1676037725
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1676037725
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 1676037725
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1676037725
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1676037725
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1676037725
transform 1 0 39744 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1676037725
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_121
timestamp 1676037725
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_122
timestamp 1676037725
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_123
timestamp 1676037725
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_124
timestamp 1676037725
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_125
timestamp 1676037725
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_126
timestamp 1676037725
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_127
timestamp 1676037725
transform 1 0 42320 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_128
timestamp 1676037725
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_129
timestamp 1676037725
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130
timestamp 1676037725
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1676037725
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1676037725
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1676037725
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1676037725
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1676037725
transform 1 0 39744 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1676037725
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1676037725
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1676037725
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1676037725
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1676037725
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1676037725
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1676037725
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1676037725
transform 1 0 42320 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1676037725
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1676037725
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1676037725
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1676037725
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1676037725
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1676037725
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1676037725
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1676037725
transform 1 0 39744 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1676037725
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1676037725
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1676037725
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1676037725
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1676037725
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1676037725
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1676037725
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1676037725
transform 1 0 42320 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1676037725
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1676037725
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1676037725
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1676037725
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1676037725
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1676037725
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1676037725
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1676037725
transform 1 0 39744 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1676037725
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1676037725
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1676037725
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1676037725
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1676037725
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1676037725
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1676037725
transform 1 0 37168 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1676037725
transform 1 0 42320 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1676037725
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1676037725
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1676037725
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1676037725
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1676037725
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1676037725
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1676037725
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1676037725
transform 1 0 39744 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1676037725
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1676037725
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1676037725
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1676037725
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1676037725
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1676037725
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1676037725
transform 1 0 37168 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1676037725
transform 1 0 42320 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1676037725
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1676037725
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1676037725
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1676037725
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1676037725
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1676037725
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1676037725
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1676037725
transform 1 0 39744 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1676037725
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1676037725
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1676037725
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1676037725
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1676037725
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1676037725
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1676037725
transform 1 0 37168 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1676037725
transform 1 0 42320 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1676037725
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1676037725
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1676037725
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1676037725
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1676037725
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1676037725
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1676037725
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1676037725
transform 1 0 39744 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1676037725
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1676037725
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1676037725
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1676037725
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1676037725
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1676037725
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1676037725
transform 1 0 37168 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1676037725
transform 1 0 42320 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1676037725
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1676037725
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1676037725
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1676037725
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1676037725
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1676037725
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1676037725
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1676037725
transform 1 0 39744 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1676037725
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1676037725
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1676037725
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1676037725
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1676037725
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1676037725
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1676037725
transform 1 0 37168 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1676037725
transform 1 0 42320 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1676037725
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1676037725
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1676037725
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1676037725
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1676037725
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1676037725
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1676037725
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1676037725
transform 1 0 39744 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1676037725
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1676037725
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1676037725
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1676037725
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1676037725
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1676037725
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1676037725
transform 1 0 37168 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1676037725
transform 1 0 42320 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1676037725
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1676037725
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1676037725
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1676037725
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1676037725
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1676037725
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1676037725
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1676037725
transform 1 0 39744 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1676037725
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1676037725
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1676037725
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1676037725
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1676037725
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1676037725
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1676037725
transform 1 0 37168 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1676037725
transform 1 0 42320 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1676037725
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1676037725
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1676037725
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1676037725
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1676037725
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1676037725
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1676037725
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1676037725
transform 1 0 39744 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1676037725
transform 1 0 3680 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1676037725
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1676037725
transform 1 0 8832 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1676037725
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1676037725
transform 1 0 13984 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1676037725
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1676037725
transform 1 0 19136 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1676037725
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1676037725
transform 1 0 24288 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1676037725
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1676037725
transform 1 0 29440 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1676037725
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1676037725
transform 1 0 34592 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1676037725
transform 1 0 37168 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1676037725
transform 1 0 39744 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1676037725
transform 1 0 42320 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0421_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 22632 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0422_
timestamp 1676037725
transform 1 0 21344 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0423_
timestamp 1676037725
transform 1 0 26404 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _0424_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 19412 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0425_
timestamp 1676037725
transform 1 0 23092 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0426_
timestamp 1676037725
transform 1 0 17664 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0427_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 24564 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0428_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 21344 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _0429_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 18308 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _0430_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 20148 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0431_
timestamp 1676037725
transform 1 0 17204 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _0432_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 18308 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__o2bb2a_1  _0433_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 17756 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _0434_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 18860 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__nand3b_1  _0435_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 20424 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__a211oi_2  _0436_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 19964 0 -1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__nand2_2  _0437_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 24932 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _0438_
timestamp 1676037725
transform 1 0 29716 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _0439_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 30360 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0440_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 23644 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _0441_
timestamp 1676037725
transform 1 0 22356 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0442_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 20608 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0443_
timestamp 1676037725
transform 1 0 18768 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0444_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 21252 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0445_
timestamp 1676037725
transform 1 0 23276 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__a21boi_1  _0446_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 24564 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _0447_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 23552 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0448_
timestamp 1676037725
transform 1 0 23828 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__a221oi_1  _0449_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 23920 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _0450_
timestamp 1676037725
transform 1 0 25760 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0451_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 19780 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0452_
timestamp 1676037725
transform 1 0 19964 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0453_
timestamp 1676037725
transform 1 0 21620 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _0454_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 18400 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _0455_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 17756 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0456_
timestamp 1676037725
transform 1 0 16928 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0457_
timestamp 1676037725
transform 1 0 17664 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _0458_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 13432 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0459_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 12788 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _0460_
timestamp 1676037725
transform 1 0 12696 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _0461_
timestamp 1676037725
transform 1 0 15732 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0462_
timestamp 1676037725
transform 1 0 14996 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0463_
timestamp 1676037725
transform 1 0 14076 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _0464_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 24564 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _0465_
timestamp 1676037725
transform 1 0 23736 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0466_
timestamp 1676037725
transform 1 0 23000 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _0467_
timestamp 1676037725
transform 1 0 29716 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0468_
timestamp 1676037725
transform 1 0 28612 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _0469_
timestamp 1676037725
transform 1 0 29072 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0470_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 12604 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0471_
timestamp 1676037725
transform 1 0 13892 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0472_
timestamp 1676037725
transform 1 0 10396 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0473_
timestamp 1676037725
transform 1 0 10948 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0474_
timestamp 1676037725
transform 1 0 12420 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0475_
timestamp 1676037725
transform 1 0 11684 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0476_
timestamp 1676037725
transform 1 0 10396 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0477_
timestamp 1676037725
transform 1 0 9752 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0478_
timestamp 1676037725
transform 1 0 17112 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0479_
timestamp 1676037725
transform 1 0 16468 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0480_
timestamp 1676037725
transform 1 0 20700 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0481_
timestamp 1676037725
transform 1 0 20056 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0482_
timestamp 1676037725
transform 1 0 21988 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0483_
timestamp 1676037725
transform 1 0 20792 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0484_
timestamp 1676037725
transform 1 0 22816 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0485_
timestamp 1676037725
transform 1 0 19320 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0486_
timestamp 1676037725
transform 1 0 16836 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0487_
timestamp 1676037725
transform 1 0 20240 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _0488_
timestamp 1676037725
transform 1 0 16928 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _0489_
timestamp 1676037725
transform 1 0 16100 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0490_
timestamp 1676037725
transform 1 0 14720 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0491_
timestamp 1676037725
transform 1 0 15180 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0492_
timestamp 1676037725
transform 1 0 13340 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _0493_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 25392 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _0494_
timestamp 1676037725
transform 1 0 16836 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _0495_
timestamp 1676037725
transform 1 0 13432 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0496_
timestamp 1676037725
transform 1 0 9384 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0497_
timestamp 1676037725
transform 1 0 13156 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0498_
timestamp 1676037725
transform 1 0 11776 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0499_
timestamp 1676037725
transform 1 0 7360 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0500_
timestamp 1676037725
transform 1 0 13524 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0501_
timestamp 1676037725
transform 1 0 20700 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0502_
timestamp 1676037725
transform 1 0 11960 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0503_
timestamp 1676037725
transform 1 0 7636 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _0504_
timestamp 1676037725
transform 1 0 10580 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0505_
timestamp 1676037725
transform 1 0 11868 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _0506_
timestamp 1676037725
transform 1 0 12972 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0507_
timestamp 1676037725
transform 1 0 10948 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_1  _0508_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 10580 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _0509_
timestamp 1676037725
transform 1 0 20700 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0510_
timestamp 1676037725
transform 1 0 14812 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_1  _0511_
timestamp 1676037725
transform 1 0 11684 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _0512_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 12512 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _0513_
timestamp 1676037725
transform 1 0 10764 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__xor2_1  _0514_
timestamp 1676037725
transform 1 0 9568 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__o2bb2a_1  _0515_
timestamp 1676037725
transform 1 0 14260 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _0516_
timestamp 1676037725
transform 1 0 11960 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__or4b_4  _0517_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 12788 0 1 11968
box -38 -48 1050 592
use sky130_fd_sc_hd__mux2_1  _0518_
timestamp 1676037725
transform 1 0 23276 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0519_
timestamp 1676037725
transform 1 0 22540 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _0520_
timestamp 1676037725
transform 1 0 30268 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0521_
timestamp 1676037725
transform 1 0 31280 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0522_
timestamp 1676037725
transform 1 0 29992 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0523_
timestamp 1676037725
transform 1 0 37444 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _0524_
timestamp 1676037725
transform 1 0 41492 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__and4b_1  _0525_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 35972 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__and4_1  _0526_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 36340 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0527_
timestamp 1676037725
transform 1 0 32108 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0528_
timestamp 1676037725
transform 1 0 33212 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0529_
timestamp 1676037725
transform 1 0 31464 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0530_
timestamp 1676037725
transform 1 0 33764 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0531_
timestamp 1676037725
transform 1 0 34408 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0532_
timestamp 1676037725
transform 1 0 37352 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0533_
timestamp 1676037725
transform 1 0 36524 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0534_
timestamp 1676037725
transform 1 0 37996 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _0535_
timestamp 1676037725
transform 1 0 37812 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0536_
timestamp 1676037725
transform 1 0 30176 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0537_
timestamp 1676037725
transform 1 0 43148 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _0538_
timestamp 1676037725
transform 1 0 38456 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__and4b_1  _0539_
timestamp 1676037725
transform 1 0 38272 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__a41o_1  _0540_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 35144 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _0541_
timestamp 1676037725
transform 1 0 34684 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__and4b_1  _0542_
timestamp 1676037725
transform 1 0 40112 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__or4b_1  _0543_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 40480 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__a21bo_1  _0544_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 35328 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_2  _0545_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 37076 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0546_
timestamp 1676037725
transform 1 0 30452 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _0547_
timestamp 1676037725
transform 1 0 30636 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _0548_
timestamp 1676037725
transform 1 0 33120 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _0549_
timestamp 1676037725
transform 1 0 27692 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0550_
timestamp 1676037725
transform 1 0 28612 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0551_
timestamp 1676037725
transform 1 0 37444 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nand4_1  _0552_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 35420 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _0553_
timestamp 1676037725
transform 1 0 37444 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0554_
timestamp 1676037725
transform 1 0 37444 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__a31oi_1  _0555_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 36248 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0556_
timestamp 1676037725
transform 1 0 37444 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _0557_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 31096 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _0558_
timestamp 1676037725
transform 1 0 30268 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0559_
timestamp 1676037725
transform 1 0 26404 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _0560_
timestamp 1676037725
transform 1 0 26772 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0561_
timestamp 1676037725
transform 1 0 25576 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _0562_
timestamp 1676037725
transform 1 0 28428 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _0563_
timestamp 1676037725
transform 1 0 26772 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0564_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 5152 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _0565_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 8648 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0566_
timestamp 1676037725
transform 1 0 7360 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _0567_
timestamp 1676037725
transform 1 0 19596 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_2  _0568_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 7452 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _0569_
timestamp 1676037725
transform 1 0 8280 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _0570_
timestamp 1676037725
transform 1 0 41308 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__buf_12  _0571_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 42780 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__and2_2  _0572_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 8924 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__buf_12  _0573_
timestamp 1676037725
transform 1 0 34224 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__and2_1  _0574_
timestamp 1676037725
transform 1 0 5336 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__buf_12  _0575_
timestamp 1676037725
transform 1 0 6900 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__and2_2  _0576_
timestamp 1676037725
transform 1 0 5796 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__buf_12  _0577_
timestamp 1676037725
transform 1 0 42780 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__and2_1  _0578_
timestamp 1676037725
transform 1 0 4600 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__buf_12  _0579_
timestamp 1676037725
transform 1 0 5612 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__and2_1  _0580_
timestamp 1676037725
transform 1 0 5152 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__buf_12  _0581_
timestamp 1676037725
transform 1 0 7176 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__and2_1  _0582_
timestamp 1676037725
transform 1 0 3128 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__buf_12  _0583_
timestamp 1676037725
transform 1 0 2852 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  _0584_
timestamp 1676037725
transform 1 0 41216 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0585_
timestamp 1676037725
transform 1 0 41400 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__buf_12  _0586_
timestamp 1676037725
transform 1 0 41032 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  _0587_
timestamp 1676037725
transform 1 0 15272 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0588_
timestamp 1676037725
transform 1 0 19504 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__buf_12  _0589_
timestamp 1676037725
transform 1 0 19964 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  _0590_
timestamp 1676037725
transform 1 0 32292 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_2  _0591_
timestamp 1676037725
transform 1 0 30912 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__buf_12  _0592_
timestamp 1676037725
transform 1 0 1932 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  _0593_
timestamp 1676037725
transform 1 0 23276 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0594_
timestamp 1676037725
transform 1 0 23276 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__buf_12  _0595_
timestamp 1676037725
transform 1 0 22908 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__and2_1  _0596_
timestamp 1676037725
transform 1 0 32292 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0597_
timestamp 1676037725
transform 1 0 34132 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0598_
timestamp 1676037725
transform 1 0 30268 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0599_
timestamp 1676037725
transform 1 0 27140 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_12  _0600_
timestamp 1676037725
transform 1 0 27232 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__and2_1  _0601_
timestamp 1676037725
transform 1 0 27324 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0602_
timestamp 1676037725
transform 1 0 27140 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0603_
timestamp 1676037725
transform 1 0 27416 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0604_
timestamp 1676037725
transform 1 0 26404 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0605_
timestamp 1676037725
transform 1 0 35788 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _0606_
timestamp 1676037725
transform 1 0 38088 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _0607_
timestamp 1676037725
transform 1 0 40020 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0608_
timestamp 1676037725
transform 1 0 40848 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _0609_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 32292 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0610_
timestamp 1676037725
transform 1 0 32568 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _0611_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 9844 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0612_
timestamp 1676037725
transform 1 0 9752 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _0613_
timestamp 1676037725
transform 1 0 23000 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0614_
timestamp 1676037725
transform 1 0 22540 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0615_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 26128 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0616_
timestamp 1676037725
transform 1 0 25208 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0617_
timestamp 1676037725
transform 1 0 24564 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _0618_
timestamp 1676037725
transform 1 0 25208 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _0619_
timestamp 1676037725
transform 1 0 25024 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0620_
timestamp 1676037725
transform 1 0 23276 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0621_
timestamp 1676037725
transform 1 0 23276 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0622_
timestamp 1676037725
transform 1 0 19412 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0623_
timestamp 1676037725
transform 1 0 21712 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0624_
timestamp 1676037725
transform 1 0 20608 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0625_
timestamp 1676037725
transform 1 0 19504 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0626_
timestamp 1676037725
transform 1 0 17756 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0627_
timestamp 1676037725
transform 1 0 18032 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0628_
timestamp 1676037725
transform 1 0 15088 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0629_
timestamp 1676037725
transform 1 0 16652 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0630_
timestamp 1676037725
transform 1 0 15088 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0631_
timestamp 1676037725
transform 1 0 14260 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0632_
timestamp 1676037725
transform 1 0 12972 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0633_
timestamp 1676037725
transform 1 0 12328 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0634_
timestamp 1676037725
transform 1 0 17112 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0635_
timestamp 1676037725
transform 1 0 15548 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0636__1
timestamp 1676037725
transform 1 0 13524 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0637_
timestamp 1676037725
transform 1 0 13616 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0638__2
timestamp 1676037725
transform 1 0 18124 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0639_
timestamp 1676037725
transform 1 0 16836 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0640__3
timestamp 1676037725
transform 1 0 15364 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0641_
timestamp 1676037725
transform 1 0 16008 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _0642_
timestamp 1676037725
transform 1 0 28612 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _0643_
timestamp 1676037725
transform 1 0 27784 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _0644_
timestamp 1676037725
transform 1 0 33396 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _0645_
timestamp 1676037725
transform 1 0 33120 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _0646_
timestamp 1676037725
transform 1 0 32200 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _0647_
timestamp 1676037725
transform 1 0 32384 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _0648_
timestamp 1676037725
transform 1 0 26312 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _0649_
timestamp 1676037725
transform 1 0 26128 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0650_
timestamp 1676037725
transform 1 0 35604 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0651_
timestamp 1676037725
transform 1 0 38180 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _0652_
timestamp 1676037725
transform 1 0 33396 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _0653_
timestamp 1676037725
transform 1 0 33764 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _0654_
timestamp 1676037725
transform 1 0 28888 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _0655_
timestamp 1676037725
transform 1 0 30176 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0656_
timestamp 1676037725
transform 1 0 29624 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0657_
timestamp 1676037725
transform 1 0 26588 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_8  _0658_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 27232 0 -1 8704
box -38 -48 1050 592
use sky130_fd_sc_hd__inv_2  _0659_
timestamp 1676037725
transform 1 0 27140 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0660_
timestamp 1676037725
transform 1 0 26404 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _0661_
timestamp 1676037725
transform 1 0 27508 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _0662_
timestamp 1676037725
transform 1 0 28244 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0663_
timestamp 1676037725
transform 1 0 38180 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0664_
timestamp 1676037725
transform 1 0 40020 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _0665_
timestamp 1676037725
transform 1 0 35052 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _0666_
timestamp 1676037725
transform 1 0 34132 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _0667_
timestamp 1676037725
transform 1 0 35880 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _0668_
timestamp 1676037725
transform 1 0 36616 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _0669_
timestamp 1676037725
transform 1 0 19964 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _0670_
timestamp 1676037725
transform 1 0 20148 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _0671_
timestamp 1676037725
transform 1 0 21436 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _0672_
timestamp 1676037725
transform 1 0 22172 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _0673_
timestamp 1676037725
transform 1 0 23184 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _0674_
timestamp 1676037725
transform 1 0 20056 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _0675_
timestamp 1676037725
transform 1 0 16008 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _0676_
timestamp 1676037725
transform 1 0 15364 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0677_
timestamp 1676037725
transform 1 0 14260 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0678_
timestamp 1676037725
transform 1 0 14904 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0679_
timestamp 1676037725
transform 1 0 25944 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0680_
timestamp 1676037725
transform 1 0 10948 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0681_
timestamp 1676037725
transform 1 0 11684 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0682_
timestamp 1676037725
transform 1 0 9660 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0683_
timestamp 1676037725
transform 1 0 10304 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0684_
timestamp 1676037725
transform 1 0 12328 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0685_
timestamp 1676037725
transform 1 0 14260 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0686_
timestamp 1676037725
transform 1 0 37444 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0687_
timestamp 1676037725
transform 1 0 35880 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0688_
timestamp 1676037725
transform 1 0 35236 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0689_
timestamp 1676037725
transform 1 0 36708 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0690_
timestamp 1676037725
transform 1 0 33580 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0691_
timestamp 1676037725
transform 1 0 33948 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0692_
timestamp 1676037725
transform 1 0 35696 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0693_
timestamp 1676037725
transform 1 0 35604 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0694_
timestamp 1676037725
transform 1 0 36432 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0695_
timestamp 1676037725
transform 1 0 26220 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0696_
timestamp 1676037725
transform 1 0 25024 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0697_
timestamp 1676037725
transform 1 0 25024 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0698_
timestamp 1676037725
transform 1 0 23828 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0699_
timestamp 1676037725
transform 1 0 21620 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0700_
timestamp 1676037725
transform 1 0 21896 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0701_
timestamp 1676037725
transform 1 0 20332 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0702_
timestamp 1676037725
transform 1 0 19412 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0703_
timestamp 1676037725
transform 1 0 17848 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0704_
timestamp 1676037725
transform 1 0 19412 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0705_
timestamp 1676037725
transform 1 0 18124 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0706_
timestamp 1676037725
transform 1 0 17480 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__o211ai_1  _0707_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 36432 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _0708_
timestamp 1676037725
transform 1 0 36248 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0709_
timestamp 1676037725
transform 1 0 39192 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _0710_
timestamp 1676037725
transform 1 0 39376 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _0711_
timestamp 1676037725
transform 1 0 38548 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0712_
timestamp 1676037725
transform 1 0 39376 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0713_
timestamp 1676037725
transform 1 0 39836 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__nor3_1  _0714_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 42780 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _0715_
timestamp 1676037725
transform 1 0 42596 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0716_
timestamp 1676037725
transform 1 0 39100 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0717_
timestamp 1676037725
transform 1 0 40020 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _0718_
timestamp 1676037725
transform 1 0 40020 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0719_
timestamp 1676037725
transform 1 0 39192 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0720_
timestamp 1676037725
transform 1 0 42596 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0721_
timestamp 1676037725
transform 1 0 41584 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _0722_
timestamp 1676037725
transform 1 0 42596 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _0723_
timestamp 1676037725
transform 1 0 42320 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _0724_
timestamp 1676037725
transform 1 0 40572 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0725_
timestamp 1676037725
transform 1 0 41308 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _0726_
timestamp 1676037725
transform 1 0 42596 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0727_
timestamp 1676037725
transform 1 0 33948 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0728_
timestamp 1676037725
transform 1 0 37444 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _0729_
timestamp 1676037725
transform 1 0 34960 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__a211oi_1  _0730_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 33856 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0731_
timestamp 1676037725
transform 1 0 34316 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_1  _0732_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 35236 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__or3b_1  _0733_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 35328 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__nor3b_1  _0734_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 36248 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0735_
timestamp 1676037725
transform 1 0 34868 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0736_
timestamp 1676037725
transform 1 0 33212 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0737_
timestamp 1676037725
transform 1 0 36708 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__a221oi_1  _0738_
timestamp 1676037725
transform 1 0 33856 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _0739_
timestamp 1676037725
transform 1 0 32936 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__a31oi_1  _0740_
timestamp 1676037725
transform 1 0 31004 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__a41o_1  _0741_
timestamp 1676037725
transform 1 0 31004 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _0742_
timestamp 1676037725
transform 1 0 31096 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0743_
timestamp 1676037725
transform 1 0 30452 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0744_
timestamp 1676037725
transform 1 0 33396 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _0745_
timestamp 1676037725
transform 1 0 32660 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__a41o_1  _0746_
timestamp 1676037725
transform 1 0 31556 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _0747_
timestamp 1676037725
transform 1 0 32292 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _0748_
timestamp 1676037725
transform 1 0 31096 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__o21ba_1  _0749_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 40020 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__a41o_1  _0750_
timestamp 1676037725
transform 1 0 40296 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _0751_
timestamp 1676037725
transform 1 0 42596 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0752_
timestamp 1676037725
transform 1 0 39284 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0753_
timestamp 1676037725
transform 1 0 38180 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _0754_
timestamp 1676037725
transform 1 0 38548 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__a41o_1  _0755_
timestamp 1676037725
transform 1 0 39192 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _0756_
timestamp 1676037725
transform 1 0 38824 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _0757_
timestamp 1676037725
transform 1 0 41400 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0758_
timestamp 1676037725
transform 1 0 37444 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _0759_
timestamp 1676037725
transform 1 0 34040 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _0760_
timestamp 1676037725
transform 1 0 36984 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0761_
timestamp 1676037725
transform 1 0 36248 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0762_
timestamp 1676037725
transform 1 0 37812 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0763_
timestamp 1676037725
transform 1 0 28428 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0764_
timestamp 1676037725
transform 1 0 29716 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0765_
timestamp 1676037725
transform 1 0 29716 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0766_
timestamp 1676037725
transform 1 0 31188 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0767_
timestamp 1676037725
transform 1 0 29808 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0768_
timestamp 1676037725
transform 1 0 30544 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0769_
timestamp 1676037725
transform 1 0 39836 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0770_
timestamp 1676037725
transform 1 0 39284 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0771_
timestamp 1676037725
transform 1 0 17572 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0772_
timestamp 1676037725
transform 1 0 20792 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0773_
timestamp 1676037725
transform 1 0 18308 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0774_
timestamp 1676037725
transform 1 0 18676 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0775_
timestamp 1676037725
transform 1 0 16468 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0776_
timestamp 1676037725
transform 1 0 18032 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0777_
timestamp 1676037725
transform 1 0 17296 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0778_
timestamp 1676037725
transform 1 0 17848 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0779_
timestamp 1676037725
transform 1 0 5244 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0780_
timestamp 1676037725
transform 1 0 6348 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0781_
timestamp 1676037725
transform 1 0 6532 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0782_
timestamp 1676037725
transform 1 0 7728 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0783_
timestamp 1676037725
transform 1 0 7820 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0784_
timestamp 1676037725
transform 1 0 7084 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0785_
timestamp 1676037725
transform 1 0 3956 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0786_
timestamp 1676037725
transform 1 0 2668 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0787_
timestamp 1676037725
transform 1 0 4784 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0788_
timestamp 1676037725
transform 1 0 1932 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0789_
timestamp 1676037725
transform 1 0 3956 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0790_
timestamp 1676037725
transform 1 0 5796 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0791_
timestamp 1676037725
transform 1 0 2668 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0792_
timestamp 1676037725
transform 1 0 2760 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0793_
timestamp 1676037725
transform 1 0 3956 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0794_
timestamp 1676037725
transform 1 0 2852 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _0795_
timestamp 1676037725
transform 1 0 9200 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _0796_
timestamp 1676037725
transform 1 0 8280 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _0797_
timestamp 1676037725
transform 1 0 9660 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _0798_
timestamp 1676037725
transform 1 0 10396 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _0799_
timestamp 1676037725
transform 1 0 9660 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _0800_
timestamp 1676037725
transform 1 0 10764 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _0801_
timestamp 1676037725
transform 1 0 28336 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_2  _0802_
timestamp 1676037725
transform 1 0 16560 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0803_
timestamp 1676037725
transform 1 0 12696 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0804_
timestamp 1676037725
transform 1 0 11868 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0805_
timestamp 1676037725
transform 1 0 14260 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0806_
timestamp 1676037725
transform 1 0 14260 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0807_
timestamp 1676037725
transform 1 0 15088 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0808_
timestamp 1676037725
transform 1 0 15364 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0809_
timestamp 1676037725
transform 1 0 11224 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0810_
timestamp 1676037725
transform 1 0 10948 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _0811_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 11684 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _0812_
timestamp 1676037725
transform 1 0 10856 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0813_
timestamp 1676037725
transform 1 0 7636 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0814_
timestamp 1676037725
transform 1 0 8372 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _0815_
timestamp 1676037725
transform 1 0 6624 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _0816_
timestamp 1676037725
transform 1 0 7176 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0817_
timestamp 1676037725
transform 1 0 6256 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _0818_
timestamp 1676037725
transform 1 0 5704 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0819_
timestamp 1676037725
transform 1 0 5612 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0820_
timestamp 1676037725
transform 1 0 6532 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0821_
timestamp 1676037725
transform 1 0 5796 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _0822_
timestamp 1676037725
transform 1 0 4968 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0823_
timestamp 1676037725
transform 1 0 4692 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0824_
timestamp 1676037725
transform 1 0 3220 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0825_
timestamp 1676037725
transform 1 0 4324 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0826_
timestamp 1676037725
transform 1 0 6532 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0827_
timestamp 1676037725
transform 1 0 5612 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0828_
timestamp 1676037725
transform 1 0 4968 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0829_
timestamp 1676037725
transform 1 0 3956 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0830_
timestamp 1676037725
transform 1 0 5612 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _0831_
timestamp 1676037725
transform 1 0 4600 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0832_
timestamp 1676037725
transform 1 0 3220 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0833_
timestamp 1676037725
transform 1 0 27508 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0834_
timestamp 1676037725
transform 1 0 28428 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _0835_
timestamp 1676037725
transform 1 0 25852 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _0836_
timestamp 1676037725
transform 1 0 25760 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _0837_
timestamp 1676037725
transform 1 0 14260 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _0838_
timestamp 1676037725
transform 1 0 16100 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0839_
timestamp 1676037725
transform 1 0 12604 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0840_
timestamp 1676037725
transform 1 0 12144 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0841_
timestamp 1676037725
transform 1 0 19136 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0842_
timestamp 1676037725
transform 1 0 19412 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _0843_
timestamp 1676037725
transform 1 0 20792 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _0844_
timestamp 1676037725
transform 1 0 20424 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _0845_
timestamp 1676037725
transform 1 0 27140 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _0846_
timestamp 1676037725
transform 1 0 26772 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _0847_
timestamp 1676037725
transform 1 0 24656 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _0848_
timestamp 1676037725
transform 1 0 25852 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0849_
timestamp 1676037725
transform 1 0 28336 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0850_
timestamp 1676037725
transform 1 0 29716 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0851_
timestamp 1676037725
transform 1 0 30176 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _0852_
timestamp 1676037725
transform 1 0 37168 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _0853_
timestamp 1676037725
transform 1 0 38824 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _0854_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 23184 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0855_
timestamp 1676037725
transform 1 0 24564 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfxtp_1  _0856_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 23092 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0857_
timestamp 1676037725
transform 1 0 19872 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0858_
timestamp 1676037725
transform 1 0 19872 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0859_
timestamp 1676037725
transform 1 0 17204 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0860_
timestamp 1676037725
transform 1 0 14812 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0861_
timestamp 1676037725
transform 1 0 14260 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0862_
timestamp 1676037725
transform 1 0 13248 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0863_
timestamp 1676037725
transform 1 0 15272 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0864_
timestamp 1676037725
transform 1 0 27784 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0865_
timestamp 1676037725
transform 1 0 27784 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0866_
timestamp 1676037725
transform 1 0 28520 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0867_
timestamp 1676037725
transform 1 0 38732 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0868_
timestamp 1676037725
transform 1 0 14904 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0869_
timestamp 1676037725
transform 1 0 16192 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0870_
timestamp 1676037725
transform 1 0 14904 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0871_
timestamp 1676037725
transform 1 0 16836 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _0872__27 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 14536 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__dfstp_1  _0872_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 14444 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_1  _0873_
timestamp 1676037725
transform 1 0 15824 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_4  _0874_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 17664 0 -1 3264
box -38 -48 2246 592
use sky130_fd_sc_hd__dfstp_2  _0875_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 26220 0 1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _0876_
timestamp 1676037725
transform 1 0 31188 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0877_
timestamp 1676037725
transform 1 0 30912 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0878_
timestamp 1676037725
transform 1 0 25116 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0879_
timestamp 1676037725
transform 1 0 37168 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0880_
timestamp 1676037725
transform 1 0 32476 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0881_
timestamp 1676037725
transform 1 0 27968 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _0882_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 27140 0 -1 7616
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _0883_
timestamp 1676037725
transform 1 0 26128 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _0884_
timestamp 1676037725
transform 1 0 27140 0 -1 10880
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _0885_
timestamp 1676037725
transform 1 0 38364 0 -1 13056
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _0886_
timestamp 1676037725
transform 1 0 34868 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0887_
timestamp 1676037725
transform 1 0 34868 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0888_
timestamp 1676037725
transform 1 0 20792 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0889_
timestamp 1676037725
transform 1 0 20700 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  _0890_
timestamp 1676037725
transform 1 0 20516 0 1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _0891_
timestamp 1676037725
transform 1 0 16836 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  _0892_
timestamp 1676037725
transform 1 0 10304 0 1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _0893_
timestamp 1676037725
transform 1 0 11684 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0894_
timestamp 1676037725
transform 1 0 10396 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0895_
timestamp 1676037725
transform 1 0 11684 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfxtp_1  _0896_
timestamp 1676037725
transform 1 0 36340 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0897_
timestamp 1676037725
transform 1 0 34592 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0898_
timestamp 1676037725
transform 1 0 34868 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0899_
timestamp 1676037725
transform 1 0 24840 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0900_
timestamp 1676037725
transform 1 0 21988 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0901_
timestamp 1676037725
transform 1 0 18492 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0902_
timestamp 1676037725
transform 1 0 17112 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0903_
timestamp 1676037725
transform 1 0 40664 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0904_
timestamp 1676037725
transform 1 0 40664 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0905_
timestamp 1676037725
transform 1 0 40940 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0906_
timestamp 1676037725
transform 1 0 42504 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0907_
timestamp 1676037725
transform 1 0 40756 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0908_
timestamp 1676037725
transform 1 0 34868 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0909_
timestamp 1676037725
transform 1 0 35420 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0910_
timestamp 1676037725
transform 1 0 33580 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0911_
timestamp 1676037725
transform 1 0 30268 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0912_
timestamp 1676037725
transform 1 0 29716 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0913_
timestamp 1676037725
transform 1 0 41308 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0914_
timestamp 1676037725
transform 1 0 40480 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0915_
timestamp 1676037725
transform 1 0 35144 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0916_
timestamp 1676037725
transform 1 0 40664 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0917_
timestamp 1676037725
transform 1 0 18952 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0918_
timestamp 1676037725
transform 1 0 30728 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0919_
timestamp 1676037725
transform 1 0 24748 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0920_
timestamp 1676037725
transform 1 0 29256 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0921_
timestamp 1676037725
transform 1 0 33028 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0922_
timestamp 1676037725
transform 1 0 31004 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0923_
timestamp 1676037725
transform 1 0 40020 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0924_
timestamp 1676037725
transform 1 0 23000 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0925_
timestamp 1676037725
transform 1 0 19320 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0926_
timestamp 1676037725
transform 1 0 17480 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0927_
timestamp 1676037725
transform 1 0 17480 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0928_
timestamp 1676037725
transform 1 0 6532 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0929_
timestamp 1676037725
transform 1 0 6532 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0930_
timestamp 1676037725
transform 1 0 6532 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0931_
timestamp 1676037725
transform 1 0 2116 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0932_
timestamp 1676037725
transform 1 0 3956 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0933_
timestamp 1676037725
transform 1 0 3956 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0934_
timestamp 1676037725
transform 1 0 2024 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0935_
timestamp 1676037725
transform 1 0 2484 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0936_
timestamp 1676037725
transform 1 0 8372 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0937_
timestamp 1676037725
transform 1 0 5888 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0938_
timestamp 1676037725
transform 1 0 7728 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0939_
timestamp 1676037725
transform 1 0 3312 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0940_
timestamp 1676037725
transform 1 0 3956 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0941_
timestamp 1676037725
transform 1 0 2024 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0942_
timestamp 1676037725
transform 1 0 3956 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0943_
timestamp 1676037725
transform 1 0 2024 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfrtp_1  _0944_
timestamp 1676037725
transform 1 0 6900 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0945_
timestamp 1676037725
transform 1 0 9108 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0946_
timestamp 1676037725
transform 1 0 9108 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfxtp_2  _0947_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 10488 0 1 7616
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _0948_
timestamp 1676037725
transform 1 0 12972 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0949_
timestamp 1676037725
transform 1 0 13524 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0950_
timestamp 1676037725
transform 1 0 11500 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0951_
timestamp 1676037725
transform 1 0 7084 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0952_
timestamp 1676037725
transform 1 0 6532 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0953_
timestamp 1676037725
transform 1 0 3956 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0954_
timestamp 1676037725
transform 1 0 5520 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0955_
timestamp 1676037725
transform 1 0 3772 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _0956_
timestamp 1676037725
transform 1 0 22172 0 -1 8704
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _0957_
timestamp 1676037725
transform 1 0 10120 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0958_
timestamp 1676037725
transform 1 0 11868 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0959_
timestamp 1676037725
transform 1 0 22264 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfrtp_1  _0960_
timestamp 1676037725
transform 1 0 28060 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0961_
timestamp 1676037725
transform 1 0 24564 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0962_
timestamp 1676037725
transform 1 0 13524 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0963_
timestamp 1676037725
transform 1 0 11776 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0964_
timestamp 1676037725
transform 1 0 17112 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0965_
timestamp 1676037725
transform 1 0 19412 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0966_
timestamp 1676037725
transform 1 0 25576 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0967_
timestamp 1676037725
transform 1 0 23644 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _0968_
timestamp 1676037725
transform 1 0 29348 0 -1 4352
box -38 -48 2154 592
use sky130_fd_sc_hd__dfxtp_1  _0969_
timestamp 1676037725
transform 1 0 38364 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  _1009_
timestamp 1676037725
transform 1 0 42780 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 22172 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_scan_clk_in
timestamp 1676037725
transform 1 0 5244 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_scan_clk_in
timestamp 1676037725
transform 1 0 2576 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_scan_clk_in
timestamp 1676037725
transform 1 0 5244 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_0__f_clk
timestamp 1676037725
transform 1 0 10396 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_1__f_clk
timestamp 1676037725
transform 1 0 12972 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_2__f_clk
timestamp 1676037725
transform 1 0 7820 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_3__f_clk
timestamp 1676037725
transform 1 0 12972 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_4__f_clk
timestamp 1676037725
transform 1 0 28612 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_5__f_clk
timestamp 1676037725
transform 1 0 31188 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_6__f_clk
timestamp 1676037725
transform 1 0 29624 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_7__f_clk
timestamp 1676037725
transform 1 0 34684 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 11960 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  input1
timestamp 1676037725
transform 1 0 1564 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1676037725
transform 1 0 43884 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1676037725
transform 1 0 44160 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1676037725
transform 1 0 37444 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1676037725
transform 1 0 31004 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1676037725
transform 1 0 25852 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1676037725
transform 1 0 44160 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input8 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 2300 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input9
timestamp 1676037725
transform 1 0 3128 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input10
timestamp 1676037725
transform 1 0 27140 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input11
timestamp 1676037725
transform 1 0 1564 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input12
timestamp 1676037725
transform 1 0 32292 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input13
timestamp 1676037725
transform 1 0 11684 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input14 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 32292 0 -1 17408
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input15
timestamp 1676037725
transform 1 0 38732 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input16
timestamp 1676037725
transform 1 0 4600 0 -1 17408
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input17
timestamp 1676037725
transform 1 0 12880 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input18
timestamp 1676037725
transform 1 0 1564 0 -1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input19
timestamp 1676037725
transform 1 0 42596 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input20
timestamp 1676037725
transform 1 0 44160 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input21
timestamp 1676037725
transform 1 0 1564 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input22
timestamp 1676037725
transform 1 0 24564 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input23
timestamp 1676037725
transform 1 0 34868 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input24
timestamp 1676037725
transform 1 0 17480 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  input25
timestamp 1676037725
transform 1 0 16836 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input26
timestamp 1676037725
transform 1 0 9752 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  scan_controller_28
timestamp 1676037725
transform 1 0 12972 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  scan_controller_29
timestamp 1676037725
transform 1 0 13524 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  scan_controller_30
timestamp 1676037725
transform 1 0 44160 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  scan_controller_31
timestamp 1676037725
transform 1 0 35512 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  scan_controller_32
timestamp 1676037725
transform 1 0 44160 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  scan_controller_33
timestamp 1676037725
transform 1 0 19412 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  scan_controller_34
timestamp 1676037725
transform 1 0 4600 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  scan_controller_35
timestamp 1676037725
transform 1 0 1564 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  scan_controller_36
timestamp 1676037725
transform 1 0 43240 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  scan_controller_37
timestamp 1676037725
transform 1 0 1564 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  scan_controller_38
timestamp 1676037725
transform 1 0 20700 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  scan_controller_39
timestamp 1676037725
transform 1 0 44160 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  scan_controller_40
timestamp 1676037725
transform 1 0 44160 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  scan_controller_41
timestamp 1676037725
transform 1 0 29716 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  scan_controller_42
timestamp 1676037725
transform 1 0 37444 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  scan_controller_43
timestamp 1676037725
transform 1 0 3956 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  scan_controller_44
timestamp 1676037725
transform 1 0 7820 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  scan_controller_45
timestamp 1676037725
transform 1 0 11684 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  scan_controller_46
timestamp 1676037725
transform 1 0 43884 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  scan_controller_47
timestamp 1676037725
transform 1 0 44160 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  scan_controller_48
timestamp 1676037725
transform 1 0 42596 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  scan_controller_49
timestamp 1676037725
transform 1 0 7820 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  scan_controller_50
timestamp 1676037725
transform 1 0 24564 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  scan_controller_51
timestamp 1676037725
transform 1 0 40020 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  scan_controller_52
timestamp 1676037725
transform 1 0 6532 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  scan_controller_53
timestamp 1676037725
transform 1 0 19412 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  scan_controller_54
timestamp 1676037725
transform 1 0 14260 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  scan_controller_55
timestamp 1676037725
transform 1 0 30360 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  scan_controller_56
timestamp 1676037725
transform 1 0 25852 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  scan_controller_57
timestamp 1676037725
transform 1 0 38732 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  scan_controller_58
timestamp 1676037725
transform 1 0 1564 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  scan_controller_59
timestamp 1676037725
transform 1 0 1564 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  scan_controller_60
timestamp 1676037725
transform 1 0 22632 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  scan_controller_61
timestamp 1676037725
transform 1 0 29716 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  scan_controller_62
timestamp 1676037725
transform 1 0 1564 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  scan_controller_63
timestamp 1676037725
transform 1 0 2208 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  scan_controller_64
timestamp 1676037725
transform 1 0 1564 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  scan_controller_65
timestamp 1676037725
transform 1 0 27784 0 -1 17408
box -38 -48 314 592
<< labels >>
flabel metal2 s 1278 19200 1390 20000 0 FreeSans 448 90 0 0 active_select[0]
port 0 nsew signal input
flabel metal2 s 43782 0 43894 800 0 FreeSans 448 90 0 0 active_select[1]
port 1 nsew signal input
flabel metal2 s 45070 0 45182 800 0 FreeSans 448 90 0 0 active_select[2]
port 2 nsew signal input
flabel metal2 s 36698 0 36810 800 0 FreeSans 448 90 0 0 active_select[3]
port 3 nsew signal input
flabel metal2 s 30902 19200 31014 20000 0 FreeSans 448 90 0 0 active_select[4]
port 4 nsew signal input
flabel metal2 s 25750 0 25862 800 0 FreeSans 448 90 0 0 active_select[5]
port 5 nsew signal input
flabel metal3 s 45200 7428 46000 7668 0 FreeSans 960 0 0 0 active_select[6]
port 6 nsew signal input
flabel metal3 s 0 16948 800 17188 0 FreeSans 960 0 0 0 active_select[7]
port 7 nsew signal input
flabel metal2 s 3210 19200 3322 20000 0 FreeSans 448 90 0 0 active_select[8]
port 8 nsew signal input
flabel metal2 s 33478 0 33590 800 0 FreeSans 448 90 0 0 clk
port 9 nsew signal input
flabel metal2 s 27038 0 27150 800 0 FreeSans 448 90 0 0 driver_sel[0]
port 10 nsew signal input
flabel metal2 s -10 19200 102 20000 0 FreeSans 448 90 0 0 driver_sel[1]
port 11 nsew signal input
flabel metal2 s 32190 0 32302 800 0 FreeSans 448 90 0 0 inputs[0]
port 12 nsew signal input
flabel metal2 s 10938 19200 11050 20000 0 FreeSans 448 90 0 0 inputs[1]
port 13 nsew signal input
flabel metal2 s 32190 19200 32302 20000 0 FreeSans 448 90 0 0 inputs[2]
port 14 nsew signal input
flabel metal2 s 38630 19200 38742 20000 0 FreeSans 448 90 0 0 inputs[3]
port 15 nsew signal input
flabel metal2 s 4498 19200 4610 20000 0 FreeSans 448 90 0 0 inputs[4]
port 16 nsew signal input
flabel metal2 s 12870 0 12982 800 0 FreeSans 448 90 0 0 inputs[5]
port 17 nsew signal input
flabel metal3 s 0 4708 800 4948 0 FreeSans 960 0 0 0 inputs[6]
port 18 nsew signal input
flabel metal2 s 41850 0 41962 800 0 FreeSans 448 90 0 0 inputs[7]
port 19 nsew signal input
flabel metal3 s 45200 8788 46000 9028 0 FreeSans 960 0 0 0 la_scan_clk_in
port 20 nsew signal input
flabel metal3 s 0 8108 800 8348 0 FreeSans 960 0 0 0 la_scan_data_in
port 21 nsew signal input
flabel metal3 s 45200 14228 46000 14468 0 FreeSans 960 0 0 0 la_scan_data_out
port 22 nsew signal tristate
flabel metal2 s 23818 19200 23930 20000 0 FreeSans 448 90 0 0 la_scan_latch_en
port 23 nsew signal input
flabel metal2 s 34122 19200 34234 20000 0 FreeSans 448 90 0 0 la_scan_select
port 24 nsew signal input
flabel metal2 s 12870 19200 12982 20000 0 FreeSans 448 90 0 0 oeb[0]
port 25 nsew signal tristate
flabel metal2 s 20598 0 20710 800 0 FreeSans 448 90 0 0 oeb[10]
port 26 nsew signal tristate
flabel metal3 s 45200 12188 46000 12428 0 FreeSans 960 0 0 0 oeb[11]
port 27 nsew signal tristate
flabel metal3 s 45200 15588 46000 15828 0 FreeSans 960 0 0 0 oeb[12]
port 28 nsew signal tristate
flabel metal2 s 28970 0 29082 800 0 FreeSans 448 90 0 0 oeb[13]
port 29 nsew signal tristate
flabel metal2 s 37342 19200 37454 20000 0 FreeSans 448 90 0 0 oeb[14]
port 30 nsew signal tristate
flabel metal2 s 3210 0 3322 800 0 FreeSans 448 90 0 0 oeb[15]
port 31 nsew signal tristate
flabel metal2 s 7718 19200 7830 20000 0 FreeSans 448 90 0 0 oeb[16]
port 32 nsew signal tristate
flabel metal2 s 10938 0 11050 800 0 FreeSans 448 90 0 0 oeb[17]
port 33 nsew signal tristate
flabel metal2 s 43782 19200 43894 20000 0 FreeSans 448 90 0 0 oeb[18]
port 34 nsew signal tristate
flabel metal3 s 45200 10828 46000 11068 0 FreeSans 960 0 0 0 oeb[19]
port 35 nsew signal tristate
flabel metal2 s 16090 0 16202 800 0 FreeSans 448 90 0 0 oeb[1]
port 36 nsew signal tristate
flabel metal2 s 41850 19200 41962 20000 0 FreeSans 448 90 0 0 oeb[20]
port 37 nsew signal tristate
flabel metal2 s 7718 0 7830 800 0 FreeSans 448 90 0 0 oeb[21]
port 38 nsew signal tristate
flabel metal2 s 23818 0 23930 800 0 FreeSans 448 90 0 0 oeb[22]
port 39 nsew signal tristate
flabel metal2 s 39918 0 40030 800 0 FreeSans 448 90 0 0 oeb[23]
port 40 nsew signal tristate
flabel metal2 s 6430 19200 6542 20000 0 FreeSans 448 90 0 0 oeb[24]
port 41 nsew signal tristate
flabel metal2 s 19310 0 19422 800 0 FreeSans 448 90 0 0 oeb[25]
port 42 nsew signal tristate
flabel metal2 s 14158 19200 14270 20000 0 FreeSans 448 90 0 0 oeb[26]
port 43 nsew signal tristate
flabel metal2 s 30258 0 30370 800 0 FreeSans 448 90 0 0 oeb[27]
port 44 nsew signal tristate
flabel metal2 s 25750 19200 25862 20000 0 FreeSans 448 90 0 0 oeb[28]
port 45 nsew signal tristate
flabel metal2 s 38630 0 38742 800 0 FreeSans 448 90 0 0 oeb[29]
port 46 nsew signal tristate
flabel metal3 s 45200 628 46000 868 0 FreeSans 960 0 0 0 oeb[2]
port 47 nsew signal tristate
flabel metal3 s 0 6748 800 6988 0 FreeSans 960 0 0 0 oeb[30]
port 48 nsew signal tristate
flabel metal3 s 0 1308 800 1548 0 FreeSans 960 0 0 0 oeb[31]
port 49 nsew signal tristate
flabel metal2 s 22530 19200 22642 20000 0 FreeSans 448 90 0 0 oeb[32]
port 50 nsew signal tristate
flabel metal2 s 28970 19200 29082 20000 0 FreeSans 448 90 0 0 oeb[33]
port 51 nsew signal tristate
flabel metal3 s 0 3348 800 3588 0 FreeSans 960 0 0 0 oeb[34]
port 52 nsew signal tristate
flabel metal2 s -10 0 102 800 0 FreeSans 448 90 0 0 oeb[35]
port 53 nsew signal tristate
flabel metal3 s 0 18308 800 18548 0 FreeSans 960 0 0 0 oeb[36]
port 54 nsew signal tristate
flabel metal2 s 27682 19200 27794 20000 0 FreeSans 448 90 0 0 oeb[37]
port 55 nsew signal tristate
flabel metal2 s 35410 19200 35522 20000 0 FreeSans 448 90 0 0 oeb[3]
port 56 nsew signal tristate
flabel metal2 s 45070 19200 45182 20000 0 FreeSans 448 90 0 0 oeb[4]
port 57 nsew signal tristate
flabel metal2 s 19310 19200 19422 20000 0 FreeSans 448 90 0 0 oeb[5]
port 58 nsew signal tristate
flabel metal2 s 4498 0 4610 800 0 FreeSans 448 90 0 0 oeb[6]
port 59 nsew signal tristate
flabel metal2 s 1278 0 1390 800 0 FreeSans 448 90 0 0 oeb[7]
port 60 nsew signal tristate
flabel metal3 s 45200 18988 46000 19228 0 FreeSans 960 0 0 0 oeb[8]
port 61 nsew signal tristate
flabel metal3 s 0 13548 800 13788 0 FreeSans 960 0 0 0 oeb[9]
port 62 nsew signal tristate
flabel metal2 s 14158 0 14270 800 0 FreeSans 448 90 0 0 outputs[0]
port 63 nsew signal tristate
flabel metal3 s 45200 17628 46000 17868 0 FreeSans 960 0 0 0 outputs[1]
port 64 nsew signal tristate
flabel metal2 s 35410 0 35522 800 0 FreeSans 448 90 0 0 outputs[2]
port 65 nsew signal tristate
flabel metal2 s 17378 19200 17490 20000 0 FreeSans 448 90 0 0 outputs[3]
port 66 nsew signal tristate
flabel metal3 s 45200 4028 46000 4268 0 FreeSans 960 0 0 0 outputs[4]
port 67 nsew signal tristate
flabel metal2 s 6430 0 6542 800 0 FreeSans 448 90 0 0 outputs[5]
port 68 nsew signal tristate
flabel metal2 s 9650 0 9762 800 0 FreeSans 448 90 0 0 outputs[6]
port 69 nsew signal tristate
flabel metal3 s 0 14908 800 15148 0 FreeSans 960 0 0 0 outputs[7]
port 70 nsew signal tristate
flabel metal3 s 45200 5388 46000 5628 0 FreeSans 960 0 0 0 ready
port 71 nsew signal tristate
flabel metal2 s 17378 0 17490 800 0 FreeSans 448 90 0 0 reset
port 72 nsew signal input
flabel metal3 s 0 11508 800 11748 0 FreeSans 960 0 0 0 scan_clk_in
port 73 nsew signal input
flabel metal2 s 40562 19200 40674 20000 0 FreeSans 448 90 0 0 scan_clk_out
port 74 nsew signal tristate
flabel metal2 s 16090 19200 16202 20000 0 FreeSans 448 90 0 0 scan_data_in
port 75 nsew signal input
flabel metal2 s 20598 19200 20710 20000 0 FreeSans 448 90 0 0 scan_data_out
port 76 nsew signal tristate
flabel metal2 s 22530 0 22642 800 0 FreeSans 448 90 0 0 scan_latch_en
port 77 nsew signal tristate
flabel metal3 s 0 10148 800 10388 0 FreeSans 960 0 0 0 scan_select
port 78 nsew signal tristate
flabel metal2 s 9650 19200 9762 20000 0 FreeSans 448 90 0 0 set_clk_div
port 79 nsew signal input
flabel metal3 s 45200 1988 46000 2228 0 FreeSans 960 0 0 0 slow_clk
port 80 nsew signal tristate
flabel metal4 s 6417 2128 6737 17456 0 FreeSans 1920 90 0 0 vccd1
port 81 nsew power bidirectional
flabel metal4 s 17364 2128 17684 17456 0 FreeSans 1920 90 0 0 vccd1
port 81 nsew power bidirectional
flabel metal4 s 28311 2128 28631 17456 0 FreeSans 1920 90 0 0 vccd1
port 81 nsew power bidirectional
flabel metal4 s 39258 2128 39578 17456 0 FreeSans 1920 90 0 0 vccd1
port 81 nsew power bidirectional
flabel metal4 s 11890 2128 12210 17456 0 FreeSans 1920 90 0 0 vssd1
port 82 nsew ground bidirectional
flabel metal4 s 22837 2128 23157 17456 0 FreeSans 1920 90 0 0 vssd1
port 82 nsew ground bidirectional
flabel metal4 s 33784 2128 34104 17456 0 FreeSans 1920 90 0 0 vssd1
port 82 nsew ground bidirectional
flabel metal4 s 44731 2128 45051 17456 0 FreeSans 1920 90 0 0 vssd1
port 82 nsew ground bidirectional
rlabel metal1 23000 16864 23000 16864 0 vccd1
rlabel via1 23077 17408 23077 17408 0 vssd1
rlabel metal1 40940 12614 40940 12614 0 _0000_
rlabel metal1 32614 13192 32614 13192 0 _0001_
rlabel metal1 10288 7786 10288 7786 0 _0002_
rlabel metal2 7222 5406 7222 5406 0 _0003_
rlabel metal2 26450 12002 26450 12002 0 _0004_
rlabel metal1 27324 9690 27324 9690 0 _0005_
rlabel metal1 35190 12104 35190 12104 0 _0006_
rlabel metal1 26404 7854 26404 7854 0 _0007_
rlabel metal1 31372 14042 31372 14042 0 _0008_
rlabel metal1 30774 11186 30774 11186 0 _0009_
rlabel metal2 26818 10710 26818 10710 0 _0010_
rlabel metal2 37490 12376 37490 12376 0 _0011_
rlabel metal1 32982 10574 32982 10574 0 _0012_
rlabel metal2 28290 13022 28290 13022 0 _0013_
rlabel metal1 22540 8058 22540 8058 0 _0014_
rlabel metal2 24610 12614 24610 12614 0 _0015_
rlabel metal1 25208 9350 25208 9350 0 _0016_
rlabel metal2 15226 3230 15226 3230 0 _0017_
rlabel metal1 14490 2924 14490 2924 0 _0018_
rlabel metal1 16376 3910 16376 3910 0 _0019_
rlabel metal1 16606 3162 16606 3162 0 _0020_
rlabel metal1 19090 2985 19090 2985 0 _0021_
rlabel metal1 16698 2618 16698 2618 0 _0022_
rlabel metal1 27745 7786 27745 7786 0 _0023_
rlabel metal1 32943 12138 32943 12138 0 _0024_
rlabel metal1 32384 9418 32384 9418 0 _0025_
rlabel metal1 26312 10234 26312 10234 0 _0026_
rlabel metal1 38180 13158 38180 13158 0 _0027_
rlabel metal1 33672 10982 33672 10982 0 _0028_
rlabel metal1 30222 12920 30222 12920 0 _0029_
rlabel metal1 27278 6630 27278 6630 0 _0030_
rlabel metal1 26680 12614 26680 12614 0 _0031_
rlabel metal1 28244 10234 28244 10234 0 _0032_
rlabel metal1 39981 12886 39981 12886 0 _0033_
rlabel metal1 34730 9894 34730 9894 0 _0034_
rlabel metal1 36616 12614 36616 12614 0 _0035_
rlabel metal1 20700 8806 20700 8806 0 _0036_
rlabel metal2 22126 11594 22126 11594 0 _0037_
rlabel metal1 20700 10506 20700 10506 0 _0038_
rlabel metal1 16192 10778 16192 10778 0 _0039_
rlabel metal1 14950 9928 14950 9928 0 _0040_
rlabel metal1 11684 6630 11684 6630 0 _0041_
rlabel metal2 10350 8704 10350 8704 0 _0042_
rlabel metal1 13708 9146 13708 9146 0 _0043_
rlabel metal2 8326 5644 8326 5644 0 _0044_
rlabel metal2 10442 5032 10442 5032 0 _0045_
rlabel metal1 10764 6426 10764 6426 0 _0046_
rlabel metal2 29026 5678 29026 5678 0 _0047_
rlabel metal1 25852 6630 25852 6630 0 _0048_
rlabel metal1 16008 5542 16008 5542 0 _0049_
rlabel metal2 12190 4760 12190 4760 0 _0050_
rlabel metal2 19458 4114 19458 4114 0 _0051_
rlabel metal1 20608 3706 20608 3706 0 _0052_
rlabel metal1 26864 3706 26864 3706 0 _0053_
rlabel metal1 25898 4216 25898 4216 0 _0054_
rlabel metal1 29939 4182 29939 4182 0 _0055_
rlabel metal1 23046 12750 23046 12750 0 _0056_
rlabel via1 23409 7446 23409 7446 0 _0057_
rlabel metal1 20971 7446 20971 7446 0 _0058_
rlabel metal1 19862 7854 19862 7854 0 _0059_
rlabel metal1 17797 8466 17797 8466 0 _0060_
rlabel metal1 15911 7786 15911 7786 0 _0061_
rlabel via1 14577 5610 14577 5610 0 _0062_
rlabel metal2 13386 7174 13386 7174 0 _0063_
rlabel metal2 15594 6562 15594 6562 0 _0064_
rlabel metal1 21022 9010 21022 9010 0 _0065_
rlabel metal2 21022 11628 21022 11628 0 _0066_
rlabel metal1 20884 10030 20884 10030 0 _0067_
rlabel metal2 16514 10404 16514 10404 0 _0068_
rlabel metal2 10718 10540 10718 10540 0 _0069_
rlabel metal1 11776 7514 11776 7514 0 _0070_
rlabel metal2 10994 8738 10994 8738 0 _0071_
rlabel metal1 13938 9418 13938 9418 0 _0072_
rlabel via1 36652 13294 36652 13294 0 _0073_
rlabel metal1 34438 15062 34438 15062 0 _0074_
rlabel metal1 35829 14314 35829 14314 0 _0075_
rlabel via1 25157 14994 25157 14994 0 _0076_
rlabel metal2 21942 14110 21942 14110 0 _0077_
rlabel metal1 18338 13974 18338 13974 0 _0078_
rlabel metal1 17388 14586 17388 14586 0 _0079_
rlabel metal1 40142 8874 40142 8874 0 _0080_
rlabel metal1 42642 10744 42642 10744 0 _0081_
rlabel metal1 40930 10030 40930 10030 0 _0082_
rlabel metal1 42596 8058 42596 8058 0 _0083_
rlabel metal2 42642 5882 42642 5882 0 _0084_
rlabel metal1 34996 5678 34996 5678 0 _0085_
rlabel metal1 35236 4794 35236 4794 0 _0086_
rlabel metal1 33800 5202 33800 5202 0 _0087_
rlabel metal1 30544 6426 30544 6426 0 _0088_
rlabel metal1 31096 6426 31096 6426 0 _0089_
rlabel metal1 39330 6664 39330 6664 0 _0090_
rlabel metal2 41446 7650 41446 7650 0 _0091_
rlabel metal1 36657 7786 36657 7786 0 _0092_
rlabel via1 29573 9554 29573 9554 0 _0093_
rlabel metal2 31234 14382 31234 14382 0 _0094_
rlabel metal1 31224 14382 31224 14382 0 _0095_
rlabel metal1 39820 14314 39820 14314 0 _0096_
rlabel metal1 23220 14994 23220 14994 0 _0097_
rlabel metal1 19540 12818 19540 12818 0 _0098_
rlabel metal1 17935 12818 17935 12818 0 _0099_
rlabel via1 17797 13226 17797 13226 0 _0100_
rlabel metal1 6624 6630 6624 6630 0 _0101_
rlabel metal1 7774 11186 7774 11186 0 _0102_
rlabel metal1 7948 7378 7948 7378 0 _0103_
rlabel metal1 3158 10710 3158 10710 0 _0104_
rlabel via1 4273 6358 4273 6358 0 _0105_
rlabel metal1 3123 6290 3123 6290 0 _0106_
rlabel metal1 3526 5610 3526 5610 0 _0107_
rlabel metal2 2898 10642 2898 10642 0 _0108_
rlabel metal1 12834 13192 12834 13192 0 _0109_
rlabel metal1 14623 13974 14623 13974 0 _0110_
rlabel metal1 11346 14314 11346 14314 0 _0111_
rlabel metal1 7304 14382 7304 14382 0 _0112_
rlabel via1 6849 13974 6849 13974 0 _0113_
rlabel metal1 3756 13226 3756 13226 0 _0114_
rlabel viali 5837 12206 5837 12206 0 _0115_
rlabel metal1 3992 11730 3992 11730 0 _0116_
rlabel metal1 28750 5134 28750 5134 0 _0117_
rlabel metal2 23046 6018 23046 6018 0 _0118_
rlabel metal1 13984 4250 13984 4250 0 _0119_
rlabel metal2 12742 4454 12742 4454 0 _0120_
rlabel metal1 17572 4250 17572 4250 0 _0121_
rlabel metal1 21666 4692 21666 4692 0 _0122_
rlabel metal2 25898 4760 25898 4760 0 _0123_
rlabel metal1 23920 3706 23920 3706 0 _0124_
rlabel metal1 30038 4046 30038 4046 0 _0125_
rlabel metal1 38778 11322 38778 11322 0 _0126_
rlabel metal1 20470 6324 20470 6324 0 _0127_
rlabel metal1 19642 5678 19642 5678 0 _0128_
rlabel metal1 19458 5746 19458 5746 0 _0129_
rlabel metal1 20102 5882 20102 5882 0 _0130_
rlabel metal1 21252 6698 21252 6698 0 _0131_
rlabel metal1 18814 6766 18814 6766 0 _0132_
rlabel metal1 21390 6800 21390 6800 0 _0133_
rlabel metal1 20562 5712 20562 5712 0 _0134_
rlabel metal1 19550 6766 19550 6766 0 _0135_
rlabel metal2 20746 6154 20746 6154 0 _0136_
rlabel metal2 17986 6800 17986 6800 0 _0137_
rlabel metal1 18860 5882 18860 5882 0 _0138_
rlabel metal1 19550 6222 19550 6222 0 _0139_
rlabel metal2 20654 5882 20654 5882 0 _0140_
rlabel metal1 20654 5882 20654 5882 0 _0141_
rlabel metal1 24426 5168 24426 5168 0 _0142_
rlabel metal2 30038 4896 30038 4896 0 _0143_
rlabel metal1 30452 3638 30452 3638 0 _0144_
rlabel via1 20562 5355 20562 5355 0 _0145_
rlabel metal2 22494 5440 22494 5440 0 _0146_
rlabel metal1 15824 4590 15824 4590 0 _0147_
rlabel metal1 19136 4998 19136 4998 0 _0148_
rlabel metal2 21390 4522 21390 4522 0 _0149_
rlabel metal1 24518 4726 24518 4726 0 _0150_
rlabel metal1 23782 4556 23782 4556 0 _0151_
rlabel metal2 24058 3978 24058 3978 0 _0152_
rlabel metal1 25990 5168 25990 5168 0 _0153_
rlabel via1 20204 4250 20204 4250 0 _0154_
rlabel metal1 21114 3978 21114 3978 0 _0155_
rlabel metal1 17158 5032 17158 5032 0 _0156_
rlabel metal1 17493 5338 17493 5338 0 _0157_
rlabel metal1 17848 4114 17848 4114 0 _0158_
rlabel metal2 12834 5406 12834 5406 0 _0159_
rlabel metal2 12926 4556 12926 4556 0 _0160_
rlabel metal1 15042 4624 15042 4624 0 _0161_
rlabel metal1 14720 4114 14720 4114 0 _0162_
rlabel metal2 24610 6120 24610 6120 0 _0163_
rlabel metal1 23690 5678 23690 5678 0 _0164_
rlabel metal1 28658 5712 28658 5712 0 _0165_
rlabel metal2 29302 6086 29302 6086 0 _0166_
rlabel metal1 13386 9078 13386 9078 0 _0167_
rlabel metal2 11178 8908 11178 8908 0 _0168_
rlabel metal1 12098 7378 12098 7378 0 _0169_
rlabel metal1 10212 10778 10212 10778 0 _0170_
rlabel metal1 16928 10030 16928 10030 0 _0171_
rlabel metal2 20746 10200 20746 10200 0 _0172_
rlabel metal1 21712 11866 21712 11866 0 _0173_
rlabel metal2 20930 9860 20930 9860 0 _0174_
rlabel metal1 17940 2550 17940 2550 0 _0175_
rlabel metal1 16330 4080 16330 4080 0 _0176_
rlabel metal1 15134 2618 15134 2618 0 _0177_
rlabel metal1 11454 13362 11454 13362 0 _0178_
rlabel metal1 21390 11628 21390 11628 0 _0179_
rlabel metal2 14490 11968 14490 11968 0 _0180_
rlabel metal2 13478 11798 13478 11798 0 _0181_
rlabel metal1 12282 12920 12282 12920 0 _0182_
rlabel metal2 12374 12274 12374 12274 0 _0183_
rlabel metal1 11132 12206 11132 12206 0 _0184_
rlabel metal2 10810 12478 10810 12478 0 _0185_
rlabel metal1 11454 12274 11454 12274 0 _0186_
rlabel metal1 12006 12172 12006 12172 0 _0187_
rlabel metal1 12144 11730 12144 11730 0 _0188_
rlabel metal1 9200 11730 9200 11730 0 _0189_
rlabel metal1 11224 11866 11224 11866 0 _0190_
rlabel metal1 12696 12954 12696 12954 0 _0191_
rlabel metal1 11408 12138 11408 12138 0 _0192_
rlabel metal2 11086 13226 11086 13226 0 _0193_
rlabel metal1 11086 12410 11086 12410 0 _0194_
rlabel metal1 14950 12138 14950 12138 0 _0195_
rlabel metal1 14904 12614 14904 12614 0 _0196_
rlabel metal1 12144 12410 12144 12410 0 _0197_
rlabel metal1 13156 12410 13156 12410 0 _0198_
rlabel metal1 10350 11322 10350 11322 0 _0199_
rlabel metal1 11684 12342 11684 12342 0 _0200_
rlabel viali 12006 11729 12006 11729 0 _0201_
rlabel metal2 12742 12036 12742 12036 0 _0202_
rlabel metal1 16928 12206 16928 12206 0 _0203_
rlabel metal1 23046 12410 23046 12410 0 _0204_
rlabel metal1 30912 13906 30912 13906 0 _0205_
rlabel metal2 27646 11424 27646 11424 0 _0206_
rlabel metal2 36432 6698 36432 6698 0 _0207_
rlabel metal2 41538 5814 41538 5814 0 _0208_
rlabel metal1 36708 6766 36708 6766 0 _0209_
rlabel metal2 36938 6817 36938 6817 0 _0210_
rlabel metal1 33120 9554 33120 9554 0 _0211_
rlabel metal1 34914 9520 34914 9520 0 _0212_
rlabel metal1 35466 9044 35466 9044 0 _0213_
rlabel metal1 34960 8806 34960 8806 0 _0214_
rlabel metal1 35650 8534 35650 8534 0 _0215_
rlabel metal2 35466 6834 35466 6834 0 _0216_
rlabel metal1 37582 4794 37582 4794 0 _0217_
rlabel metal1 38318 5236 38318 5236 0 _0218_
rlabel metal1 38456 4794 38456 4794 0 _0219_
rlabel metal1 34914 5032 34914 5032 0 _0220_
rlabel metal2 43746 6528 43746 6528 0 _0221_
rlabel via1 38790 5270 38790 5270 0 _0222_
rlabel metal1 35880 8942 35880 8942 0 _0223_
rlabel metal1 34730 9588 34730 9588 0 _0224_
rlabel metal1 36478 9486 36478 9486 0 _0225_
rlabel metal2 37582 9724 37582 9724 0 _0226_
rlabel metal1 39744 8330 39744 8330 0 _0227_
rlabel metal2 36754 9792 36754 9792 0 _0228_
rlabel metal1 36570 10098 36570 10098 0 _0229_
rlabel metal1 30728 10234 30728 10234 0 _0230_
rlabel metal2 32246 11356 32246 11356 0 _0231_
rlabel metal1 28842 13260 28842 13260 0 _0232_
rlabel metal1 25576 14450 25576 14450 0 _0233_
rlabel metal1 36662 8602 36662 8602 0 _0234_
rlabel metal2 36386 10982 36386 10982 0 _0235_
rlabel metal1 37444 11118 37444 11118 0 _0236_
rlabel metal1 37122 11866 37122 11866 0 _0237_
rlabel metal1 30820 10166 30820 10166 0 _0238_
rlabel metal1 27186 8942 27186 8942 0 _0239_
rlabel metal1 25806 7888 25806 7888 0 _0240_
rlabel metal1 27002 10064 27002 10064 0 _0241_
rlabel metal1 4968 5202 4968 5202 0 _0242_
rlabel metal1 7912 5678 7912 5678 0 _0243_
rlabel metal1 41906 13804 41906 13804 0 _0244_
rlabel metal1 7958 6766 7958 6766 0 _0245_
rlabel metal2 41446 14756 41446 14756 0 _0246_
rlabel metal2 9338 4624 9338 4624 0 _0247_
rlabel metal2 7038 13668 7038 13668 0 _0248_
rlabel metal2 6210 5389 6210 5389 0 _0249_
rlabel metal2 5658 3978 5658 3978 0 _0250_
rlabel metal2 7222 4012 7222 4012 0 _0251_
rlabel metal1 3312 12954 3312 12954 0 _0252_
rlabel metal2 41814 10234 41814 10234 0 _0253_
rlabel metal2 41446 11764 41446 11764 0 _0254_
rlabel metal1 15594 14518 15594 14518 0 _0255_
rlabel metal2 19550 16116 19550 16116 0 _0256_
rlabel metal2 32062 13974 32062 13974 0 _0257_
rlabel metal2 2162 11951 2162 11951 0 _0258_
rlabel metal1 23644 13294 23644 13294 0 _0259_
rlabel metal1 23000 13158 23000 13158 0 _0260_
rlabel metal1 33534 12682 33534 12682 0 _0261_
rlabel metal1 42642 8296 42642 8296 0 _0262_
rlabel metal2 27278 6596 27278 6596 0 _0263_
rlabel metal2 27370 10115 27370 10115 0 _0264_
rlabel viali 26634 11729 26634 11729 0 _0265_
rlabel metal2 38134 10404 38134 10404 0 _0266_
rlabel metal1 39054 10234 39054 10234 0 _0267_
rlabel metal1 40756 11322 40756 11322 0 _0268_
rlabel metal1 32752 11866 32752 11866 0 _0269_
rlabel metal1 10166 6426 10166 6426 0 _0270_
rlabel metal1 23092 7854 23092 7854 0 _0271_
rlabel metal1 25438 8500 25438 8500 0 _0272_
rlabel metal1 24794 12240 24794 12240 0 _0273_
rlabel metal2 25254 9078 25254 9078 0 _0274_
rlabel metal1 23460 6630 23460 6630 0 _0275_
rlabel metal2 21942 8092 21942 8092 0 _0276_
rlabel metal1 20424 8602 20424 8602 0 _0277_
rlabel metal1 18032 8058 18032 8058 0 _0278_
rlabel metal2 16882 8092 16882 8092 0 _0279_
rlabel metal1 14812 6766 14812 6766 0 _0280_
rlabel metal1 12788 6766 12788 6766 0 _0281_
rlabel metal1 16468 6290 16468 6290 0 _0282_
rlabel metal1 28336 8058 28336 8058 0 _0286_
rlabel metal1 33396 12410 33396 12410 0 _0287_
rlabel metal1 32430 9554 32430 9554 0 _0288_
rlabel metal2 26358 10234 26358 10234 0 _0289_
rlabel metal1 37766 13226 37766 13226 0 _0290_
rlabel metal2 33626 10676 33626 10676 0 _0291_
rlabel metal1 29808 11798 29808 11798 0 _0292_
rlabel metal1 26818 6800 26818 6800 0 _0293_
rlabel metal1 20194 9622 20194 9622 0 _0294_
rlabel metal1 26634 12784 26634 12784 0 _0295_
rlabel metal1 28152 10030 28152 10030 0 _0296_
rlabel metal1 39284 11254 39284 11254 0 _0297_
rlabel metal1 34454 10030 34454 10030 0 _0298_
rlabel metal1 36524 12818 36524 12818 0 _0299_
rlabel metal2 20378 9146 20378 9146 0 _0300_
rlabel metal1 22080 12206 22080 12206 0 _0301_
rlabel metal1 20838 11288 20838 11288 0 _0302_
rlabel viali 15594 10644 15594 10644 0 _0303_
rlabel metal1 14766 10030 14766 10030 0 _0304_
rlabel metal1 9660 4114 9660 4114 0 _0305_
rlabel metal1 11500 6766 11500 6766 0 _0306_
rlabel metal1 10166 8058 10166 8058 0 _0307_
rlabel metal1 13478 7514 13478 7514 0 _0308_
rlabel metal1 36938 14042 36938 14042 0 _0309_
rlabel metal1 35696 13906 35696 13906 0 _0310_
rlabel metal1 34086 14518 34086 14518 0 _0311_
rlabel metal2 33626 14790 33626 14790 0 _0312_
rlabel metal2 35742 15844 35742 15844 0 _0313_
rlabel metal2 36662 15436 36662 15436 0 _0314_
rlabel metal1 25898 14246 25898 14246 0 _0315_
rlabel metal1 25162 14586 25162 14586 0 _0316_
rlabel metal1 22586 13294 22586 13294 0 _0317_
rlabel metal2 22218 13940 22218 13940 0 _0318_
rlabel metal1 20148 13294 20148 13294 0 _0319_
rlabel metal1 19412 13498 19412 13498 0 _0320_
rlabel metal1 19044 14246 19044 14246 0 _0321_
rlabel metal1 17940 14382 17940 14382 0 _0322_
rlabel metal2 37030 7514 37030 7514 0 _0323_
rlabel metal1 33350 7854 33350 7854 0 _0324_
rlabel metal1 40020 8466 40020 8466 0 _0325_
rlabel metal2 39422 8772 39422 8772 0 _0326_
rlabel metal2 42918 9826 42918 9826 0 _0327_
rlabel metal1 42826 9996 42826 9996 0 _0328_
rlabel metal2 42826 10438 42826 10438 0 _0329_
rlabel metal2 42642 9452 42642 9452 0 _0330_
rlabel metal1 40158 9146 40158 9146 0 _0331_
rlabel metal1 40020 10234 40020 10234 0 _0332_
rlabel metal2 42918 8976 42918 8976 0 _0333_
rlabel metal1 42504 8534 42504 8534 0 _0334_
rlabel metal1 42872 7854 42872 7854 0 _0335_
rlabel metal1 41124 6358 41124 6358 0 _0336_
rlabel metal1 42826 6256 42826 6256 0 _0337_
rlabel metal1 34040 6290 34040 6290 0 _0338_
rlabel metal1 35144 6766 35144 6766 0 _0339_
rlabel metal1 34224 5882 34224 5882 0 _0340_
rlabel metal2 34362 6630 34362 6630 0 _0341_
rlabel metal1 35972 6222 35972 6222 0 _0342_
rlabel metal1 35650 6630 35650 6630 0 _0343_
rlabel metal1 35696 4590 35696 4590 0 _0344_
rlabel metal1 33810 6358 33810 6358 0 _0345_
rlabel metal1 34178 6256 34178 6256 0 _0346_
rlabel metal1 33304 5202 33304 5202 0 _0347_
rlabel metal2 31326 9078 31326 9078 0 _0348_
rlabel metal1 31096 7514 31096 7514 0 _0349_
rlabel metal1 30728 6290 30728 6290 0 _0350_
rlabel metal2 33810 6970 33810 6970 0 _0351_
rlabel metal1 33442 6630 33442 6630 0 _0352_
rlabel metal2 32798 7174 32798 7174 0 _0353_
rlabel metal2 32338 6732 32338 6732 0 _0354_
rlabel metal1 42136 7310 42136 7310 0 _0355_
rlabel metal1 42642 7412 42642 7412 0 _0356_
rlabel metal2 40158 6970 40158 6970 0 _0357_
rlabel metal2 38594 7990 38594 7990 0 _0358_
rlabel metal1 36202 7854 36202 7854 0 _0359_
rlabel metal1 39284 7514 39284 7514 0 _0360_
rlabel metal2 41630 7548 41630 7548 0 _0361_
rlabel metal1 35972 7514 35972 7514 0 _0362_
rlabel metal1 35374 8058 35374 8058 0 _0363_
rlabel metal2 37398 8296 37398 8296 0 _0364_
rlabel metal2 38042 8092 38042 8092 0 _0365_
rlabel metal1 28934 9486 28934 9486 0 _0366_
rlabel metal1 30774 14586 30774 14586 0 _0367_
rlabel metal2 30222 14518 30222 14518 0 _0368_
rlabel metal1 39606 14382 39606 14382 0 _0369_
rlabel metal1 20424 14994 20424 14994 0 _0370_
rlabel metal1 18814 10234 18814 10234 0 _0371_
rlabel metal1 17572 11254 17572 11254 0 _0372_
rlabel metal1 17756 11322 17756 11322 0 _0373_
rlabel metal1 6394 6766 6394 6766 0 _0374_
rlabel metal2 7958 11322 7958 11322 0 _0375_
rlabel metal2 7314 7548 7314 7548 0 _0376_
rlabel metal1 3634 10234 3634 10234 0 _0377_
rlabel metal1 3496 7378 3496 7378 0 _0378_
rlabel metal1 4278 5066 4278 5066 0 _0379_
rlabel metal1 2852 7718 2852 7718 0 _0380_
rlabel metal1 3542 10030 3542 10030 0 _0381_
rlabel metal2 8510 5134 8510 5134 0 _0382_
rlabel metal1 10304 4590 10304 4590 0 _0383_
rlabel metal1 10442 7174 10442 7174 0 _0384_
rlabel metal1 24702 12376 24702 12376 0 _0385_
rlabel via1 5290 12886 5290 12886 0 _0386_
rlabel metal2 12742 13498 12742 13498 0 _0387_
rlabel metal1 14996 13498 14996 13498 0 _0388_
rlabel metal1 11316 13294 11316 13294 0 _0389_
rlabel metal1 15548 13498 15548 13498 0 _0390_
rlabel metal1 8326 13974 8326 13974 0 _0391_
rlabel metal1 11592 13702 11592 13702 0 _0392_
rlabel metal2 12282 14212 12282 14212 0 _0393_
rlabel via1 6034 13226 6034 13226 0 _0394_
rlabel metal1 7912 13498 7912 13498 0 _0395_
rlabel metal1 7314 13430 7314 13430 0 _0396_
rlabel metal1 5842 14416 5842 14416 0 _0397_
rlabel metal1 5842 14042 5842 14042 0 _0398_
rlabel metal2 5658 14790 5658 14790 0 _0399_
rlabel metal2 4370 13566 4370 13566 0 _0400_
rlabel metal1 5014 14042 5014 14042 0 _0401_
rlabel metal1 3450 13396 3450 13396 0 _0402_
rlabel metal2 5842 12172 5842 12172 0 _0403_
rlabel metal1 6410 12886 6410 12886 0 _0404_
rlabel metal1 5612 12818 5612 12818 0 _0405_
rlabel metal1 5152 12206 5152 12206 0 _0406_
rlabel metal1 5520 11866 5520 11866 0 _0407_
rlabel metal1 3450 12172 3450 12172 0 _0408_
rlabel metal2 27646 6086 27646 6086 0 _0409_
rlabel metal2 26082 6324 26082 6324 0 _0410_
rlabel metal1 15410 4794 15410 4794 0 _0411_
rlabel metal2 12742 5372 12742 5372 0 _0412_
rlabel metal2 19642 3706 19642 3706 0 _0413_
rlabel metal2 20654 3706 20654 3706 0 _0414_
rlabel metal2 27002 3706 27002 3706 0 _0415_
rlabel metal1 25484 3706 25484 3706 0 _0416_
rlabel metal1 28750 4114 28750 4114 0 _0417_
rlabel metal1 34270 8908 34270 8908 0 _0418_
rlabel metal1 39054 11152 39054 11152 0 _0419_
rlabel metal2 26358 9350 26358 9350 0 active
rlabel metal1 1472 17170 1472 17170 0 active_select[0]
rlabel metal2 43838 1588 43838 1588 0 active_select[1]
rlabel metal2 45126 1894 45126 1894 0 active_select[2]
rlabel metal2 36754 840 36754 840 0 active_select[3]
rlabel metal1 31096 17170 31096 17170 0 active_select[4]
rlabel metal2 25806 1588 25806 1588 0 active_select[5]
rlabel via2 44390 7837 44390 7837 0 active_select[6]
rlabel metal3 820 17068 820 17068 0 active_select[7]
rlabel metal2 3266 18234 3266 18234 0 active_select[8]
rlabel metal2 30590 9146 30590 9146 0 aio_input_reg\[0\]
rlabel metal1 35374 14042 35374 14042 0 aio_input_reg\[1\]
rlabel metal1 33212 14314 33212 14314 0 aio_input_reg\[2\]
rlabel metal1 41538 14586 41538 14586 0 aio_input_reg\[3\]
rlabel metal1 24932 14382 24932 14382 0 aio_input_reg\[4\]
rlabel metal1 21390 12682 21390 12682 0 aio_input_reg\[5\]
rlabel metal2 18906 13056 18906 13056 0 aio_input_reg\[6\]
rlabel metal1 18722 13498 18722 13498 0 aio_input_reg\[7\]
rlabel metal1 24518 13804 24518 13804 0 aio_input_sh
rlabel metal2 37490 11288 37490 11288 0 aio_input_shift\[0\]
rlabel metal2 37858 14144 37858 14144 0 aio_input_shift\[1\]
rlabel metal1 36570 14858 36570 14858 0 aio_input_shift\[2\]
rlabel metal1 26726 14518 26726 14518 0 aio_input_shift\[3\]
rlabel metal2 26634 14586 26634 14586 0 aio_input_shift\[4\]
rlabel metal1 23828 14042 23828 14042 0 aio_input_shift\[5\]
rlabel metal2 19918 14144 19918 14144 0 aio_input_shift\[6\]
rlabel metal1 18890 15062 18890 15062 0 aio_input_shift\[7\]
rlabel metal2 29210 9350 29210 9350 0 aio_input_sync\[0\]
rlabel metal1 29946 14416 29946 14416 0 aio_input_sync\[1\]
rlabel metal2 30038 14348 30038 14348 0 aio_input_sync\[2\]
rlabel metal2 40158 14518 40158 14518 0 aio_input_sync\[3\]
rlabel metal1 17066 15130 17066 15130 0 aio_input_sync\[4\]
rlabel metal1 18078 9146 18078 9146 0 aio_input_sync\[5\]
rlabel metal2 16330 10234 16330 10234 0 aio_input_sync\[6\]
rlabel metal2 18262 10234 18262 10234 0 aio_input_sync\[7\]
rlabel metal1 4876 5134 4876 5134 0 aio_output_cap
rlabel metal2 5658 9248 5658 9248 0 aio_output_reg\[0\]
rlabel metal2 41814 12801 41814 12801 0 aio_output_reg\[1\]
rlabel metal1 9108 6290 9108 6290 0 aio_output_reg\[2\]
rlabel metal1 5152 10506 5152 10506 0 aio_output_reg\[3\]
rlabel metal1 5290 6426 5290 6426 0 aio_output_reg\[4\]
rlabel metal2 4370 5882 4370 5882 0 aio_output_reg\[5\]
rlabel metal1 5336 5882 5336 5882 0 aio_output_reg\[6\]
rlabel metal2 3450 12070 3450 12070 0 aio_output_reg\[7\]
rlabel metal2 7958 9758 7958 9758 0 aio_output_shift\[0\]
rlabel metal1 7820 9418 7820 9418 0 aio_output_shift\[1\]
rlabel metal1 4646 8534 4646 8534 0 aio_output_shift\[2\]
rlabel metal1 4365 8534 4365 8534 0 aio_output_shift\[3\]
rlabel metal1 4825 6766 4825 6766 0 aio_output_shift\[4\]
rlabel metal1 5382 6664 5382 6664 0 aio_output_shift\[5\]
rlabel metal2 3174 8738 3174 8738 0 aio_output_shift\[6\]
rlabel metal2 3910 10234 3910 10234 0 aio_output_shift\[7\]
rlabel metal1 40986 8398 40986 8398 0 bit_cnt\[0\]
rlabel metal1 40112 10710 40112 10710 0 bit_cnt\[1\]
rlabel metal2 40526 10098 40526 10098 0 bit_cnt\[2\]
rlabel metal1 42780 9554 42780 9554 0 bit_cnt\[3\]
rlabel metal2 33534 2098 33534 2098 0 clk
rlabel metal1 25484 9010 25484 9010 0 clk_divider_I.active
rlabel metal1 36708 11118 36708 11118 0 clk_divider_I.ce
rlabel metal1 24702 6800 24702 6800 0 clk_divider_I.compare\[0\]
rlabel metal1 21114 7242 21114 7242 0 clk_divider_I.compare\[1\]
rlabel metal2 21666 6834 21666 6834 0 clk_divider_I.compare\[2\]
rlabel metal1 18400 7854 18400 7854 0 clk_divider_I.compare\[3\]
rlabel metal2 16238 8262 16238 8262 0 clk_divider_I.compare\[4\]
rlabel metal1 15594 5882 15594 5882 0 clk_divider_I.compare\[5\]
rlabel metal2 19274 5967 19274 5967 0 clk_divider_I.compare\[6\]
rlabel metal1 18400 5678 18400 5678 0 clk_divider_I.compare\[7\]
rlabel metal2 29854 5610 29854 5610 0 clk_divider_I.counter\[0\]
rlabel metal1 24840 5678 24840 5678 0 clk_divider_I.counter\[1\]
rlabel metal1 15778 5168 15778 5168 0 clk_divider_I.counter\[2\]
rlabel metal1 18170 5236 18170 5236 0 clk_divider_I.counter\[3\]
rlabel via1 18262 5746 18262 5746 0 clk_divider_I.counter\[4\]
rlabel metal1 21482 5168 21482 5168 0 clk_divider_I.counter\[5\]
rlabel metal2 27370 4998 27370 4998 0 clk_divider_I.counter\[6\]
rlabel metal2 24058 4964 24058 4964 0 clk_divider_I.counter\[7\]
rlabel metal1 20102 4114 20102 4114 0 clk_divider_I.reset
rlabel metal2 15686 7140 15686 7140 0 clk_divider_I.set_now
rlabel metal1 12006 15572 12006 15572 0 clk_divider_I.set_sync\[0\]
rlabel metal1 18630 14824 18630 14824 0 clk_divider_I.set_sync\[1\]
rlabel metal1 13156 10642 13156 10642 0 clknet_0_clk
rlabel metal1 5428 7854 5428 7854 0 clknet_0_scan_clk_in
rlabel metal1 3036 6766 3036 6766 0 clknet_1_0__leaf_scan_clk_in
rlabel metal1 6440 8398 6440 8398 0 clknet_1_1__leaf_scan_clk_in
rlabel metal1 4186 5678 4186 5678 0 clknet_3_0__leaf_clk
rlabel metal1 15410 2448 15410 2448 0 clknet_3_1__leaf_clk
rlabel metal2 6578 14144 6578 14144 0 clknet_3_2__leaf_clk
rlabel metal1 11914 15028 11914 15028 0 clknet_3_3__leaf_clk
rlabel metal1 28152 5134 28152 5134 0 clknet_3_4__leaf_clk
rlabel metal2 40526 8432 40526 8432 0 clknet_3_5__leaf_clk
rlabel metal1 24886 15028 24886 15028 0 clknet_3_6__leaf_clk
rlabel metal1 38778 13940 38778 13940 0 clknet_3_7__leaf_clk
rlabel metal2 27094 1554 27094 1554 0 driver_sel[0]
rlabel metal1 874 16558 874 16558 0 driver_sel[1]
rlabel metal2 32246 1554 32246 1554 0 inputs[0]
rlabel metal1 11454 17238 11454 17238 0 inputs[1]
rlabel metal1 32292 17170 32292 17170 0 inputs[2]
rlabel metal1 38778 17238 38778 17238 0 inputs[3]
rlabel metal1 4600 17170 4600 17170 0 inputs[4]
rlabel metal2 12926 1588 12926 1588 0 inputs[5]
rlabel metal3 820 4828 820 4828 0 inputs[6]
rlabel metal2 41906 1554 41906 1554 0 inputs[7]
rlabel metal2 41906 11356 41906 11356 0 int_scan_clk_out
rlabel metal1 20194 15130 20194 15130 0 int_scan_data_out
rlabel metal1 24978 13158 24978 13158 0 int_scan_latch_en
rlabel metal2 31510 13056 31510 13056 0 int_scan_select
rlabel metal2 44390 8687 44390 8687 0 la_scan_clk_in
rlabel metal3 820 8228 820 8228 0 la_scan_data_in
rlabel metal3 45180 14348 45180 14348 0 la_scan_data_out
rlabel metal1 24334 17170 24334 17170 0 la_scan_latch_en
rlabel metal2 35098 18122 35098 18122 0 la_scan_select
rlabel metal2 1794 13209 1794 13209 0 net1
rlabel metal1 23874 14484 23874 14484 0 net10
rlabel metal1 3542 16626 3542 16626 0 net11
rlabel metal1 23414 9894 23414 9894 0 net12
rlabel metal1 23782 14348 23782 14348 0 net13
rlabel metal1 28280 14994 28280 14994 0 net14
rlabel via2 23690 14331 23690 14331 0 net15
rlabel metal1 7912 17102 7912 17102 0 net16
rlabel metal1 12880 2618 12880 2618 0 net17
rlabel metal2 1886 4930 1886 4930 0 net18
rlabel metal1 22057 2618 22057 2618 0 net19
rlabel metal2 43930 4114 43930 4114 0 net2
rlabel metal2 44206 9010 44206 9010 0 net20
rlabel metal1 4255 7990 4255 7990 0 net21
rlabel metal1 24196 16966 24196 16966 0 net22
rlabel metal1 33166 14994 33166 14994 0 net23
rlabel metal1 17802 2380 17802 2380 0 net24
rlabel via2 41722 13957 41722 13957 0 net25
rlabel metal1 10028 16966 10028 16966 0 net26
rlabel metal2 14858 3264 14858 3264 0 net27
rlabel metal1 13064 17170 13064 17170 0 net28
rlabel metal2 16146 1656 16146 1656 0 net29
rlabel metal2 44206 3910 44206 3910 0 net3
rlabel metal1 44528 3502 44528 3502 0 net30
rlabel metal1 35604 17170 35604 17170 0 net31
rlabel metal1 44758 16762 44758 16762 0 net32
rlabel metal1 19504 17170 19504 17170 0 net33
rlabel metal2 4554 1588 4554 1588 0 net34
rlabel metal2 1334 1588 1334 1588 0 net35
rlabel metal2 43470 17612 43470 17612 0 net36
rlabel metal3 820 13668 820 13668 0 net37
rlabel metal2 20654 823 20654 823 0 net38
rlabel metal1 44712 12614 44712 12614 0 net39
rlabel metal1 37168 4590 37168 4590 0 net4
rlabel metal2 44390 15793 44390 15793 0 net40
rlabel metal2 29026 1588 29026 1588 0 net41
rlabel metal1 37536 17170 37536 17170 0 net42
rlabel metal2 3266 840 3266 840 0 net43
rlabel metal1 7912 17170 7912 17170 0 net44
rlabel metal2 10994 823 10994 823 0 net45
rlabel metal1 43976 17170 43976 17170 0 net46
rlabel metal1 44712 11118 44712 11118 0 net47
rlabel metal2 42826 18122 42826 18122 0 net48
rlabel metal2 7774 1588 7774 1588 0 net49
rlabel metal1 31188 16966 31188 16966 0 net5
rlabel metal2 23874 1588 23874 1588 0 net50
rlabel metal2 39974 823 39974 823 0 net51
rlabel metal1 6624 17170 6624 17170 0 net52
rlabel metal2 19366 1588 19366 1588 0 net53
rlabel metal1 14352 17170 14352 17170 0 net54
rlabel metal2 30314 823 30314 823 0 net55
rlabel metal1 25944 17170 25944 17170 0 net56
rlabel metal2 38686 1588 38686 1588 0 net57
rlabel metal1 1380 5882 1380 5882 0 net58
rlabel metal3 820 1428 820 1428 0 net59
rlabel metal1 28290 2278 28290 2278 0 net6
rlabel metal1 22724 17170 22724 17170 0 net60
rlabel metal1 29486 17170 29486 17170 0 net61
rlabel metal3 820 3468 820 3468 0 net62
rlabel metal2 46 1622 46 1622 0 net63
rlabel metal3 866 18428 866 18428 0 net64
rlabel metal1 27876 17170 27876 17170 0 net65
rlabel metal2 13662 3196 13662 3196 0 net66
rlabel metal1 17342 3026 17342 3026 0 net67
rlabel metal1 15778 2414 15778 2414 0 net68
rlabel metal2 12650 15164 12650 15164 0 net69
rlabel metal1 43838 7718 43838 7718 0 net7
rlabel metal1 3036 9622 3036 9622 0 net8
rlabel metal1 3542 17034 3542 17034 0 net9
rlabel metal1 9660 6630 9660 6630 0 outputs[0]
rlabel metal1 44528 17510 44528 17510 0 outputs[1]
rlabel metal2 35466 1860 35466 1860 0 outputs[2]
rlabel metal2 17250 16915 17250 16915 0 outputs[3]
rlabel metal1 44344 5134 44344 5134 0 outputs[4]
rlabel metal2 6486 1231 6486 1231 0 outputs[5]
rlabel metal2 9706 1860 9706 1860 0 outputs[6]
rlabel metal3 866 15028 866 15028 0 outputs[7]
rlabel metal2 41722 5372 41722 5372 0 proj_cnt\[0\]
rlabel metal2 36570 6324 36570 6324 0 proj_cnt\[1\]
rlabel metal1 37352 5202 37352 5202 0 proj_cnt\[2\]
rlabel metal2 35006 5542 35006 5542 0 proj_cnt\[3\]
rlabel metal1 31878 6868 31878 6868 0 proj_cnt\[4\]
rlabel metal1 30774 6630 30774 6630 0 proj_cnt\[5\]
rlabel metal1 43056 6630 43056 6630 0 proj_cnt\[6\]
rlabel metal2 36294 7820 36294 7820 0 proj_cnt\[7\]
rlabel metal2 36570 8228 36570 8228 0 proj_cnt\[8\]
rlabel via2 41446 5219 41446 5219 0 ready
rlabel metal2 17434 1588 17434 1588 0 reset
rlabel via1 16261 3026 16261 3026 0 rst_shift\[0\]
rlabel metal2 18078 3230 18078 3230 0 rst_shift\[1\]
rlabel metal3 2384 11628 2384 11628 0 scan_clk_in
rlabel metal2 41538 14144 41538 14144 0 scan_clk_out
rlabel metal2 16882 18122 16882 18122 0 scan_data_in
rlabel metal1 20792 16558 20792 16558 0 scan_data_out
rlabel metal1 23000 2958 23000 2958 0 scan_latch_en
rlabel metal3 820 10268 820 10268 0 scan_select
rlabel metal1 9844 17170 9844 17170 0 set_clk_div
rlabel metal2 41446 3213 41446 3213 0 slow_clk
rlabel metal1 41906 10200 41906 10200 0 state\[0\]
rlabel metal2 36018 11390 36018 11390 0 state\[12\]
rlabel metal1 37904 12070 37904 12070 0 state\[13\]
rlabel metal2 32522 11900 32522 11900 0 state\[1\]
rlabel metal2 31602 10642 31602 10642 0 state\[2\]
rlabel metal1 21735 10574 21735 10574 0 state\[3\]
rlabel metal1 38824 12410 38824 12410 0 state\[4\]
rlabel metal2 35190 10268 35190 10268 0 state\[5\]
rlabel metal1 29762 12648 29762 12648 0 state\[6\]
rlabel metal1 17158 12172 17158 12172 0 state\[8\]
rlabel metal1 25640 13226 25640 13226 0 state\[9\]
rlabel metal1 21643 10642 21643 10642 0 ws_cfg\[0\]
rlabel metal2 21206 11220 21206 11220 0 ws_cfg\[1\]
rlabel metal1 18170 11696 18170 11696 0 ws_cfg\[2\]
rlabel metal1 15456 11730 15456 11730 0 ws_cfg\[3\]
rlabel metal2 11270 11356 11270 11356 0 ws_cfg\[4\]
rlabel metal1 11730 10642 11730 10642 0 ws_cfg\[5\]
rlabel metal1 12236 10778 12236 10778 0 ws_cfg\[6\]
rlabel metal2 13202 10540 13202 10540 0 ws_cfg\[7\]
rlabel metal2 14490 13838 14490 13838 0 ws_cnt\[0\]
rlabel metal1 14628 14042 14628 14042 0 ws_cnt\[1\]
rlabel metal1 13156 14382 13156 14382 0 ws_cnt\[2\]
rlabel metal1 9016 13906 9016 13906 0 ws_cnt\[3\]
rlabel metal1 5796 13906 5796 13906 0 ws_cnt\[4\]
rlabel metal1 6440 13498 6440 13498 0 ws_cnt\[5\]
rlabel metal1 5934 12648 5934 12648 0 ws_cnt\[6\]
rlabel metal1 5750 11764 5750 11764 0 ws_cnt\[7\]
rlabel metal1 11914 7956 11914 7956 0 ws_set_now
rlabel metal1 9062 5134 9062 5134 0 ws_set_sync\[0\]
rlabel metal1 10580 6154 10580 6154 0 ws_set_sync\[1\]
rlabel metal1 10396 6358 10396 6358 0 ws_set_sync\[2\]
<< properties >>
string FIXED_BBOX 0 0 46000 20000
<< end >>
