module MichaelBell_6bit_fifo (vccd1,
    vssd1,
    io_in,
    io_out);
 input vccd1;
 input vssd1;
 input [7:0] io_in;
 output [7:0] io_out;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire _203_;
 wire _204_;
 wire _205_;
 wire _206_;
 wire _207_;
 wire _208_;
 wire _209_;
 wire _210_;
 wire _211_;
 wire _212_;
 wire _213_;
 wire _214_;
 wire _215_;
 wire _216_;
 wire _217_;
 wire _218_;
 wire _219_;
 wire _220_;
 wire _221_;
 wire _222_;
 wire _223_;
 wire _224_;
 wire _225_;
 wire _226_;
 wire _227_;
 wire _228_;
 wire _229_;
 wire _230_;
 wire _231_;
 wire _232_;
 wire _233_;
 wire _234_;
 wire _235_;
 wire _236_;
 wire _237_;
 wire _238_;
 wire _239_;
 wire _240_;
 wire _241_;
 wire _242_;
 wire _243_;
 wire _244_;
 wire _245_;
 wire _246_;
 wire _247_;
 wire _248_;
 wire _249_;
 wire _250_;
 wire _251_;
 wire \data_in_buffer[0].A ;
 wire \data_in_buffer[0].X ;
 wire \data_in_buffer[0].b[0] ;
 wire \data_in_buffer[0].genblk1[0].mid ;
 wire \data_in_buffer[0].genblk1[1].mid ;
 wire \data_in_buffer[1].A ;
 wire \data_in_buffer[1].X ;
 wire \data_in_buffer[1].b[0] ;
 wire \data_in_buffer[1].genblk1[0].mid ;
 wire \data_in_buffer[1].genblk1[1].mid ;
 wire \data_in_buffer[2].A ;
 wire \data_in_buffer[2].X ;
 wire \data_in_buffer[2].b[0] ;
 wire \data_in_buffer[2].genblk1[0].mid ;
 wire \data_in_buffer[2].genblk1[1].mid ;
 wire \data_in_buffer[3].A ;
 wire \data_in_buffer[3].X ;
 wire \data_in_buffer[3].b[0] ;
 wire \data_in_buffer[3].genblk1[0].mid ;
 wire \data_in_buffer[3].genblk1[1].mid ;
 wire \data_in_buffer[4].A ;
 wire \data_in_buffer[4].X ;
 wire \data_in_buffer[4].b[0] ;
 wire \data_in_buffer[4].genblk1[0].mid ;
 wire \data_in_buffer[4].genblk1[1].mid ;
 wire \data_in_buffer[5].A ;
 wire \data_in_buffer[5].X ;
 wire \data_in_buffer[5].b[0] ;
 wire \data_in_buffer[5].genblk1[0].mid ;
 wire \data_in_buffer[5].genblk1[1].mid ;
 wire \f_fifo.data_in[0] ;
 wire \f_fifo.data_in[1] ;
 wire \f_fifo.data_in[2] ;
 wire \f_fifo.data_in[3] ;
 wire \f_fifo.data_in[4] ;
 wire \f_fifo.data_in[5] ;
 wire \f_fifo.empty_n ;
 wire \f_fifo.fifo_data[0][0] ;
 wire \f_fifo.fifo_data[0][1] ;
 wire \f_fifo.fifo_data[0][2] ;
 wire \f_fifo.fifo_data[0][3] ;
 wire \f_fifo.fifo_data[0][4] ;
 wire \f_fifo.fifo_data[0][5] ;
 wire \f_fifo.fifo_data[1][0] ;
 wire \f_fifo.fifo_data[1][1] ;
 wire \f_fifo.fifo_data[1][2] ;
 wire \f_fifo.fifo_data[1][3] ;
 wire \f_fifo.fifo_data[1][4] ;
 wire \f_fifo.fifo_data[1][5] ;
 wire \f_fifo.fifo_data[2][0] ;
 wire \f_fifo.fifo_data[2][1] ;
 wire \f_fifo.fifo_data[2][2] ;
 wire \f_fifo.fifo_data[2][3] ;
 wire \f_fifo.fifo_data[2][4] ;
 wire \f_fifo.fifo_data[2][5] ;
 wire \f_fifo.fifo_data[3][0] ;
 wire \f_fifo.fifo_data[3][1] ;
 wire \f_fifo.fifo_data[3][2] ;
 wire \f_fifo.fifo_data[3][3] ;
 wire \f_fifo.fifo_data[3][4] ;
 wire \f_fifo.fifo_data[3][5] ;
 wire \f_fifo.read_addr[0] ;
 wire \f_fifo.read_addr[1] ;
 wire \f_fifo.reset_n ;
 wire \f_fifo.write_addr[0] ;
 wire \f_fifo.write_addr[1] ;
 wire \l_fifo.genblk1[0].entry.empty ;
 wire \l_fifo.genblk1[0].entry.input_buf[0].A ;
 wire \l_fifo.genblk1[0].entry.input_buf[0].X ;
 wire \l_fifo.genblk1[0].entry.input_buf[0].genblk1[0].mid ;
 wire \l_fifo.genblk1[0].entry.input_buf[1].A ;
 wire \l_fifo.genblk1[0].entry.input_buf[1].X ;
 wire \l_fifo.genblk1[0].entry.input_buf[1].genblk1[0].mid ;
 wire \l_fifo.genblk1[0].entry.input_buf[2].A ;
 wire \l_fifo.genblk1[0].entry.input_buf[2].X ;
 wire \l_fifo.genblk1[0].entry.input_buf[2].genblk1[0].mid ;
 wire \l_fifo.genblk1[0].entry.input_buf[3].A ;
 wire \l_fifo.genblk1[0].entry.input_buf[3].X ;
 wire \l_fifo.genblk1[0].entry.input_buf[3].genblk1[0].mid ;
 wire \l_fifo.genblk1[0].entry.input_buf[4].A ;
 wire \l_fifo.genblk1[0].entry.input_buf[4].X ;
 wire \l_fifo.genblk1[0].entry.input_buf[4].genblk1[0].mid ;
 wire \l_fifo.genblk1[0].entry.input_buf[5].A ;
 wire \l_fifo.genblk1[0].entry.input_buf[5].X ;
 wire \l_fifo.genblk1[0].entry.input_buf[5].genblk1[0].mid ;
 wire \l_fifo.genblk1[10].entry.empty ;
 wire \l_fifo.genblk1[10].entry.input_buf[0].A ;
 wire \l_fifo.genblk1[10].entry.input_buf[0].X ;
 wire \l_fifo.genblk1[10].entry.input_buf[0].genblk1[0].mid ;
 wire \l_fifo.genblk1[10].entry.input_buf[1].A ;
 wire \l_fifo.genblk1[10].entry.input_buf[1].X ;
 wire \l_fifo.genblk1[10].entry.input_buf[1].genblk1[0].mid ;
 wire \l_fifo.genblk1[10].entry.input_buf[2].A ;
 wire \l_fifo.genblk1[10].entry.input_buf[2].X ;
 wire \l_fifo.genblk1[10].entry.input_buf[2].genblk1[0].mid ;
 wire \l_fifo.genblk1[10].entry.input_buf[3].A ;
 wire \l_fifo.genblk1[10].entry.input_buf[3].X ;
 wire \l_fifo.genblk1[10].entry.input_buf[3].genblk1[0].mid ;
 wire \l_fifo.genblk1[10].entry.input_buf[4].A ;
 wire \l_fifo.genblk1[10].entry.input_buf[4].X ;
 wire \l_fifo.genblk1[10].entry.input_buf[4].genblk1[0].mid ;
 wire \l_fifo.genblk1[10].entry.input_buf[5].A ;
 wire \l_fifo.genblk1[10].entry.input_buf[5].X ;
 wire \l_fifo.genblk1[10].entry.input_buf[5].genblk1[0].mid ;
 wire \l_fifo.genblk1[10].entry.next_is_empty ;
 wire \l_fifo.genblk1[11].entry.empty ;
 wire \l_fifo.genblk1[11].entry.input_buf[0].A ;
 wire \l_fifo.genblk1[11].entry.input_buf[0].X ;
 wire \l_fifo.genblk1[11].entry.input_buf[0].genblk1[0].mid ;
 wire \l_fifo.genblk1[11].entry.input_buf[1].A ;
 wire \l_fifo.genblk1[11].entry.input_buf[1].X ;
 wire \l_fifo.genblk1[11].entry.input_buf[1].genblk1[0].mid ;
 wire \l_fifo.genblk1[11].entry.input_buf[2].A ;
 wire \l_fifo.genblk1[11].entry.input_buf[2].X ;
 wire \l_fifo.genblk1[11].entry.input_buf[2].genblk1[0].mid ;
 wire \l_fifo.genblk1[11].entry.input_buf[3].A ;
 wire \l_fifo.genblk1[11].entry.input_buf[3].X ;
 wire \l_fifo.genblk1[11].entry.input_buf[3].genblk1[0].mid ;
 wire \l_fifo.genblk1[11].entry.input_buf[4].A ;
 wire \l_fifo.genblk1[11].entry.input_buf[4].X ;
 wire \l_fifo.genblk1[11].entry.input_buf[4].genblk1[0].mid ;
 wire \l_fifo.genblk1[11].entry.input_buf[5].A ;
 wire \l_fifo.genblk1[11].entry.input_buf[5].X ;
 wire \l_fifo.genblk1[11].entry.input_buf[5].genblk1[0].mid ;
 wire \l_fifo.genblk1[12].entry.empty ;
 wire \l_fifo.genblk1[12].entry.input_buf[0].A ;
 wire \l_fifo.genblk1[12].entry.input_buf[0].X ;
 wire \l_fifo.genblk1[12].entry.input_buf[0].genblk1[0].mid ;
 wire \l_fifo.genblk1[12].entry.input_buf[1].A ;
 wire \l_fifo.genblk1[12].entry.input_buf[1].X ;
 wire \l_fifo.genblk1[12].entry.input_buf[1].genblk1[0].mid ;
 wire \l_fifo.genblk1[12].entry.input_buf[2].A ;
 wire \l_fifo.genblk1[12].entry.input_buf[2].X ;
 wire \l_fifo.genblk1[12].entry.input_buf[2].genblk1[0].mid ;
 wire \l_fifo.genblk1[12].entry.input_buf[3].A ;
 wire \l_fifo.genblk1[12].entry.input_buf[3].X ;
 wire \l_fifo.genblk1[12].entry.input_buf[3].genblk1[0].mid ;
 wire \l_fifo.genblk1[12].entry.input_buf[4].A ;
 wire \l_fifo.genblk1[12].entry.input_buf[4].X ;
 wire \l_fifo.genblk1[12].entry.input_buf[4].genblk1[0].mid ;
 wire \l_fifo.genblk1[12].entry.input_buf[5].A ;
 wire \l_fifo.genblk1[12].entry.input_buf[5].X ;
 wire \l_fifo.genblk1[12].entry.input_buf[5].genblk1[0].mid ;
 wire \l_fifo.genblk1[13].entry.empty ;
 wire \l_fifo.genblk1[13].entry.input_buf[0].A ;
 wire \l_fifo.genblk1[13].entry.input_buf[0].X ;
 wire \l_fifo.genblk1[13].entry.input_buf[0].genblk1[0].mid ;
 wire \l_fifo.genblk1[13].entry.input_buf[1].A ;
 wire \l_fifo.genblk1[13].entry.input_buf[1].X ;
 wire \l_fifo.genblk1[13].entry.input_buf[1].genblk1[0].mid ;
 wire \l_fifo.genblk1[13].entry.input_buf[2].A ;
 wire \l_fifo.genblk1[13].entry.input_buf[2].X ;
 wire \l_fifo.genblk1[13].entry.input_buf[2].genblk1[0].mid ;
 wire \l_fifo.genblk1[13].entry.input_buf[3].A ;
 wire \l_fifo.genblk1[13].entry.input_buf[3].X ;
 wire \l_fifo.genblk1[13].entry.input_buf[3].genblk1[0].mid ;
 wire \l_fifo.genblk1[13].entry.input_buf[4].A ;
 wire \l_fifo.genblk1[13].entry.input_buf[4].X ;
 wire \l_fifo.genblk1[13].entry.input_buf[4].genblk1[0].mid ;
 wire \l_fifo.genblk1[13].entry.input_buf[5].A ;
 wire \l_fifo.genblk1[13].entry.input_buf[5].X ;
 wire \l_fifo.genblk1[13].entry.input_buf[5].genblk1[0].mid ;
 wire \l_fifo.genblk1[14].entry.empty ;
 wire \l_fifo.genblk1[14].entry.input_buf[0].A ;
 wire \l_fifo.genblk1[14].entry.input_buf[0].X ;
 wire \l_fifo.genblk1[14].entry.input_buf[0].genblk1[0].mid ;
 wire \l_fifo.genblk1[14].entry.input_buf[1].A ;
 wire \l_fifo.genblk1[14].entry.input_buf[1].X ;
 wire \l_fifo.genblk1[14].entry.input_buf[1].genblk1[0].mid ;
 wire \l_fifo.genblk1[14].entry.input_buf[2].A ;
 wire \l_fifo.genblk1[14].entry.input_buf[2].X ;
 wire \l_fifo.genblk1[14].entry.input_buf[2].genblk1[0].mid ;
 wire \l_fifo.genblk1[14].entry.input_buf[3].A ;
 wire \l_fifo.genblk1[14].entry.input_buf[3].X ;
 wire \l_fifo.genblk1[14].entry.input_buf[3].genblk1[0].mid ;
 wire \l_fifo.genblk1[14].entry.input_buf[4].A ;
 wire \l_fifo.genblk1[14].entry.input_buf[4].X ;
 wire \l_fifo.genblk1[14].entry.input_buf[4].genblk1[0].mid ;
 wire \l_fifo.genblk1[14].entry.input_buf[5].A ;
 wire \l_fifo.genblk1[14].entry.input_buf[5].X ;
 wire \l_fifo.genblk1[14].entry.input_buf[5].genblk1[0].mid ;
 wire \l_fifo.genblk1[15].entry.empty ;
 wire \l_fifo.genblk1[15].entry.input_buf[0].A ;
 wire \l_fifo.genblk1[15].entry.input_buf[0].X ;
 wire \l_fifo.genblk1[15].entry.input_buf[0].genblk1[0].mid ;
 wire \l_fifo.genblk1[15].entry.input_buf[1].A ;
 wire \l_fifo.genblk1[15].entry.input_buf[1].X ;
 wire \l_fifo.genblk1[15].entry.input_buf[1].genblk1[0].mid ;
 wire \l_fifo.genblk1[15].entry.input_buf[2].A ;
 wire \l_fifo.genblk1[15].entry.input_buf[2].X ;
 wire \l_fifo.genblk1[15].entry.input_buf[2].genblk1[0].mid ;
 wire \l_fifo.genblk1[15].entry.input_buf[3].A ;
 wire \l_fifo.genblk1[15].entry.input_buf[3].X ;
 wire \l_fifo.genblk1[15].entry.input_buf[3].genblk1[0].mid ;
 wire \l_fifo.genblk1[15].entry.input_buf[4].A ;
 wire \l_fifo.genblk1[15].entry.input_buf[4].X ;
 wire \l_fifo.genblk1[15].entry.input_buf[4].genblk1[0].mid ;
 wire \l_fifo.genblk1[15].entry.input_buf[5].A ;
 wire \l_fifo.genblk1[15].entry.input_buf[5].X ;
 wire \l_fifo.genblk1[15].entry.input_buf[5].genblk1[0].mid ;
 wire \l_fifo.genblk1[16].entry.empty ;
 wire \l_fifo.genblk1[16].entry.input_buf[0].A ;
 wire \l_fifo.genblk1[16].entry.input_buf[0].X ;
 wire \l_fifo.genblk1[16].entry.input_buf[0].genblk1[0].mid ;
 wire \l_fifo.genblk1[16].entry.input_buf[1].A ;
 wire \l_fifo.genblk1[16].entry.input_buf[1].X ;
 wire \l_fifo.genblk1[16].entry.input_buf[1].genblk1[0].mid ;
 wire \l_fifo.genblk1[16].entry.input_buf[2].A ;
 wire \l_fifo.genblk1[16].entry.input_buf[2].X ;
 wire \l_fifo.genblk1[16].entry.input_buf[2].genblk1[0].mid ;
 wire \l_fifo.genblk1[16].entry.input_buf[3].A ;
 wire \l_fifo.genblk1[16].entry.input_buf[3].X ;
 wire \l_fifo.genblk1[16].entry.input_buf[3].genblk1[0].mid ;
 wire \l_fifo.genblk1[16].entry.input_buf[4].A ;
 wire \l_fifo.genblk1[16].entry.input_buf[4].X ;
 wire \l_fifo.genblk1[16].entry.input_buf[4].genblk1[0].mid ;
 wire \l_fifo.genblk1[16].entry.input_buf[5].A ;
 wire \l_fifo.genblk1[16].entry.input_buf[5].X ;
 wire \l_fifo.genblk1[16].entry.input_buf[5].genblk1[0].mid ;
 wire \l_fifo.genblk1[17].entry.empty ;
 wire \l_fifo.genblk1[17].entry.input_buf[0].A ;
 wire \l_fifo.genblk1[17].entry.input_buf[0].X ;
 wire \l_fifo.genblk1[17].entry.input_buf[0].genblk1[0].mid ;
 wire \l_fifo.genblk1[17].entry.input_buf[1].A ;
 wire \l_fifo.genblk1[17].entry.input_buf[1].X ;
 wire \l_fifo.genblk1[17].entry.input_buf[1].genblk1[0].mid ;
 wire \l_fifo.genblk1[17].entry.input_buf[2].A ;
 wire \l_fifo.genblk1[17].entry.input_buf[2].X ;
 wire \l_fifo.genblk1[17].entry.input_buf[2].genblk1[0].mid ;
 wire \l_fifo.genblk1[17].entry.input_buf[3].A ;
 wire \l_fifo.genblk1[17].entry.input_buf[3].X ;
 wire \l_fifo.genblk1[17].entry.input_buf[3].genblk1[0].mid ;
 wire \l_fifo.genblk1[17].entry.input_buf[4].A ;
 wire \l_fifo.genblk1[17].entry.input_buf[4].X ;
 wire \l_fifo.genblk1[17].entry.input_buf[4].genblk1[0].mid ;
 wire \l_fifo.genblk1[17].entry.input_buf[5].A ;
 wire \l_fifo.genblk1[17].entry.input_buf[5].X ;
 wire \l_fifo.genblk1[17].entry.input_buf[5].genblk1[0].mid ;
 wire \l_fifo.genblk1[18].entry.empty ;
 wire \l_fifo.genblk1[18].entry.input_buf[0].A ;
 wire \l_fifo.genblk1[18].entry.input_buf[0].X ;
 wire \l_fifo.genblk1[18].entry.input_buf[0].genblk1[0].mid ;
 wire \l_fifo.genblk1[18].entry.input_buf[1].A ;
 wire \l_fifo.genblk1[18].entry.input_buf[1].X ;
 wire \l_fifo.genblk1[18].entry.input_buf[1].genblk1[0].mid ;
 wire \l_fifo.genblk1[18].entry.input_buf[2].A ;
 wire \l_fifo.genblk1[18].entry.input_buf[2].X ;
 wire \l_fifo.genblk1[18].entry.input_buf[2].genblk1[0].mid ;
 wire \l_fifo.genblk1[18].entry.input_buf[3].A ;
 wire \l_fifo.genblk1[18].entry.input_buf[3].X ;
 wire \l_fifo.genblk1[18].entry.input_buf[3].genblk1[0].mid ;
 wire \l_fifo.genblk1[18].entry.input_buf[4].A ;
 wire \l_fifo.genblk1[18].entry.input_buf[4].X ;
 wire \l_fifo.genblk1[18].entry.input_buf[4].genblk1[0].mid ;
 wire \l_fifo.genblk1[18].entry.input_buf[5].A ;
 wire \l_fifo.genblk1[18].entry.input_buf[5].X ;
 wire \l_fifo.genblk1[18].entry.input_buf[5].genblk1[0].mid ;
 wire \l_fifo.genblk1[19].entry.empty ;
 wire \l_fifo.genblk1[19].entry.input_buf[0].A ;
 wire \l_fifo.genblk1[19].entry.input_buf[0].X ;
 wire \l_fifo.genblk1[19].entry.input_buf[0].genblk1[0].mid ;
 wire \l_fifo.genblk1[19].entry.input_buf[1].A ;
 wire \l_fifo.genblk1[19].entry.input_buf[1].X ;
 wire \l_fifo.genblk1[19].entry.input_buf[1].genblk1[0].mid ;
 wire \l_fifo.genblk1[19].entry.input_buf[2].A ;
 wire \l_fifo.genblk1[19].entry.input_buf[2].X ;
 wire \l_fifo.genblk1[19].entry.input_buf[2].genblk1[0].mid ;
 wire \l_fifo.genblk1[19].entry.input_buf[3].A ;
 wire \l_fifo.genblk1[19].entry.input_buf[3].X ;
 wire \l_fifo.genblk1[19].entry.input_buf[3].genblk1[0].mid ;
 wire \l_fifo.genblk1[19].entry.input_buf[4].A ;
 wire \l_fifo.genblk1[19].entry.input_buf[4].X ;
 wire \l_fifo.genblk1[19].entry.input_buf[4].genblk1[0].mid ;
 wire \l_fifo.genblk1[19].entry.input_buf[5].A ;
 wire \l_fifo.genblk1[19].entry.input_buf[5].X ;
 wire \l_fifo.genblk1[19].entry.input_buf[5].genblk1[0].mid ;
 wire \l_fifo.genblk1[1].entry.empty ;
 wire \l_fifo.genblk1[1].entry.input_buf[0].A ;
 wire \l_fifo.genblk1[1].entry.input_buf[0].X ;
 wire \l_fifo.genblk1[1].entry.input_buf[0].genblk1[0].mid ;
 wire \l_fifo.genblk1[1].entry.input_buf[1].A ;
 wire \l_fifo.genblk1[1].entry.input_buf[1].X ;
 wire \l_fifo.genblk1[1].entry.input_buf[1].genblk1[0].mid ;
 wire \l_fifo.genblk1[1].entry.input_buf[2].A ;
 wire \l_fifo.genblk1[1].entry.input_buf[2].X ;
 wire \l_fifo.genblk1[1].entry.input_buf[2].genblk1[0].mid ;
 wire \l_fifo.genblk1[1].entry.input_buf[3].A ;
 wire \l_fifo.genblk1[1].entry.input_buf[3].X ;
 wire \l_fifo.genblk1[1].entry.input_buf[3].genblk1[0].mid ;
 wire \l_fifo.genblk1[1].entry.input_buf[4].A ;
 wire \l_fifo.genblk1[1].entry.input_buf[4].X ;
 wire \l_fifo.genblk1[1].entry.input_buf[4].genblk1[0].mid ;
 wire \l_fifo.genblk1[1].entry.input_buf[5].A ;
 wire \l_fifo.genblk1[1].entry.input_buf[5].X ;
 wire \l_fifo.genblk1[1].entry.input_buf[5].genblk1[0].mid ;
 wire \l_fifo.genblk1[20].entry.empty ;
 wire \l_fifo.genblk1[20].entry.input_buf[0].A ;
 wire \l_fifo.genblk1[20].entry.input_buf[0].X ;
 wire \l_fifo.genblk1[20].entry.input_buf[0].genblk1[0].mid ;
 wire \l_fifo.genblk1[20].entry.input_buf[1].A ;
 wire \l_fifo.genblk1[20].entry.input_buf[1].X ;
 wire \l_fifo.genblk1[20].entry.input_buf[1].genblk1[0].mid ;
 wire \l_fifo.genblk1[20].entry.input_buf[2].A ;
 wire \l_fifo.genblk1[20].entry.input_buf[2].X ;
 wire \l_fifo.genblk1[20].entry.input_buf[2].genblk1[0].mid ;
 wire \l_fifo.genblk1[20].entry.input_buf[3].A ;
 wire \l_fifo.genblk1[20].entry.input_buf[3].X ;
 wire \l_fifo.genblk1[20].entry.input_buf[3].genblk1[0].mid ;
 wire \l_fifo.genblk1[20].entry.input_buf[4].A ;
 wire \l_fifo.genblk1[20].entry.input_buf[4].X ;
 wire \l_fifo.genblk1[20].entry.input_buf[4].genblk1[0].mid ;
 wire \l_fifo.genblk1[20].entry.input_buf[5].A ;
 wire \l_fifo.genblk1[20].entry.input_buf[5].X ;
 wire \l_fifo.genblk1[20].entry.input_buf[5].genblk1[0].mid ;
 wire \l_fifo.genblk1[21].entry.empty ;
 wire \l_fifo.genblk1[21].entry.input_buf[0].A ;
 wire \l_fifo.genblk1[21].entry.input_buf[0].X ;
 wire \l_fifo.genblk1[21].entry.input_buf[0].genblk1[0].mid ;
 wire \l_fifo.genblk1[21].entry.input_buf[1].A ;
 wire \l_fifo.genblk1[21].entry.input_buf[1].X ;
 wire \l_fifo.genblk1[21].entry.input_buf[1].genblk1[0].mid ;
 wire \l_fifo.genblk1[21].entry.input_buf[2].A ;
 wire \l_fifo.genblk1[21].entry.input_buf[2].X ;
 wire \l_fifo.genblk1[21].entry.input_buf[2].genblk1[0].mid ;
 wire \l_fifo.genblk1[21].entry.input_buf[3].A ;
 wire \l_fifo.genblk1[21].entry.input_buf[3].X ;
 wire \l_fifo.genblk1[21].entry.input_buf[3].genblk1[0].mid ;
 wire \l_fifo.genblk1[21].entry.input_buf[4].A ;
 wire \l_fifo.genblk1[21].entry.input_buf[4].X ;
 wire \l_fifo.genblk1[21].entry.input_buf[4].genblk1[0].mid ;
 wire \l_fifo.genblk1[21].entry.input_buf[5].A ;
 wire \l_fifo.genblk1[21].entry.input_buf[5].X ;
 wire \l_fifo.genblk1[21].entry.input_buf[5].genblk1[0].mid ;
 wire \l_fifo.genblk1[22].entry.empty ;
 wire \l_fifo.genblk1[22].entry.input_buf[0].A ;
 wire \l_fifo.genblk1[22].entry.input_buf[0].X ;
 wire \l_fifo.genblk1[22].entry.input_buf[0].genblk1[0].mid ;
 wire \l_fifo.genblk1[22].entry.input_buf[1].A ;
 wire \l_fifo.genblk1[22].entry.input_buf[1].X ;
 wire \l_fifo.genblk1[22].entry.input_buf[1].genblk1[0].mid ;
 wire \l_fifo.genblk1[22].entry.input_buf[2].A ;
 wire \l_fifo.genblk1[22].entry.input_buf[2].X ;
 wire \l_fifo.genblk1[22].entry.input_buf[2].genblk1[0].mid ;
 wire \l_fifo.genblk1[22].entry.input_buf[3].A ;
 wire \l_fifo.genblk1[22].entry.input_buf[3].X ;
 wire \l_fifo.genblk1[22].entry.input_buf[3].genblk1[0].mid ;
 wire \l_fifo.genblk1[22].entry.input_buf[4].A ;
 wire \l_fifo.genblk1[22].entry.input_buf[4].X ;
 wire \l_fifo.genblk1[22].entry.input_buf[4].genblk1[0].mid ;
 wire \l_fifo.genblk1[22].entry.input_buf[5].A ;
 wire \l_fifo.genblk1[22].entry.input_buf[5].X ;
 wire \l_fifo.genblk1[22].entry.input_buf[5].genblk1[0].mid ;
 wire \l_fifo.genblk1[23].entry.empty ;
 wire \l_fifo.genblk1[23].entry.input_buf[0].A ;
 wire \l_fifo.genblk1[23].entry.input_buf[0].X ;
 wire \l_fifo.genblk1[23].entry.input_buf[0].genblk1[0].mid ;
 wire \l_fifo.genblk1[23].entry.input_buf[1].A ;
 wire \l_fifo.genblk1[23].entry.input_buf[1].X ;
 wire \l_fifo.genblk1[23].entry.input_buf[1].genblk1[0].mid ;
 wire \l_fifo.genblk1[23].entry.input_buf[2].A ;
 wire \l_fifo.genblk1[23].entry.input_buf[2].X ;
 wire \l_fifo.genblk1[23].entry.input_buf[2].genblk1[0].mid ;
 wire \l_fifo.genblk1[23].entry.input_buf[3].A ;
 wire \l_fifo.genblk1[23].entry.input_buf[3].X ;
 wire \l_fifo.genblk1[23].entry.input_buf[3].genblk1[0].mid ;
 wire \l_fifo.genblk1[23].entry.input_buf[4].A ;
 wire \l_fifo.genblk1[23].entry.input_buf[4].X ;
 wire \l_fifo.genblk1[23].entry.input_buf[4].genblk1[0].mid ;
 wire \l_fifo.genblk1[23].entry.input_buf[5].A ;
 wire \l_fifo.genblk1[23].entry.input_buf[5].X ;
 wire \l_fifo.genblk1[23].entry.input_buf[5].genblk1[0].mid ;
 wire \l_fifo.genblk1[24].entry.empty ;
 wire \l_fifo.genblk1[24].entry.input_buf[0].A ;
 wire \l_fifo.genblk1[24].entry.input_buf[0].X ;
 wire \l_fifo.genblk1[24].entry.input_buf[0].genblk1[0].mid ;
 wire \l_fifo.genblk1[24].entry.input_buf[1].A ;
 wire \l_fifo.genblk1[24].entry.input_buf[1].X ;
 wire \l_fifo.genblk1[24].entry.input_buf[1].genblk1[0].mid ;
 wire \l_fifo.genblk1[24].entry.input_buf[2].A ;
 wire \l_fifo.genblk1[24].entry.input_buf[2].X ;
 wire \l_fifo.genblk1[24].entry.input_buf[2].genblk1[0].mid ;
 wire \l_fifo.genblk1[24].entry.input_buf[3].A ;
 wire \l_fifo.genblk1[24].entry.input_buf[3].X ;
 wire \l_fifo.genblk1[24].entry.input_buf[3].genblk1[0].mid ;
 wire \l_fifo.genblk1[24].entry.input_buf[4].A ;
 wire \l_fifo.genblk1[24].entry.input_buf[4].X ;
 wire \l_fifo.genblk1[24].entry.input_buf[4].genblk1[0].mid ;
 wire \l_fifo.genblk1[24].entry.input_buf[5].A ;
 wire \l_fifo.genblk1[24].entry.input_buf[5].X ;
 wire \l_fifo.genblk1[24].entry.input_buf[5].genblk1[0].mid ;
 wire \l_fifo.genblk1[25].entry.empty ;
 wire \l_fifo.genblk1[25].entry.input_buf[0].A ;
 wire \l_fifo.genblk1[25].entry.input_buf[0].X ;
 wire \l_fifo.genblk1[25].entry.input_buf[0].genblk1[0].mid ;
 wire \l_fifo.genblk1[25].entry.input_buf[1].A ;
 wire \l_fifo.genblk1[25].entry.input_buf[1].X ;
 wire \l_fifo.genblk1[25].entry.input_buf[1].genblk1[0].mid ;
 wire \l_fifo.genblk1[25].entry.input_buf[2].A ;
 wire \l_fifo.genblk1[25].entry.input_buf[2].X ;
 wire \l_fifo.genblk1[25].entry.input_buf[2].genblk1[0].mid ;
 wire \l_fifo.genblk1[25].entry.input_buf[3].A ;
 wire \l_fifo.genblk1[25].entry.input_buf[3].X ;
 wire \l_fifo.genblk1[25].entry.input_buf[3].genblk1[0].mid ;
 wire \l_fifo.genblk1[25].entry.input_buf[4].A ;
 wire \l_fifo.genblk1[25].entry.input_buf[4].X ;
 wire \l_fifo.genblk1[25].entry.input_buf[4].genblk1[0].mid ;
 wire \l_fifo.genblk1[25].entry.input_buf[5].A ;
 wire \l_fifo.genblk1[25].entry.input_buf[5].X ;
 wire \l_fifo.genblk1[25].entry.input_buf[5].genblk1[0].mid ;
 wire \l_fifo.genblk1[26].entry.empty ;
 wire \l_fifo.genblk1[26].entry.input_buf[0].A ;
 wire \l_fifo.genblk1[26].entry.input_buf[0].X ;
 wire \l_fifo.genblk1[26].entry.input_buf[0].genblk1[0].mid ;
 wire \l_fifo.genblk1[26].entry.input_buf[1].A ;
 wire \l_fifo.genblk1[26].entry.input_buf[1].X ;
 wire \l_fifo.genblk1[26].entry.input_buf[1].genblk1[0].mid ;
 wire \l_fifo.genblk1[26].entry.input_buf[2].A ;
 wire \l_fifo.genblk1[26].entry.input_buf[2].X ;
 wire \l_fifo.genblk1[26].entry.input_buf[2].genblk1[0].mid ;
 wire \l_fifo.genblk1[26].entry.input_buf[3].A ;
 wire \l_fifo.genblk1[26].entry.input_buf[3].X ;
 wire \l_fifo.genblk1[26].entry.input_buf[3].genblk1[0].mid ;
 wire \l_fifo.genblk1[26].entry.input_buf[4].A ;
 wire \l_fifo.genblk1[26].entry.input_buf[4].X ;
 wire \l_fifo.genblk1[26].entry.input_buf[4].genblk1[0].mid ;
 wire \l_fifo.genblk1[26].entry.input_buf[5].A ;
 wire \l_fifo.genblk1[26].entry.input_buf[5].X ;
 wire \l_fifo.genblk1[26].entry.input_buf[5].genblk1[0].mid ;
 wire \l_fifo.genblk1[27].entry.empty ;
 wire \l_fifo.genblk1[27].entry.input_buf[0].A ;
 wire \l_fifo.genblk1[27].entry.input_buf[0].X ;
 wire \l_fifo.genblk1[27].entry.input_buf[0].genblk1[0].mid ;
 wire \l_fifo.genblk1[27].entry.input_buf[1].A ;
 wire \l_fifo.genblk1[27].entry.input_buf[1].X ;
 wire \l_fifo.genblk1[27].entry.input_buf[1].genblk1[0].mid ;
 wire \l_fifo.genblk1[27].entry.input_buf[2].A ;
 wire \l_fifo.genblk1[27].entry.input_buf[2].X ;
 wire \l_fifo.genblk1[27].entry.input_buf[2].genblk1[0].mid ;
 wire \l_fifo.genblk1[27].entry.input_buf[3].A ;
 wire \l_fifo.genblk1[27].entry.input_buf[3].X ;
 wire \l_fifo.genblk1[27].entry.input_buf[3].genblk1[0].mid ;
 wire \l_fifo.genblk1[27].entry.input_buf[4].A ;
 wire \l_fifo.genblk1[27].entry.input_buf[4].X ;
 wire \l_fifo.genblk1[27].entry.input_buf[4].genblk1[0].mid ;
 wire \l_fifo.genblk1[27].entry.input_buf[5].A ;
 wire \l_fifo.genblk1[27].entry.input_buf[5].X ;
 wire \l_fifo.genblk1[27].entry.input_buf[5].genblk1[0].mid ;
 wire \l_fifo.genblk1[28].entry.empty ;
 wire \l_fifo.genblk1[28].entry.input_buf[0].A ;
 wire \l_fifo.genblk1[28].entry.input_buf[0].X ;
 wire \l_fifo.genblk1[28].entry.input_buf[0].genblk1[0].mid ;
 wire \l_fifo.genblk1[28].entry.input_buf[1].A ;
 wire \l_fifo.genblk1[28].entry.input_buf[1].X ;
 wire \l_fifo.genblk1[28].entry.input_buf[1].genblk1[0].mid ;
 wire \l_fifo.genblk1[28].entry.input_buf[2].A ;
 wire \l_fifo.genblk1[28].entry.input_buf[2].X ;
 wire \l_fifo.genblk1[28].entry.input_buf[2].genblk1[0].mid ;
 wire \l_fifo.genblk1[28].entry.input_buf[3].A ;
 wire \l_fifo.genblk1[28].entry.input_buf[3].X ;
 wire \l_fifo.genblk1[28].entry.input_buf[3].genblk1[0].mid ;
 wire \l_fifo.genblk1[28].entry.input_buf[4].A ;
 wire \l_fifo.genblk1[28].entry.input_buf[4].X ;
 wire \l_fifo.genblk1[28].entry.input_buf[4].genblk1[0].mid ;
 wire \l_fifo.genblk1[28].entry.input_buf[5].A ;
 wire \l_fifo.genblk1[28].entry.input_buf[5].X ;
 wire \l_fifo.genblk1[28].entry.input_buf[5].genblk1[0].mid ;
 wire \l_fifo.genblk1[29].entry.empty ;
 wire \l_fifo.genblk1[29].entry.input_buf[0].A ;
 wire \l_fifo.genblk1[29].entry.input_buf[0].X ;
 wire \l_fifo.genblk1[29].entry.input_buf[0].genblk1[0].mid ;
 wire \l_fifo.genblk1[29].entry.input_buf[1].A ;
 wire \l_fifo.genblk1[29].entry.input_buf[1].X ;
 wire \l_fifo.genblk1[29].entry.input_buf[1].genblk1[0].mid ;
 wire \l_fifo.genblk1[29].entry.input_buf[2].A ;
 wire \l_fifo.genblk1[29].entry.input_buf[2].X ;
 wire \l_fifo.genblk1[29].entry.input_buf[2].genblk1[0].mid ;
 wire \l_fifo.genblk1[29].entry.input_buf[3].A ;
 wire \l_fifo.genblk1[29].entry.input_buf[3].X ;
 wire \l_fifo.genblk1[29].entry.input_buf[3].genblk1[0].mid ;
 wire \l_fifo.genblk1[29].entry.input_buf[4].A ;
 wire \l_fifo.genblk1[29].entry.input_buf[4].X ;
 wire \l_fifo.genblk1[29].entry.input_buf[4].genblk1[0].mid ;
 wire \l_fifo.genblk1[29].entry.input_buf[5].A ;
 wire \l_fifo.genblk1[29].entry.input_buf[5].X ;
 wire \l_fifo.genblk1[29].entry.input_buf[5].genblk1[0].mid ;
 wire \l_fifo.genblk1[2].entry.empty ;
 wire \l_fifo.genblk1[2].entry.input_buf[0].A ;
 wire \l_fifo.genblk1[2].entry.input_buf[0].X ;
 wire \l_fifo.genblk1[2].entry.input_buf[0].genblk1[0].mid ;
 wire \l_fifo.genblk1[2].entry.input_buf[1].A ;
 wire \l_fifo.genblk1[2].entry.input_buf[1].X ;
 wire \l_fifo.genblk1[2].entry.input_buf[1].genblk1[0].mid ;
 wire \l_fifo.genblk1[2].entry.input_buf[2].A ;
 wire \l_fifo.genblk1[2].entry.input_buf[2].X ;
 wire \l_fifo.genblk1[2].entry.input_buf[2].genblk1[0].mid ;
 wire \l_fifo.genblk1[2].entry.input_buf[3].A ;
 wire \l_fifo.genblk1[2].entry.input_buf[3].X ;
 wire \l_fifo.genblk1[2].entry.input_buf[3].genblk1[0].mid ;
 wire \l_fifo.genblk1[2].entry.input_buf[4].A ;
 wire \l_fifo.genblk1[2].entry.input_buf[4].X ;
 wire \l_fifo.genblk1[2].entry.input_buf[4].genblk1[0].mid ;
 wire \l_fifo.genblk1[2].entry.input_buf[5].A ;
 wire \l_fifo.genblk1[2].entry.input_buf[5].X ;
 wire \l_fifo.genblk1[2].entry.input_buf[5].genblk1[0].mid ;
 wire \l_fifo.genblk1[30].entry.empty ;
 wire \l_fifo.genblk1[30].entry.input_buf[0].A ;
 wire \l_fifo.genblk1[30].entry.input_buf[0].X ;
 wire \l_fifo.genblk1[30].entry.input_buf[0].genblk1[0].mid ;
 wire \l_fifo.genblk1[30].entry.input_buf[1].A ;
 wire \l_fifo.genblk1[30].entry.input_buf[1].X ;
 wire \l_fifo.genblk1[30].entry.input_buf[1].genblk1[0].mid ;
 wire \l_fifo.genblk1[30].entry.input_buf[2].A ;
 wire \l_fifo.genblk1[30].entry.input_buf[2].X ;
 wire \l_fifo.genblk1[30].entry.input_buf[2].genblk1[0].mid ;
 wire \l_fifo.genblk1[30].entry.input_buf[3].A ;
 wire \l_fifo.genblk1[30].entry.input_buf[3].X ;
 wire \l_fifo.genblk1[30].entry.input_buf[3].genblk1[0].mid ;
 wire \l_fifo.genblk1[30].entry.input_buf[4].A ;
 wire \l_fifo.genblk1[30].entry.input_buf[4].X ;
 wire \l_fifo.genblk1[30].entry.input_buf[4].genblk1[0].mid ;
 wire \l_fifo.genblk1[30].entry.input_buf[5].A ;
 wire \l_fifo.genblk1[30].entry.input_buf[5].X ;
 wire \l_fifo.genblk1[30].entry.input_buf[5].genblk1[0].mid ;
 wire \l_fifo.genblk1[31].entry.empty ;
 wire \l_fifo.genblk1[31].entry.input_buf[0].A ;
 wire \l_fifo.genblk1[31].entry.input_buf[0].X ;
 wire \l_fifo.genblk1[31].entry.input_buf[0].genblk1[0].mid ;
 wire \l_fifo.genblk1[31].entry.input_buf[1].A ;
 wire \l_fifo.genblk1[31].entry.input_buf[1].X ;
 wire \l_fifo.genblk1[31].entry.input_buf[1].genblk1[0].mid ;
 wire \l_fifo.genblk1[31].entry.input_buf[2].A ;
 wire \l_fifo.genblk1[31].entry.input_buf[2].X ;
 wire \l_fifo.genblk1[31].entry.input_buf[2].genblk1[0].mid ;
 wire \l_fifo.genblk1[31].entry.input_buf[3].A ;
 wire \l_fifo.genblk1[31].entry.input_buf[3].X ;
 wire \l_fifo.genblk1[31].entry.input_buf[3].genblk1[0].mid ;
 wire \l_fifo.genblk1[31].entry.input_buf[4].A ;
 wire \l_fifo.genblk1[31].entry.input_buf[4].X ;
 wire \l_fifo.genblk1[31].entry.input_buf[4].genblk1[0].mid ;
 wire \l_fifo.genblk1[31].entry.input_buf[5].A ;
 wire \l_fifo.genblk1[31].entry.input_buf[5].X ;
 wire \l_fifo.genblk1[31].entry.input_buf[5].genblk1[0].mid ;
 wire \l_fifo.genblk1[32].entry.empty ;
 wire \l_fifo.genblk1[32].entry.input_buf[0].A ;
 wire \l_fifo.genblk1[32].entry.input_buf[0].X ;
 wire \l_fifo.genblk1[32].entry.input_buf[0].genblk1[0].mid ;
 wire \l_fifo.genblk1[32].entry.input_buf[1].A ;
 wire \l_fifo.genblk1[32].entry.input_buf[1].X ;
 wire \l_fifo.genblk1[32].entry.input_buf[1].genblk1[0].mid ;
 wire \l_fifo.genblk1[32].entry.input_buf[2].A ;
 wire \l_fifo.genblk1[32].entry.input_buf[2].X ;
 wire \l_fifo.genblk1[32].entry.input_buf[2].genblk1[0].mid ;
 wire \l_fifo.genblk1[32].entry.input_buf[3].A ;
 wire \l_fifo.genblk1[32].entry.input_buf[3].X ;
 wire \l_fifo.genblk1[32].entry.input_buf[3].genblk1[0].mid ;
 wire \l_fifo.genblk1[32].entry.input_buf[4].A ;
 wire \l_fifo.genblk1[32].entry.input_buf[4].X ;
 wire \l_fifo.genblk1[32].entry.input_buf[4].genblk1[0].mid ;
 wire \l_fifo.genblk1[32].entry.input_buf[5].A ;
 wire \l_fifo.genblk1[32].entry.input_buf[5].X ;
 wire \l_fifo.genblk1[32].entry.input_buf[5].genblk1[0].mid ;
 wire \l_fifo.genblk1[33].entry.empty ;
 wire \l_fifo.genblk1[33].entry.input_buf[0].A ;
 wire \l_fifo.genblk1[33].entry.input_buf[0].X ;
 wire \l_fifo.genblk1[33].entry.input_buf[0].genblk1[0].mid ;
 wire \l_fifo.genblk1[33].entry.input_buf[1].A ;
 wire \l_fifo.genblk1[33].entry.input_buf[1].X ;
 wire \l_fifo.genblk1[33].entry.input_buf[1].genblk1[0].mid ;
 wire \l_fifo.genblk1[33].entry.input_buf[2].A ;
 wire \l_fifo.genblk1[33].entry.input_buf[2].X ;
 wire \l_fifo.genblk1[33].entry.input_buf[2].genblk1[0].mid ;
 wire \l_fifo.genblk1[33].entry.input_buf[3].A ;
 wire \l_fifo.genblk1[33].entry.input_buf[3].X ;
 wire \l_fifo.genblk1[33].entry.input_buf[3].genblk1[0].mid ;
 wire \l_fifo.genblk1[33].entry.input_buf[4].A ;
 wire \l_fifo.genblk1[33].entry.input_buf[4].X ;
 wire \l_fifo.genblk1[33].entry.input_buf[4].genblk1[0].mid ;
 wire \l_fifo.genblk1[33].entry.input_buf[5].A ;
 wire \l_fifo.genblk1[33].entry.input_buf[5].X ;
 wire \l_fifo.genblk1[33].entry.input_buf[5].genblk1[0].mid ;
 wire \l_fifo.genblk1[34].entry.empty ;
 wire \l_fifo.genblk1[34].entry.input_buf[0].A ;
 wire \l_fifo.genblk1[34].entry.input_buf[0].X ;
 wire \l_fifo.genblk1[34].entry.input_buf[0].genblk1[0].mid ;
 wire \l_fifo.genblk1[34].entry.input_buf[1].A ;
 wire \l_fifo.genblk1[34].entry.input_buf[1].X ;
 wire \l_fifo.genblk1[34].entry.input_buf[1].genblk1[0].mid ;
 wire \l_fifo.genblk1[34].entry.input_buf[2].A ;
 wire \l_fifo.genblk1[34].entry.input_buf[2].X ;
 wire \l_fifo.genblk1[34].entry.input_buf[2].genblk1[0].mid ;
 wire \l_fifo.genblk1[34].entry.input_buf[3].A ;
 wire \l_fifo.genblk1[34].entry.input_buf[3].X ;
 wire \l_fifo.genblk1[34].entry.input_buf[3].genblk1[0].mid ;
 wire \l_fifo.genblk1[34].entry.input_buf[4].A ;
 wire \l_fifo.genblk1[34].entry.input_buf[4].X ;
 wire \l_fifo.genblk1[34].entry.input_buf[4].genblk1[0].mid ;
 wire \l_fifo.genblk1[34].entry.input_buf[5].A ;
 wire \l_fifo.genblk1[34].entry.input_buf[5].X ;
 wire \l_fifo.genblk1[34].entry.input_buf[5].genblk1[0].mid ;
 wire \l_fifo.genblk1[35].entry.empty ;
 wire \l_fifo.genblk1[35].entry.input_buf[0].A ;
 wire \l_fifo.genblk1[35].entry.input_buf[0].X ;
 wire \l_fifo.genblk1[35].entry.input_buf[0].genblk1[0].mid ;
 wire \l_fifo.genblk1[35].entry.input_buf[1].A ;
 wire \l_fifo.genblk1[35].entry.input_buf[1].X ;
 wire \l_fifo.genblk1[35].entry.input_buf[1].genblk1[0].mid ;
 wire \l_fifo.genblk1[35].entry.input_buf[2].A ;
 wire \l_fifo.genblk1[35].entry.input_buf[2].X ;
 wire \l_fifo.genblk1[35].entry.input_buf[2].genblk1[0].mid ;
 wire \l_fifo.genblk1[35].entry.input_buf[3].A ;
 wire \l_fifo.genblk1[35].entry.input_buf[3].X ;
 wire \l_fifo.genblk1[35].entry.input_buf[3].genblk1[0].mid ;
 wire \l_fifo.genblk1[35].entry.input_buf[4].A ;
 wire \l_fifo.genblk1[35].entry.input_buf[4].X ;
 wire \l_fifo.genblk1[35].entry.input_buf[4].genblk1[0].mid ;
 wire \l_fifo.genblk1[35].entry.input_buf[5].A ;
 wire \l_fifo.genblk1[35].entry.input_buf[5].X ;
 wire \l_fifo.genblk1[35].entry.input_buf[5].genblk1[0].mid ;
 wire \l_fifo.genblk1[36].entry.empty ;
 wire \l_fifo.genblk1[36].entry.input_buf[0].A ;
 wire \l_fifo.genblk1[36].entry.input_buf[0].X ;
 wire \l_fifo.genblk1[36].entry.input_buf[0].genblk1[0].mid ;
 wire \l_fifo.genblk1[36].entry.input_buf[1].A ;
 wire \l_fifo.genblk1[36].entry.input_buf[1].X ;
 wire \l_fifo.genblk1[36].entry.input_buf[1].genblk1[0].mid ;
 wire \l_fifo.genblk1[36].entry.input_buf[2].A ;
 wire \l_fifo.genblk1[36].entry.input_buf[2].X ;
 wire \l_fifo.genblk1[36].entry.input_buf[2].genblk1[0].mid ;
 wire \l_fifo.genblk1[36].entry.input_buf[3].A ;
 wire \l_fifo.genblk1[36].entry.input_buf[3].X ;
 wire \l_fifo.genblk1[36].entry.input_buf[3].genblk1[0].mid ;
 wire \l_fifo.genblk1[36].entry.input_buf[4].A ;
 wire \l_fifo.genblk1[36].entry.input_buf[4].X ;
 wire \l_fifo.genblk1[36].entry.input_buf[4].genblk1[0].mid ;
 wire \l_fifo.genblk1[36].entry.input_buf[5].A ;
 wire \l_fifo.genblk1[36].entry.input_buf[5].X ;
 wire \l_fifo.genblk1[36].entry.input_buf[5].genblk1[0].mid ;
 wire \l_fifo.genblk1[37].entry.empty ;
 wire \l_fifo.genblk1[37].entry.input_buf[0].A ;
 wire \l_fifo.genblk1[37].entry.input_buf[0].X ;
 wire \l_fifo.genblk1[37].entry.input_buf[0].genblk1[0].mid ;
 wire \l_fifo.genblk1[37].entry.input_buf[1].A ;
 wire \l_fifo.genblk1[37].entry.input_buf[1].X ;
 wire \l_fifo.genblk1[37].entry.input_buf[1].genblk1[0].mid ;
 wire \l_fifo.genblk1[37].entry.input_buf[2].A ;
 wire \l_fifo.genblk1[37].entry.input_buf[2].X ;
 wire \l_fifo.genblk1[37].entry.input_buf[2].genblk1[0].mid ;
 wire \l_fifo.genblk1[37].entry.input_buf[3].A ;
 wire \l_fifo.genblk1[37].entry.input_buf[3].X ;
 wire \l_fifo.genblk1[37].entry.input_buf[3].genblk1[0].mid ;
 wire \l_fifo.genblk1[37].entry.input_buf[4].A ;
 wire \l_fifo.genblk1[37].entry.input_buf[4].X ;
 wire \l_fifo.genblk1[37].entry.input_buf[4].genblk1[0].mid ;
 wire \l_fifo.genblk1[37].entry.input_buf[5].A ;
 wire \l_fifo.genblk1[37].entry.input_buf[5].X ;
 wire \l_fifo.genblk1[37].entry.input_buf[5].genblk1[0].mid ;
 wire \l_fifo.genblk1[38].entry.empty ;
 wire \l_fifo.genblk1[38].entry.input_buf[0].A ;
 wire \l_fifo.genblk1[38].entry.input_buf[0].X ;
 wire \l_fifo.genblk1[38].entry.input_buf[0].genblk1[0].mid ;
 wire \l_fifo.genblk1[38].entry.input_buf[1].A ;
 wire \l_fifo.genblk1[38].entry.input_buf[1].X ;
 wire \l_fifo.genblk1[38].entry.input_buf[1].genblk1[0].mid ;
 wire \l_fifo.genblk1[38].entry.input_buf[2].A ;
 wire \l_fifo.genblk1[38].entry.input_buf[2].X ;
 wire \l_fifo.genblk1[38].entry.input_buf[2].genblk1[0].mid ;
 wire \l_fifo.genblk1[38].entry.input_buf[3].A ;
 wire \l_fifo.genblk1[38].entry.input_buf[3].X ;
 wire \l_fifo.genblk1[38].entry.input_buf[3].genblk1[0].mid ;
 wire \l_fifo.genblk1[38].entry.input_buf[4].A ;
 wire \l_fifo.genblk1[38].entry.input_buf[4].X ;
 wire \l_fifo.genblk1[38].entry.input_buf[4].genblk1[0].mid ;
 wire \l_fifo.genblk1[38].entry.input_buf[5].A ;
 wire \l_fifo.genblk1[38].entry.input_buf[5].X ;
 wire \l_fifo.genblk1[38].entry.input_buf[5].genblk1[0].mid ;
 wire \l_fifo.genblk1[39].entry.empty ;
 wire \l_fifo.genblk1[39].entry.input_buf[0].A ;
 wire \l_fifo.genblk1[39].entry.input_buf[0].X ;
 wire \l_fifo.genblk1[39].entry.input_buf[0].genblk1[0].mid ;
 wire \l_fifo.genblk1[39].entry.input_buf[1].A ;
 wire \l_fifo.genblk1[39].entry.input_buf[1].X ;
 wire \l_fifo.genblk1[39].entry.input_buf[1].genblk1[0].mid ;
 wire \l_fifo.genblk1[39].entry.input_buf[2].A ;
 wire \l_fifo.genblk1[39].entry.input_buf[2].X ;
 wire \l_fifo.genblk1[39].entry.input_buf[2].genblk1[0].mid ;
 wire \l_fifo.genblk1[39].entry.input_buf[3].A ;
 wire \l_fifo.genblk1[39].entry.input_buf[3].X ;
 wire \l_fifo.genblk1[39].entry.input_buf[3].genblk1[0].mid ;
 wire \l_fifo.genblk1[39].entry.input_buf[4].A ;
 wire \l_fifo.genblk1[39].entry.input_buf[4].X ;
 wire \l_fifo.genblk1[39].entry.input_buf[4].genblk1[0].mid ;
 wire \l_fifo.genblk1[39].entry.input_buf[5].A ;
 wire \l_fifo.genblk1[39].entry.input_buf[5].X ;
 wire \l_fifo.genblk1[39].entry.input_buf[5].genblk1[0].mid ;
 wire \l_fifo.genblk1[3].entry.empty ;
 wire \l_fifo.genblk1[3].entry.input_buf[0].A ;
 wire \l_fifo.genblk1[3].entry.input_buf[0].X ;
 wire \l_fifo.genblk1[3].entry.input_buf[0].genblk1[0].mid ;
 wire \l_fifo.genblk1[3].entry.input_buf[1].A ;
 wire \l_fifo.genblk1[3].entry.input_buf[1].X ;
 wire \l_fifo.genblk1[3].entry.input_buf[1].genblk1[0].mid ;
 wire \l_fifo.genblk1[3].entry.input_buf[2].A ;
 wire \l_fifo.genblk1[3].entry.input_buf[2].X ;
 wire \l_fifo.genblk1[3].entry.input_buf[2].genblk1[0].mid ;
 wire \l_fifo.genblk1[3].entry.input_buf[3].A ;
 wire \l_fifo.genblk1[3].entry.input_buf[3].X ;
 wire \l_fifo.genblk1[3].entry.input_buf[3].genblk1[0].mid ;
 wire \l_fifo.genblk1[3].entry.input_buf[4].A ;
 wire \l_fifo.genblk1[3].entry.input_buf[4].X ;
 wire \l_fifo.genblk1[3].entry.input_buf[4].genblk1[0].mid ;
 wire \l_fifo.genblk1[3].entry.input_buf[5].A ;
 wire \l_fifo.genblk1[3].entry.input_buf[5].X ;
 wire \l_fifo.genblk1[3].entry.input_buf[5].genblk1[0].mid ;
 wire \l_fifo.genblk1[40].entry.empty ;
 wire \l_fifo.genblk1[40].entry.input_buf[0].A ;
 wire \l_fifo.genblk1[40].entry.input_buf[0].X ;
 wire \l_fifo.genblk1[40].entry.input_buf[0].genblk1[0].mid ;
 wire \l_fifo.genblk1[40].entry.input_buf[1].A ;
 wire \l_fifo.genblk1[40].entry.input_buf[1].X ;
 wire \l_fifo.genblk1[40].entry.input_buf[1].genblk1[0].mid ;
 wire \l_fifo.genblk1[40].entry.input_buf[2].A ;
 wire \l_fifo.genblk1[40].entry.input_buf[2].X ;
 wire \l_fifo.genblk1[40].entry.input_buf[2].genblk1[0].mid ;
 wire \l_fifo.genblk1[40].entry.input_buf[3].A ;
 wire \l_fifo.genblk1[40].entry.input_buf[3].X ;
 wire \l_fifo.genblk1[40].entry.input_buf[3].genblk1[0].mid ;
 wire \l_fifo.genblk1[40].entry.input_buf[4].A ;
 wire \l_fifo.genblk1[40].entry.input_buf[4].X ;
 wire \l_fifo.genblk1[40].entry.input_buf[4].genblk1[0].mid ;
 wire \l_fifo.genblk1[40].entry.input_buf[5].A ;
 wire \l_fifo.genblk1[40].entry.input_buf[5].X ;
 wire \l_fifo.genblk1[40].entry.input_buf[5].genblk1[0].mid ;
 wire \l_fifo.genblk1[41].entry.empty ;
 wire \l_fifo.genblk1[41].entry.input_buf[0].A ;
 wire \l_fifo.genblk1[41].entry.input_buf[0].X ;
 wire \l_fifo.genblk1[41].entry.input_buf[0].genblk1[0].mid ;
 wire \l_fifo.genblk1[41].entry.input_buf[1].A ;
 wire \l_fifo.genblk1[41].entry.input_buf[1].X ;
 wire \l_fifo.genblk1[41].entry.input_buf[1].genblk1[0].mid ;
 wire \l_fifo.genblk1[41].entry.input_buf[2].A ;
 wire \l_fifo.genblk1[41].entry.input_buf[2].X ;
 wire \l_fifo.genblk1[41].entry.input_buf[2].genblk1[0].mid ;
 wire \l_fifo.genblk1[41].entry.input_buf[3].A ;
 wire \l_fifo.genblk1[41].entry.input_buf[3].X ;
 wire \l_fifo.genblk1[41].entry.input_buf[3].genblk1[0].mid ;
 wire \l_fifo.genblk1[41].entry.input_buf[4].A ;
 wire \l_fifo.genblk1[41].entry.input_buf[4].X ;
 wire \l_fifo.genblk1[41].entry.input_buf[4].genblk1[0].mid ;
 wire \l_fifo.genblk1[41].entry.input_buf[5].A ;
 wire \l_fifo.genblk1[41].entry.input_buf[5].X ;
 wire \l_fifo.genblk1[41].entry.input_buf[5].genblk1[0].mid ;
 wire \l_fifo.genblk1[42].entry.empty ;
 wire \l_fifo.genblk1[42].entry.input_buf[0].A ;
 wire \l_fifo.genblk1[42].entry.input_buf[0].X ;
 wire \l_fifo.genblk1[42].entry.input_buf[0].genblk1[0].mid ;
 wire \l_fifo.genblk1[42].entry.input_buf[1].A ;
 wire \l_fifo.genblk1[42].entry.input_buf[1].X ;
 wire \l_fifo.genblk1[42].entry.input_buf[1].genblk1[0].mid ;
 wire \l_fifo.genblk1[42].entry.input_buf[2].A ;
 wire \l_fifo.genblk1[42].entry.input_buf[2].X ;
 wire \l_fifo.genblk1[42].entry.input_buf[2].genblk1[0].mid ;
 wire \l_fifo.genblk1[42].entry.input_buf[3].A ;
 wire \l_fifo.genblk1[42].entry.input_buf[3].X ;
 wire \l_fifo.genblk1[42].entry.input_buf[3].genblk1[0].mid ;
 wire \l_fifo.genblk1[42].entry.input_buf[4].A ;
 wire \l_fifo.genblk1[42].entry.input_buf[4].X ;
 wire \l_fifo.genblk1[42].entry.input_buf[4].genblk1[0].mid ;
 wire \l_fifo.genblk1[42].entry.input_buf[5].A ;
 wire \l_fifo.genblk1[42].entry.input_buf[5].X ;
 wire \l_fifo.genblk1[42].entry.input_buf[5].genblk1[0].mid ;
 wire \l_fifo.genblk1[43].entry.empty ;
 wire \l_fifo.genblk1[43].entry.input_buf[0].A ;
 wire \l_fifo.genblk1[43].entry.input_buf[0].X ;
 wire \l_fifo.genblk1[43].entry.input_buf[0].genblk1[0].mid ;
 wire \l_fifo.genblk1[43].entry.input_buf[1].A ;
 wire \l_fifo.genblk1[43].entry.input_buf[1].X ;
 wire \l_fifo.genblk1[43].entry.input_buf[1].genblk1[0].mid ;
 wire \l_fifo.genblk1[43].entry.input_buf[2].A ;
 wire \l_fifo.genblk1[43].entry.input_buf[2].X ;
 wire \l_fifo.genblk1[43].entry.input_buf[2].genblk1[0].mid ;
 wire \l_fifo.genblk1[43].entry.input_buf[3].A ;
 wire \l_fifo.genblk1[43].entry.input_buf[3].X ;
 wire \l_fifo.genblk1[43].entry.input_buf[3].genblk1[0].mid ;
 wire \l_fifo.genblk1[43].entry.input_buf[4].A ;
 wire \l_fifo.genblk1[43].entry.input_buf[4].X ;
 wire \l_fifo.genblk1[43].entry.input_buf[4].genblk1[0].mid ;
 wire \l_fifo.genblk1[43].entry.input_buf[5].A ;
 wire \l_fifo.genblk1[43].entry.input_buf[5].X ;
 wire \l_fifo.genblk1[43].entry.input_buf[5].genblk1[0].mid ;
 wire \l_fifo.genblk1[44].entry.empty ;
 wire \l_fifo.genblk1[44].entry.input_buf[0].A ;
 wire \l_fifo.genblk1[44].entry.input_buf[0].X ;
 wire \l_fifo.genblk1[44].entry.input_buf[0].genblk1[0].mid ;
 wire \l_fifo.genblk1[44].entry.input_buf[1].A ;
 wire \l_fifo.genblk1[44].entry.input_buf[1].X ;
 wire \l_fifo.genblk1[44].entry.input_buf[1].genblk1[0].mid ;
 wire \l_fifo.genblk1[44].entry.input_buf[2].A ;
 wire \l_fifo.genblk1[44].entry.input_buf[2].X ;
 wire \l_fifo.genblk1[44].entry.input_buf[2].genblk1[0].mid ;
 wire \l_fifo.genblk1[44].entry.input_buf[3].A ;
 wire \l_fifo.genblk1[44].entry.input_buf[3].X ;
 wire \l_fifo.genblk1[44].entry.input_buf[3].genblk1[0].mid ;
 wire \l_fifo.genblk1[44].entry.input_buf[4].A ;
 wire \l_fifo.genblk1[44].entry.input_buf[4].X ;
 wire \l_fifo.genblk1[44].entry.input_buf[4].genblk1[0].mid ;
 wire \l_fifo.genblk1[44].entry.input_buf[5].A ;
 wire \l_fifo.genblk1[44].entry.input_buf[5].X ;
 wire \l_fifo.genblk1[44].entry.input_buf[5].genblk1[0].mid ;
 wire \l_fifo.genblk1[45].entry.empty ;
 wire \l_fifo.genblk1[45].entry.input_buf[0].A ;
 wire \l_fifo.genblk1[45].entry.input_buf[0].X ;
 wire \l_fifo.genblk1[45].entry.input_buf[0].genblk1[0].mid ;
 wire \l_fifo.genblk1[45].entry.input_buf[1].A ;
 wire \l_fifo.genblk1[45].entry.input_buf[1].X ;
 wire \l_fifo.genblk1[45].entry.input_buf[1].genblk1[0].mid ;
 wire \l_fifo.genblk1[45].entry.input_buf[2].A ;
 wire \l_fifo.genblk1[45].entry.input_buf[2].X ;
 wire \l_fifo.genblk1[45].entry.input_buf[2].genblk1[0].mid ;
 wire \l_fifo.genblk1[45].entry.input_buf[3].A ;
 wire \l_fifo.genblk1[45].entry.input_buf[3].X ;
 wire \l_fifo.genblk1[45].entry.input_buf[3].genblk1[0].mid ;
 wire \l_fifo.genblk1[45].entry.input_buf[4].A ;
 wire \l_fifo.genblk1[45].entry.input_buf[4].X ;
 wire \l_fifo.genblk1[45].entry.input_buf[4].genblk1[0].mid ;
 wire \l_fifo.genblk1[45].entry.input_buf[5].A ;
 wire \l_fifo.genblk1[45].entry.input_buf[5].X ;
 wire \l_fifo.genblk1[45].entry.input_buf[5].genblk1[0].mid ;
 wire \l_fifo.genblk1[46].entry.empty ;
 wire \l_fifo.genblk1[46].entry.input_buf[0].A ;
 wire \l_fifo.genblk1[46].entry.input_buf[0].X ;
 wire \l_fifo.genblk1[46].entry.input_buf[0].genblk1[0].mid ;
 wire \l_fifo.genblk1[46].entry.input_buf[1].A ;
 wire \l_fifo.genblk1[46].entry.input_buf[1].X ;
 wire \l_fifo.genblk1[46].entry.input_buf[1].genblk1[0].mid ;
 wire \l_fifo.genblk1[46].entry.input_buf[2].A ;
 wire \l_fifo.genblk1[46].entry.input_buf[2].X ;
 wire \l_fifo.genblk1[46].entry.input_buf[2].genblk1[0].mid ;
 wire \l_fifo.genblk1[46].entry.input_buf[3].A ;
 wire \l_fifo.genblk1[46].entry.input_buf[3].X ;
 wire \l_fifo.genblk1[46].entry.input_buf[3].genblk1[0].mid ;
 wire \l_fifo.genblk1[46].entry.input_buf[4].A ;
 wire \l_fifo.genblk1[46].entry.input_buf[4].X ;
 wire \l_fifo.genblk1[46].entry.input_buf[4].genblk1[0].mid ;
 wire \l_fifo.genblk1[46].entry.input_buf[5].A ;
 wire \l_fifo.genblk1[46].entry.input_buf[5].X ;
 wire \l_fifo.genblk1[46].entry.input_buf[5].genblk1[0].mid ;
 wire \l_fifo.genblk1[47].entry.empty ;
 wire \l_fifo.genblk1[47].entry.input_buf[0].X ;
 wire \l_fifo.genblk1[47].entry.input_buf[0].genblk1[0].mid ;
 wire \l_fifo.genblk1[47].entry.input_buf[1].X ;
 wire \l_fifo.genblk1[47].entry.input_buf[1].genblk1[0].mid ;
 wire \l_fifo.genblk1[47].entry.input_buf[2].X ;
 wire \l_fifo.genblk1[47].entry.input_buf[2].genblk1[0].mid ;
 wire \l_fifo.genblk1[47].entry.input_buf[3].X ;
 wire \l_fifo.genblk1[47].entry.input_buf[3].genblk1[0].mid ;
 wire \l_fifo.genblk1[47].entry.input_buf[4].X ;
 wire \l_fifo.genblk1[47].entry.input_buf[4].genblk1[0].mid ;
 wire \l_fifo.genblk1[47].entry.input_buf[5].X ;
 wire \l_fifo.genblk1[47].entry.input_buf[5].genblk1[0].mid ;
 wire \l_fifo.genblk1[47].entry.write_in ;
 wire \l_fifo.genblk1[4].entry.empty ;
 wire \l_fifo.genblk1[4].entry.input_buf[0].A ;
 wire \l_fifo.genblk1[4].entry.input_buf[0].X ;
 wire \l_fifo.genblk1[4].entry.input_buf[0].genblk1[0].mid ;
 wire \l_fifo.genblk1[4].entry.input_buf[1].A ;
 wire \l_fifo.genblk1[4].entry.input_buf[1].X ;
 wire \l_fifo.genblk1[4].entry.input_buf[1].genblk1[0].mid ;
 wire \l_fifo.genblk1[4].entry.input_buf[2].A ;
 wire \l_fifo.genblk1[4].entry.input_buf[2].X ;
 wire \l_fifo.genblk1[4].entry.input_buf[2].genblk1[0].mid ;
 wire \l_fifo.genblk1[4].entry.input_buf[3].A ;
 wire \l_fifo.genblk1[4].entry.input_buf[3].X ;
 wire \l_fifo.genblk1[4].entry.input_buf[3].genblk1[0].mid ;
 wire \l_fifo.genblk1[4].entry.input_buf[4].A ;
 wire \l_fifo.genblk1[4].entry.input_buf[4].X ;
 wire \l_fifo.genblk1[4].entry.input_buf[4].genblk1[0].mid ;
 wire \l_fifo.genblk1[4].entry.input_buf[5].A ;
 wire \l_fifo.genblk1[4].entry.input_buf[5].X ;
 wire \l_fifo.genblk1[4].entry.input_buf[5].genblk1[0].mid ;
 wire \l_fifo.genblk1[5].entry.empty ;
 wire \l_fifo.genblk1[5].entry.input_buf[0].A ;
 wire \l_fifo.genblk1[5].entry.input_buf[0].X ;
 wire \l_fifo.genblk1[5].entry.input_buf[0].genblk1[0].mid ;
 wire \l_fifo.genblk1[5].entry.input_buf[1].A ;
 wire \l_fifo.genblk1[5].entry.input_buf[1].X ;
 wire \l_fifo.genblk1[5].entry.input_buf[1].genblk1[0].mid ;
 wire \l_fifo.genblk1[5].entry.input_buf[2].A ;
 wire \l_fifo.genblk1[5].entry.input_buf[2].X ;
 wire \l_fifo.genblk1[5].entry.input_buf[2].genblk1[0].mid ;
 wire \l_fifo.genblk1[5].entry.input_buf[3].A ;
 wire \l_fifo.genblk1[5].entry.input_buf[3].X ;
 wire \l_fifo.genblk1[5].entry.input_buf[3].genblk1[0].mid ;
 wire \l_fifo.genblk1[5].entry.input_buf[4].A ;
 wire \l_fifo.genblk1[5].entry.input_buf[4].X ;
 wire \l_fifo.genblk1[5].entry.input_buf[4].genblk1[0].mid ;
 wire \l_fifo.genblk1[5].entry.input_buf[5].A ;
 wire \l_fifo.genblk1[5].entry.input_buf[5].X ;
 wire \l_fifo.genblk1[5].entry.input_buf[5].genblk1[0].mid ;
 wire \l_fifo.genblk1[6].entry.empty ;
 wire \l_fifo.genblk1[6].entry.input_buf[0].A ;
 wire \l_fifo.genblk1[6].entry.input_buf[0].X ;
 wire \l_fifo.genblk1[6].entry.input_buf[0].genblk1[0].mid ;
 wire \l_fifo.genblk1[6].entry.input_buf[1].A ;
 wire \l_fifo.genblk1[6].entry.input_buf[1].X ;
 wire \l_fifo.genblk1[6].entry.input_buf[1].genblk1[0].mid ;
 wire \l_fifo.genblk1[6].entry.input_buf[2].A ;
 wire \l_fifo.genblk1[6].entry.input_buf[2].X ;
 wire \l_fifo.genblk1[6].entry.input_buf[2].genblk1[0].mid ;
 wire \l_fifo.genblk1[6].entry.input_buf[3].A ;
 wire \l_fifo.genblk1[6].entry.input_buf[3].X ;
 wire \l_fifo.genblk1[6].entry.input_buf[3].genblk1[0].mid ;
 wire \l_fifo.genblk1[6].entry.input_buf[4].A ;
 wire \l_fifo.genblk1[6].entry.input_buf[4].X ;
 wire \l_fifo.genblk1[6].entry.input_buf[4].genblk1[0].mid ;
 wire \l_fifo.genblk1[6].entry.input_buf[5].A ;
 wire \l_fifo.genblk1[6].entry.input_buf[5].X ;
 wire \l_fifo.genblk1[6].entry.input_buf[5].genblk1[0].mid ;
 wire \l_fifo.genblk1[7].entry.empty ;
 wire \l_fifo.genblk1[7].entry.input_buf[0].A ;
 wire \l_fifo.genblk1[7].entry.input_buf[0].X ;
 wire \l_fifo.genblk1[7].entry.input_buf[0].genblk1[0].mid ;
 wire \l_fifo.genblk1[7].entry.input_buf[1].A ;
 wire \l_fifo.genblk1[7].entry.input_buf[1].X ;
 wire \l_fifo.genblk1[7].entry.input_buf[1].genblk1[0].mid ;
 wire \l_fifo.genblk1[7].entry.input_buf[2].A ;
 wire \l_fifo.genblk1[7].entry.input_buf[2].X ;
 wire \l_fifo.genblk1[7].entry.input_buf[2].genblk1[0].mid ;
 wire \l_fifo.genblk1[7].entry.input_buf[3].A ;
 wire \l_fifo.genblk1[7].entry.input_buf[3].X ;
 wire \l_fifo.genblk1[7].entry.input_buf[3].genblk1[0].mid ;
 wire \l_fifo.genblk1[7].entry.input_buf[4].A ;
 wire \l_fifo.genblk1[7].entry.input_buf[4].X ;
 wire \l_fifo.genblk1[7].entry.input_buf[4].genblk1[0].mid ;
 wire \l_fifo.genblk1[7].entry.input_buf[5].A ;
 wire \l_fifo.genblk1[7].entry.input_buf[5].X ;
 wire \l_fifo.genblk1[7].entry.input_buf[5].genblk1[0].mid ;
 wire \l_fifo.genblk1[8].entry.empty ;
 wire \l_fifo.genblk1[8].entry.input_buf[0].A ;
 wire \l_fifo.genblk1[8].entry.input_buf[0].X ;
 wire \l_fifo.genblk1[8].entry.input_buf[0].genblk1[0].mid ;
 wire \l_fifo.genblk1[8].entry.input_buf[1].A ;
 wire \l_fifo.genblk1[8].entry.input_buf[1].X ;
 wire \l_fifo.genblk1[8].entry.input_buf[1].genblk1[0].mid ;
 wire \l_fifo.genblk1[8].entry.input_buf[2].A ;
 wire \l_fifo.genblk1[8].entry.input_buf[2].X ;
 wire \l_fifo.genblk1[8].entry.input_buf[2].genblk1[0].mid ;
 wire \l_fifo.genblk1[8].entry.input_buf[3].A ;
 wire \l_fifo.genblk1[8].entry.input_buf[3].X ;
 wire \l_fifo.genblk1[8].entry.input_buf[3].genblk1[0].mid ;
 wire \l_fifo.genblk1[8].entry.input_buf[4].A ;
 wire \l_fifo.genblk1[8].entry.input_buf[4].X ;
 wire \l_fifo.genblk1[8].entry.input_buf[4].genblk1[0].mid ;
 wire \l_fifo.genblk1[8].entry.input_buf[5].A ;
 wire \l_fifo.genblk1[8].entry.input_buf[5].X ;
 wire \l_fifo.genblk1[8].entry.input_buf[5].genblk1[0].mid ;
 wire \l_fifo.genblk1[9].entry.input_buf[0].A ;
 wire \l_fifo.genblk1[9].entry.input_buf[0].X ;
 wire \l_fifo.genblk1[9].entry.input_buf[0].genblk1[0].mid ;
 wire \l_fifo.genblk1[9].entry.input_buf[1].A ;
 wire \l_fifo.genblk1[9].entry.input_buf[1].X ;
 wire \l_fifo.genblk1[9].entry.input_buf[1].genblk1[0].mid ;
 wire \l_fifo.genblk1[9].entry.input_buf[2].A ;
 wire \l_fifo.genblk1[9].entry.input_buf[2].X ;
 wire \l_fifo.genblk1[9].entry.input_buf[2].genblk1[0].mid ;
 wire \l_fifo.genblk1[9].entry.input_buf[3].A ;
 wire \l_fifo.genblk1[9].entry.input_buf[3].X ;
 wire \l_fifo.genblk1[9].entry.input_buf[3].genblk1[0].mid ;
 wire \l_fifo.genblk1[9].entry.input_buf[4].A ;
 wire \l_fifo.genblk1[9].entry.input_buf[4].X ;
 wire \l_fifo.genblk1[9].entry.input_buf[4].genblk1[0].mid ;
 wire \l_fifo.genblk1[9].entry.input_buf[5].A ;
 wire \l_fifo.genblk1[9].entry.input_buf[5].X ;
 wire \l_fifo.genblk1[9].entry.input_buf[5].genblk1[0].mid ;
 wire \l_fifo.ready ;
 wire net1;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net2;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net3;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net4;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire reset_n_in;
 wire [0:0] clknet_0_io_in;
 wire [0:0] clknet_3_0__leaf_io_in;
 wire [0:0] clknet_3_1__leaf_io_in;
 wire [0:0] clknet_3_2__leaf_io_in;
 wire [0:0] clknet_3_3__leaf_io_in;
 wire [0:0] clknet_3_4__leaf_io_in;
 wire [0:0] clknet_3_5__leaf_io_in;
 wire [0:0] clknet_3_6__leaf_io_in;
 wire [0:0] clknet_3_7__leaf_io_in;

 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(_000_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_10 (.DIODE(\l_fifo.genblk1[14].entry.input_buf[0].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_11 (.DIODE(\l_fifo.genblk1[17].entry.input_buf[2].X ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_12 (.DIODE(\l_fifo.genblk1[3].entry.input_buf[3].X ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(_002_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_3 (.DIODE(_010_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_4 (.DIODE(_024_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_5 (.DIODE(_082_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_6 (.DIODE(\data_in_buffer[5].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_7 (.DIODE(\l_fifo.genblk1[18].entry.input_buf[2].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_8 (.DIODE(_053_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_9 (.DIODE(\data_in_buffer[0].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_0_106 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_113 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_119 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_0_131 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_139 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_141 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_153 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_165 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_0_169 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_179 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_0_187 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_195 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_197 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_0_203 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_209 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_0_21 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_214 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_221 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_225 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_237 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_249 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_253 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_265 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_27 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_277 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_281 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_29 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_0_293 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_0_47 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_55 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_57 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_69 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_81 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_85 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_97 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_10_103 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_10_118 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_10_131 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_10_138 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_10_141 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_10_150 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_10_161 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_10_170 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_10_179 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_10_187 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_10_194 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_10_197 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_10_212 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_10_220 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_10_24 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_10_241 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_10_248 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_10_253 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_10_258 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_10_265 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_10_272 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_10_279 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_10_286 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_10_29 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_10_293 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_10_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_10_50 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_10_58 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_10_78 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_10_85 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_11_107 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_11_111 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_11_113 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_11_123 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_11_127 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_11_131 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_11_140 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_11_147 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_11_15 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_11_159 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_11_166 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_11_169 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_11_184 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_11_201 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_11_218 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_11_225 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_11_240 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_11_247 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_11_259 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_11_266 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_11_273 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_11_279 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_11_281 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_11_285 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_11_289 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_11_293 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_11_297 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_11_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_11_36 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_11_48 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_11_57 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_11_63 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_11_81 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_11_85 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_11_89 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_11_96 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_12_108 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_12_121 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_12_129 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_12_138 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_12_141 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_12_154 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_12_163 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_12_174 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_12_181 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_12_188 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_12_197 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_12_209 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_12_216 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_12_22 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_12_223 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_12_230 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_12_247 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_12_251 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_12_253 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_12_268 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_12_275 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_12_282 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_12_289 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_12_29 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_12_293 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_12_297 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_12_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_12_34 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_12_42 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_12_65 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_12_77 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_12_82 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_12_85 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_12_91 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_12_99 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_13_109 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_13_11 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_13_113 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_13_121 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_13_125 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_13_132 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_13_139 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_13_150 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_13_156 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_13_164 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_13_169 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_13_179 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_13_200 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_13_208 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_13_222 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_13_225 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_13_240 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_13_244 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_13_249 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_13_256 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_13_263 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_13_271 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_13_278 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_13_281 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_13_286 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_13_297 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_13_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_13_30 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_13_51 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_13_55 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_13_57 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_13_77 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_13_97 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_14_103 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_14_113 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_14_123 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_14_132 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_14_141 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_14_150 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_14_157 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_14_165 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_14_180 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_14_188 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_14_197 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_14_213 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_14_220 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_14_228 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_14_233 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_14_240 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_14_247 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_14_251 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_14_253 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_14_26 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_14_274 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_14_281 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_14_288 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_14_29 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_14_295 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_14_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_14_35 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_14_53 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_14_59 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_14_76 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_14_85 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_15_110 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_15_113 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_15_122 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_15_131 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_15_135 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_15_143 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_15_147 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_15_153 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_15_164 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_15_169 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_15_176 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_15_193 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_15_200 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_15_207 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_15_21 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_15_214 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_15_221 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_15_225 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_15_230 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_15_237 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_15_244 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_15_255 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_15_261 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_15_265 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_15_274 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_15_281 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_15_286 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_15_293 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_15_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_15_42 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_15_54 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_15_57 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_15_77 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_15_97 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_16_108 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_16_116 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_16_122 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_16_133 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_16_139 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_16_141 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_16_155 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_16_172 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_16_188 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_16_197 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_16_202 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_16_208 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_16_212 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_16_22 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_16_229 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_16_246 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_16_253 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_16_268 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_16_276 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_16_281 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_16_288 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_16_29 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_16_292 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_16_296 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_16_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_16_48 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_16_57 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_16_78 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_16_85 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_16_93 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_17_100 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_17_106 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_17_110 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_17_113 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_17_121 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_17_129 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_17_141 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_17_148 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_17_152 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_17_159 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_17_166 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_17_169 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_17_176 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_17_193 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_17_197 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_17_211 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_17_218 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_17_225 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_17_232 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_17_240 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_17_247 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_17_254 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_17_261 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_17_278 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_17_281 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_17_287 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_17_293 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_17_297 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_17_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_17_36 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_17_47 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_17_54 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_17_57 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_17_8 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_17_80 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_18_102 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_18_112 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_18_121 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_18_129 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_18_138 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_18_141 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_18_152 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_18_161 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_18_168 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_18_187 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_18_194 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_18_197 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_18_202 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_18_209 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_18_228 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_18_24 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_18_245 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_18_251 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_18_253 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_18_268 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_18_275 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_18_283 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_18_29 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_18_297 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_18_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_18_33 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_18_36 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_18_55 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_18_76 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_18_85 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_18_91 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_19_104 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_19_113 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_19_119 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_19_126 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_19_134 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_19_141 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_19_145 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_19_151 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_19_157 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_19_16 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_19_166 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_19_169 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_19_184 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_19_188 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_19_202 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_19_219 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_19_223 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_19_225 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_19_244 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_19_261 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_19_278 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_19_281 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_19_286 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_19_293 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_19_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_19_34 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_19_54 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_19_57 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_19_76 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_19_8 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_19_80 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_19_84 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_19_93 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_1_102 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_1_109 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_1_113 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_1_118 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_1_128 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_1_135 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_1_139 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_1_143 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_1_160 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_1_169 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_1_184 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_1_201 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_1_205 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_1_219 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_1_223 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_1_225 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_1_23 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_1_230 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_1_239 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_1_251 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_1_263 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_1_275 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_1_279 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_1_281 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_1_293 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_1_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_1_43 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_1_55 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_1_57 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_1_63 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_1_81 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_20_103 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_20_110 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_20_117 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_20_126 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_20_138 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_20_141 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_20_152 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_20_162 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_20_169 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_20_190 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_20_197 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_20_202 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_20_209 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_20_230 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_20_237 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_20_241 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_20_246 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_20_253 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_20_259 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_20_26 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_20_273 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_20_281 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_20_288 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_20_29 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_20_295 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_20_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_20_41 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_20_67 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_20_71 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_20_75 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_20_82 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_20_85 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_20_9 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_21_106 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_21_113 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_21_123 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_21_132 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_21_136 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_21_140 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_21_151 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_21_160 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_21_169 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_21_184 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_21_192 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_21_199 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_21_206 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_21_213 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_21_217 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_21_222 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_21_225 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_21_231 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_21_248 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_21_265 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_21_27 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_21_272 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_21_281 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_21_296 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_21_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_21_34 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_21_54 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_21_57 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_21_76 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_21_84 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_21_88 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_21_9 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_21_97 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_22_101 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_22_106 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_22_117 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_22_121 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_22_126 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_22_138 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_22_141 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_22_148 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_22_157 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_22_163 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_22_167 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_22_179 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_22_186 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_22_194 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_22_197 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_22_218 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_22_22 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_22_224 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_22_238 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_22_246 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_22_253 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_22_258 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_22_265 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_22_272 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_22_279 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_22_287 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_22_29 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_22_294 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_22_298 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_22_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_22_41 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_22_65 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_22_74 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_22_82 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_22_85 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_22_91 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_22_97 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_23_101 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_23_110 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_23_113 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_23_120 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_23_135 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_23_144 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_23_150 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_23_154 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_23_163 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_23_167 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_23_169 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_23_188 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_23_192 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_23_206 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_23_213 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_23_220 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_23_225 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_23_23 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_23_235 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_23_247 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_23_254 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_23_262 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_23_276 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_23_281 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_23_286 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_23_293 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_23_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_23_43 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_23_50 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_23_57 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_23_76 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_23_85 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_23_94 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_24_100 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_24_111 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_24_119 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_24_131 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_24_138 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_24_141 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_24_152 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_24_161 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_24_178 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_24_186 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_24_193 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_24_197 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_24_212 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_24_219 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_24_226 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_24_23 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_24_233 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_24_250 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_24_253 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_24_269 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_24_27 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_24_29 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_24_290 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_24_297 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_24_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_24_48 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_24_55 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_24_80 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_24_85 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_25_101 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_25_110 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_25_113 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_25_117 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_25_131 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_25_139 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_25_144 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_25_152 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_25_166 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_25_169 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_25_188 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_25_205 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_25_222 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_25_225 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_25_231 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_25_25 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_25_252 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_25_259 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_25_267 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_25_274 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_25_281 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_25_286 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_25_29 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_25_293 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_25_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_25_34 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_25_54 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_25_57 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_25_63 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_25_7 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_25_81 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_26_105 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_26_113 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_26_128 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_26_134 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_26_138 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_26_141 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_26_148 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_26_152 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_26_157 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_26_166 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_26_174 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_26_181 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_26_188 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_26_197 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_26_203 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_26_217 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_26_23 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_26_238 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_26_246 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_26_253 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_26_258 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_26_266 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_26_27 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_26_280 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_26_288 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_26_29 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_26_296 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_26_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_26_34 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_26_41 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_26_65 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_26_72 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_26_79 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_26_83 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_26_85 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_26_89 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_26_93 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_27_110 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_27_113 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_27_119 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_27_12 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_27_133 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_27_141 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_27_155 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_27_163 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_27_167 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_27_169 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_27_188 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_27_195 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_27_199 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_27_210 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_27_217 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_27_223 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_27_225 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_27_229 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_27_240 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_27_244 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_27_258 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_27_275 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_27_279 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_27_281 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_27_296 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_27_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_27_36 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_27_44 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_27_49 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_27_55 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_27_57 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_27_76 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_27_84 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_27_88 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_27_98 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_28_109 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_28_117 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_28_129 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_28_138 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_28_141 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_28_147 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_28_161 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_28_178 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_28_186 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_28_193 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_28_197 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_28_214 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_28_218 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_28_232 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_28_249 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_28_25 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_28_253 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_28_268 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_28_275 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_28_283 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_28_29 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_28_297 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_28_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_28_49 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_28_7 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_28_70 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_28_78 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_28_82 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_28_85 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_28_91 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_28_98 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_29_104 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_29_113 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_29_123 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_29_131 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_29_137 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_29_142 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_29_150 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_29_158 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_29_166 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_29_169 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_29_181 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_29_202 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_29_209 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_29_216 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_29_22 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_29_225 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_29_229 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_29_234 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_29_241 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_29_245 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_29_250 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_29_257 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_29_264 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_29_271 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_29_278 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_29_281 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_29_287 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_29_294 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_29_298 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_29_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_29_43 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_29_50 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_29_57 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_29_63 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_29_74 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_29_79 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_29_83 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_29_88 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_29_95 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_2_109 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_2_117 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_2_123 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_2_129 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_2_137 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_2_141 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_2_153 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_2_162 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_2_169 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_2_180 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_2_187 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_2_194 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_2_197 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_2_202 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_2_209 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_2_216 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_2_22 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_2_228 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_2_235 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_2_242 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_2_250 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_2_253 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_2_265 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_2_277 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_2_289 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_2_29 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_2_297 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_2_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_2_41 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_2_61 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_2_82 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_2_85 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_2_97 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_30_104 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_30_111 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_30_121 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_30_138 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_30_141 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_30_156 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_30_160 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_30_174 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_30_180 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_30_194 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_30_197 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_30_203 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_30_217 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_30_22 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_30_234 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_30_241 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_30_248 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_30_253 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_30_259 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_30_267 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_30_274 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_30_282 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_30_29 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_30_297 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_30_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_30_34 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_30_41 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_30_48 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_30_59 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_30_82 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_30_85 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_30_91 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_30_95 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_31_103 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_31_110 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_31_113 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_31_122 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_31_129 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_31_136 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_31_153 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_31_164 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_31_169 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_31_186 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_31_193 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_31_210 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_31_217 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_31_223 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_31_225 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_31_240 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_31_257 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_31_27 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_31_274 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_31_281 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_31_296 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_31_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_31_38 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_31_45 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_31_52 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_31_57 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_31_77 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_31_85 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_31_89 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_31_9 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_31_96 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_32_100 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_32_111 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_32_115 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_32_123 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_32_127 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_32_131 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_32_138 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_32_141 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_32_146 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_32_153 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_32_170 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_32_177 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_32_194 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_32_197 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_32_202 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_32_209 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_32_216 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_32_22 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_32_223 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_32_230 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_32_237 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_32_244 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_32_253 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_32_268 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_32_285 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_32_29 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_32_293 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_32_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_32_35 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_32_44 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_32_59 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_32_79 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_32_83 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_32_85 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_32_89 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_32_93 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_33_103 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_33_11 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_33_110 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_33_113 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_33_129 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_33_146 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_33_152 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_33_166 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_33_169 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_33_174 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_33_18 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_33_182 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_33_190 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_33_197 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_33_205 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_33_222 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_33_225 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_33_240 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_33_25 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_33_257 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_33_275 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_33_279 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_33_281 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_33_287 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_33_291 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_33_296 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_33_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_33_50 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_33_57 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_33_64 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_33_7 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_33_71 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_33_82 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_33_89 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_33_96 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_34_101 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_34_112 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_34_121 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_34_138 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_34_141 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_34_157 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_34_165 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_34_186 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_34_194 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_34_197 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_34_213 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_34_220 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_34_227 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_34_23 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_34_233 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_34_238 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_34_245 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_34_251 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_34_253 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_34_268 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_34_27 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_34_276 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_34_29 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_34_297 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_34_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_34_34 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_34_41 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_34_52 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_34_64 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_34_71 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_34_82 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_34_85 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_35_10 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_35_108 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_35_113 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_35_119 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_35_123 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_35_127 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_35_134 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_35_141 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_35_145 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_35_149 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_35_166 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_35_169 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_35_188 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_35_19 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_35_205 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_35_213 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_35_217 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_35_222 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_35_225 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_35_240 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_35_247 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_35_26 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_35_264 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_35_276 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_35_281 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_35_296 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_35_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_35_32 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_35_36 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_35_43 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_35_49 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_35_53 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_35_57 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_35_76 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_35_87 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_36_101 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_36_115 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_36_132 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_36_141 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_36_145 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_36_159 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_36_163 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_36_17 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_36_177 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_36_184 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_36_188 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_36_193 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_36_197 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_36_202 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_36_219 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_36_236 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_36_240 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_36_244 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_36_253 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_36_259 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_36_26 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_36_265 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_36_279 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_36_287 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_36_29 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_36_294 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_36_298 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_36_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_36_39 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_36_45 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_36_49 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_36_56 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_36_63 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_36_72 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_36_8 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_36_82 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_36_85 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_36_97 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_37_104 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_37_113 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_37_124 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_37_141 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_37_145 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_37_159 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_37_166 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_37_169 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_37_188 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_37_20 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_37_200 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_37_207 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_37_214 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_37_222 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_37_225 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_37_230 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_37_249 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_37_255 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_37_269 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_37_276 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_37_28 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_37_281 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_37_296 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_37_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_37_33 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_37_40 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_37_47 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_37_54 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_37_57 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_37_65 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_37_76 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_37_86 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_37_9 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_37_93 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_38_100 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_38_109 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_38_11 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_38_117 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_38_124 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_38_131 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_38_138 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_38_141 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_38_145 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_38_15 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_38_150 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_38_158 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_38_166 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_38_171 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_38_177 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_38_182 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_38_189 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_38_19 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_38_195 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_38_197 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_38_212 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_38_229 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_38_241 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_38_248 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_38_253 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_38_26 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_38_268 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_38_285 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_38_29 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_38_292 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_38_298 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_38_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_38_38 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_38_44 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_38_49 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_38_56 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_38_63 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_38_74 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_38_82 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_38_85 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_39_106 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_39_113 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_39_128 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_39_149 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_39_157 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_39_162 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_39_169 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_39_184 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_39_191 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_39_195 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_39_209 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_39_22 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_39_221 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_39_225 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_39_244 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_39_252 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_39_260 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_39_264 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_39_278 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_39_281 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_39_293 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_39_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_39_34 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_39_54 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_39_57 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_39_64 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_39_79 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_39_89 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_39_9 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_39_98 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_3_109 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_3_113 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_3_119 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_3_128 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_3_135 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_3_139 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_3_145 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_3_157 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_3_166 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_3_169 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_3_182 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_3_190 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_3_204 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_3_221 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_3_225 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_3_240 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_3_247 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_3_259 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_3_27 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_3_271 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_3_279 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_3_281 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_3_293 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_3_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_3_47 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_3_55 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_3_57 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_3_65 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_3_85 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_3_9 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_3_93 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_3_97 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_40_10 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_40_109 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_40_113 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_40_117 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_40_134 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_40_141 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_40_160 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_40_168 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_40_172 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_40_177 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_40_194 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_40_197 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_40_202 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_40_206 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_40_21 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_40_220 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_40_237 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_40_241 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_40_246 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_40_253 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_40_268 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_40_27 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_40_276 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_40_29 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_40_297 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_40_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_40_41 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_40_53 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_40_61 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_40_75 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_40_82 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_40_85 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_40_92 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_41_100 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_41_109 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_41_113 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_41_129 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_41_146 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_41_15 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_41_154 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_41_166 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_41_169 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_41_184 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_41_201 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_41_208 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_41_215 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_41_222 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_41_225 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_41_242 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_41_259 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_41_26 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_41_266 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_41_273 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_41_279 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_41_281 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_41_287 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_41_294 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_41_298 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_41_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_41_32 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_41_36 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_41_47 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_41_54 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_41_57 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_41_66 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_41_81 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_41_9 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_41_92 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_42_100 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_42_107 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_42_124 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_42_13 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_42_132 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_42_141 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_42_148 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_42_155 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_42_163 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_42_180 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_42_187 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_42_194 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_42_197 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_42_21 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_42_212 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_42_220 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_42_227 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_42_248 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_42_253 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_42_259 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_42_26 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_42_265 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_42_279 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_42_29 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_42_296 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_42_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_42_38 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_42_50 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_42_54 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_42_58 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_42_65 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_42_82 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_42_85 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_43_110 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_43_113 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_43_125 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_43_13 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_43_133 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_43_148 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_43_165 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_43_169 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_43_184 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_43_201 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_43_22 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_43_222 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_43_225 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_43_230 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_43_238 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_43_243 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_43_251 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_43_258 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_43_265 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_43_272 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_43_281 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_43_286 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_43_293 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_43_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_43_30 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_43_37 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_43_43 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_43_47 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_43_54 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_43_57 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_43_67 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_43_71 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_43_76 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_43_9 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_43_93 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_44_10 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_44_103 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_44_107 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_44_118 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_44_135 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_44_139 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_44_141 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_44_146 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_44_154 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_44_166 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_44_174 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_44_181 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_44_19 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_44_193 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_44_197 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_44_212 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_44_229 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_44_246 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_44_253 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_44_26 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_44_268 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_44_276 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_44_284 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_44_29 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_44_291 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_44_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_44_36 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_44_43 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_44_50 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_44_57 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_44_74 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_44_78 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_44_82 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_44_85 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_44_95 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_45_101 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_45_110 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_45_113 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_45_120 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_45_13 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_45_137 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_45_154 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_45_161 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_45_167 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_45_169 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_45_177 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_45_18 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_45_194 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_45_211 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_45_219 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_45_22 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_45_223 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_45_225 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_45_230 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_45_251 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_45_258 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_45_264 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_45_27 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_45_278 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_45_281 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_45_296 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_45_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_45_34 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_45_45 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_45_54 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_45_57 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_45_65 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_45_69 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_45_83 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_45_87 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_45_9 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_46_105 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_46_12 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_46_122 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_46_131 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_46_138 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_46_141 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_46_147 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_46_161 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_46_178 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_46_185 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_46_19 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_46_192 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_46_197 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_46_212 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_46_220 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_46_235 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_46_242 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_46_249 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_46_253 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_46_258 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_46_26 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_46_265 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_46_272 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_46_279 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_46_286 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_46_29 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_46_293 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_46_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_46_44 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_46_63 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_46_74 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_46_78 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_46_82 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_46_85 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_46_91 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_47_105 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_47_110 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_47_113 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_47_119 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_47_133 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_47_15 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_47_150 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_47_156 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_47_161 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_47_167 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_47_169 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_47_174 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_47_181 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_47_190 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_47_197 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_47_204 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_47_208 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_47_22 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_47_222 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_47_225 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_47_230 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_47_237 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_47_244 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_47_250 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_47_264 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_47_272 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_47_281 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_47_29 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_47_297 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_47_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_47_36 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_47_53 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_47_57 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_47_65 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_47_73 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_47_8 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_47_80 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_47_97 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_48_100 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_48_108 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_48_112 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_48_12 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_48_129 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_48_138 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_48_141 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_48_147 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_48_164 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_48_185 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_48_19 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_48_192 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_48_197 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_48_203 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_48_209 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_48_223 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_48_227 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_48_232 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_48_249 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_48_253 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_48_26 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_48_269 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_48_286 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_48_29 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_48_293 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_48_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_48_35 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_48_46 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_48_54 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_48_71 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_48_82 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_48_85 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_49_109 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_49_113 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_49_132 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_49_149 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_49_15 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_49_155 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_49_159 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_49_166 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_49_169 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_49_184 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_49_201 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_49_218 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_49_22 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_49_225 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_49_230 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_49_237 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_49_258 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_49_265 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_49_275 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_49_279 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_49_281 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_49_286 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_49_293 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_49_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_49_31 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_49_39 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_49_54 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_49_57 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_49_78 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_49_8 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_49_82 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_49_87 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_49_95 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_4_103 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_4_114 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_4_127 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_4_138 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_4_141 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_4_145 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_4_154 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_4_171 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_4_179 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_4_184 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_4_191 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_4_195 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_4_197 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_4_216 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_4_224 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_4_239 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_4_246 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_4_253 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_4_26 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_4_265 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_4_277 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_4_289 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_4_29 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_4_297 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_4_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_4_48 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_4_60 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_4_78 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_4_85 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_50_100 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_50_119 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_50_12 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_50_123 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_50_127 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_50_138 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_50_141 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_50_146 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_50_152 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_50_156 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_50_173 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_50_194 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_50_197 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_50_20 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_50_202 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_50_208 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_50_213 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_50_230 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_50_247 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_50_251 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_50_253 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_50_258 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_50_265 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_50_272 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_50_279 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_50_286 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_50_29 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_50_293 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_50_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_50_44 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_50_52 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_50_61 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_50_68 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_50_75 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_50_82 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_50_85 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_51_105 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_51_111 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_51_113 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_51_117 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_51_121 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_51_128 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_51_138 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_51_155 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_51_162 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_51_169 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_51_175 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_51_183 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_51_191 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_51_208 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_51_216 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_51_225 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_51_230 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_51_238 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_51_24 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_51_243 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_51_248 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_51_252 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_51_267 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_51_274 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_51_281 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_51_296 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_51_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_51_32 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_51_46 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_51_50 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_51_54 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_51_57 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_51_63 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_51_71 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_51_77 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_51_81 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_51_88 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_51_96 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_52_100 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_52_117 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_52_12 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_52_138 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_52_141 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_52_157 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_52_174 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_52_19 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_52_191 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_52_195 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_52_197 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_52_203 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_52_207 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_52_221 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_52_229 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_52_244 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_52_253 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_52_26 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_52_268 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_52_285 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_52_29 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_52_292 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_52_298 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_52_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_52_48 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_52_65 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_52_82 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_52_85 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_53_102 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_53_109 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_53_113 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_53_117 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_53_121 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_53_128 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_53_136 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_53_143 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_53_15 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_53_151 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_53_155 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_53_166 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_53_169 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_53_174 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_53_180 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_53_185 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_53_204 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_53_218 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_53_225 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_53_230 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_53_251 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_53_258 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_53_265 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_53_272 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_53_281 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_53_286 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_53_290 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_53_294 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_53_298 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_53_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_53_30 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_53_34 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_53_49 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_53_55 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_53_57 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_53_67 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_53_78 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_53_8 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_53_85 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_54_112 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_54_12 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_54_129 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_54_136 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_54_141 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_54_147 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_54_156 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_54_173 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_54_180 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_54_187 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_54_19 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_54_194 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_54_197 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_54_205 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_54_212 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_54_219 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_54_236 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_54_244 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_54_253 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_54_259 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_54_26 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_54_266 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_54_273 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_54_280 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_54_287 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_54_29 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_54_294 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_54_298 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_54_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_54_35 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_54_52 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_54_58 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_54_63 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_54_71 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_54_82 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_54_85 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_54_95 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_55_106 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_55_110 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_55_113 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_55_119 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_55_123 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_55_14 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_55_140 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_55_154 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_55_162 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_55_166 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_55_169 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_55_174 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_55_18 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_55_191 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_55_212 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_55_219 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_55_223 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_55_225 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_55_23 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_55_240 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_55_247 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_55_254 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_55_261 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_55_268 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_55_275 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_55_279 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_55_281 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_55_286 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_55_293 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_55_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_55_30 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_55_37 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_55_45 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_55_54 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_55_57 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_55_72 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_55_83 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_55_9 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_55_90 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_55_98 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_56_100 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_56_12 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_56_121 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_56_138 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_56_141 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_56_157 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_56_174 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_56_19 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_56_191 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_56_195 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_56_197 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_56_212 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_56_229 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_56_236 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_56_243 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_56_250 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_56_253 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_56_26 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_56_268 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_56_275 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_56_282 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_56_29 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_56_291 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_56_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_56_48 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_56_65 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_56_82 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_56_85 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_57_103 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_57_110 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_57_113 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_57_119 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_57_12 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_57_123 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_57_127 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_57_131 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_57_138 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_57_141 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_57_145 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_57_149 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_57_156 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_57_163 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_57_167 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_57_169 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_57_176 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_57_184 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_57_19 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_57_190 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_57_197 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_57_202 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_57_209 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_57_218 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_57_225 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_57_230 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_57_237 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_57_244 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_57_253 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_57_258 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_57_26 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_57_265 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_57_272 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_57_281 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_57_286 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_57_29 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_57_293 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_57_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_57_33 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_57_37 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_57_45 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_57_54 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_57_57 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_57_67 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_57_71 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_57_75 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_57_82 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_57_85 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_57_96 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_5_100 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_5_104 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_5_11 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_5_110 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_5_113 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_5_124 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_5_128 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_5_136 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_5_14 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_5_147 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_5_154 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_5_158 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_5_166 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_5_169 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_5_184 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_5_201 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_5_208 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_5_215 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_5_222 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_5_225 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_5_230 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_5_237 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_5_244 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_5_251 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_5_258 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_5_265 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_5_272 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_5_281 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_5_293 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_5_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_5_33 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_5_54 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_5_57 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_5_80 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_6_109 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_6_120 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_6_131 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_6_138 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_6_141 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_6_147 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_6_158 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_6_166 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_6_173 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_6_184 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_6_193 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_6_197 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_6_201 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_6_21 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_6_215 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_6_222 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_6_230 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_6_244 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_6_253 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_6_258 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_6_265 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_6_27 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_6_272 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_6_284 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_6_29 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_6_296 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_6_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_6_47 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_6_59 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_6_76 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_6_85 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_6_91 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_6_98 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_7_110 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_7_113 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_7_120 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_7_129 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_7_140 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_7_149 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_7_15 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_7_153 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_7_161 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_7_167 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_7_169 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_7_184 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_7_188 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_7_193 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_7_199 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_7_203 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_7_210 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_7_217 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_7_223 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_7_225 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_7_231 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_7_235 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_7_240 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_7_257 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_7_264 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_7_271 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_7_278 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_7_281 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_7_286 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_7_298 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_7_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_7_36 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_7_48 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_7_57 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_7_78 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_7_86 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_7_9 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_7_90 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_7_99 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_8_110 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_8_124 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_8_135 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_8_139 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_8_141 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_8_150 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_8_163 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_8_180 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_8_188 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_8_197 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_8_212 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_8_22 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_8_229 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_8_233 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_8_247 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_8_251 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_8_253 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_8_258 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_8_265 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_8_272 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_8_281 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_8_288 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_8_29 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_8_295 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_8_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_8_41 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_8_65 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_8_77 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_8_83 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_8_85 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_8_90 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_8_97 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_9_104 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_9_110 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_9_113 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_9_128 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_9_135 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_9_139 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_9_14 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_9_145 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_9_160 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_9_169 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_9_176 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_9_193 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_9_200 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_9_204 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_9_218 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_9_225 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_9_229 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_9_243 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_9_250 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_9_257 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_9_264 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_9_271 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_9_278 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_9_281 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_9_286 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_9_293 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_9_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_9_32 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_9_54 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_9_57 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_9_78 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_9_8 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_9_98 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_0 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_1 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_10 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_100 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_101 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_102 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_103 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_104 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_105 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_106 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_107 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_108 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_109 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_11 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_110 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_111 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_112 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_113 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_114 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_115 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_12 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_13 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_14 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_15 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_16 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_17 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_18 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_19 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_2 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_20 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_21 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_22 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_23 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_24 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_25 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_26 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_27 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_28 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_29 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_30 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_31 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_32 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_33 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_34 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_35 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_36 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_37 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_38 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_39 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_4 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_40 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_41 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_42 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_43 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_44 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_45 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_46 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_47 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_48 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_49 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_5 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_50 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_51 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_52 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_53 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_54 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_55 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_56 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_57 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_58 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_59 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_6 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_60 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_61 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_62 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_63 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_64 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_65 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_66 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_67 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_68 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_69 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_7 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_70 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_71 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_72 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_73 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_74 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_75 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_76 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_77 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_78 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_79 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_8 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_80 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_81 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_82 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_83 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_84 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_85 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_86 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_87 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_88 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_89 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_9 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_90 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_91 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_92 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_93 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_94 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_95 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_96 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_97 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_98 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_99 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_116 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_117 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_118 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_119 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_120 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_121 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_122 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_123 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_124 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_125 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_126 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_127 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_128 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_129 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_130 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_131 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_132 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_133 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_134 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_135 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_136 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_137 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_138 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_139 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_140 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_141 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_142 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_143 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_144 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_145 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_146 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_147 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_148 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_149 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_150 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_151 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_152 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_153 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_154 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_155 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_156 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_157 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_158 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_159 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_160 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_161 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_162 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_163 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_164 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_165 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_166 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_167 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_168 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_169 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_170 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_171 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_172 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_173 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_174 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_175 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_176 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_177 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_178 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_179 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_180 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_181 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_182 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_183 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_184 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_185 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_186 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_187 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_188 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_189 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_190 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_191 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_192 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_193 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_194 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_195 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_196 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_197 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_198 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_199 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_200 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_201 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_202 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_203 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_204 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_205 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_206 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_207 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_208 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_209 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_210 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_211 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_212 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_213 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_214 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_215 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_216 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_217 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_218 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_219 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_220 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_221 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_222 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_223 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_224 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_225 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_226 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_227 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_228 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_229 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_230 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_231 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_232 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_233 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_234 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_235 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_236 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_237 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_238 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_239 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_240 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_241 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_242 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_243 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_244 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_245 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_246 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_247 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_248 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_249 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_250 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_251 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_252 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_253 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_254 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_255 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_256 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_257 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_258 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_259 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_260 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_261 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_262 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_263 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_264 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_265 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_266 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_267 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_268 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_269 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_270 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_271 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_272 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_273 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_274 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_275 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_276 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_277 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_278 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_279 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_280 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_281 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_282 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_283 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_284 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_285 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_286 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_287 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_288 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_289 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_290 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_291 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_292 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_293 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_294 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_295 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_296 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_297 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_298 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_299 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_300 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_301 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_302 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_303 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_304 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_305 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_306 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_307 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_308 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_309 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_310 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_311 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_312 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_313 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_314 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_315 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_316 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_317 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_318 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_319 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_320 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_321 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_322 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_323 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_324 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_325 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_326 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_327 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_328 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_329 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_330 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_331 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_332 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_333 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_334 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_335 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_336 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_337 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_338 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_339 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_340 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_341 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_342 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_343 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_344 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_345 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_346 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_347 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_348 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_349 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_350 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_351 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_352 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_353 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_354 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_355 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_356 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_357 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_358 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_359 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_360 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_361 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_362 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_363 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_364 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_365 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_366 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_367 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_368 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_369 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_370 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_371 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_372 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_373 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_374 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_375 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_376 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_377 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_378 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_379 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_380 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_381 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_382 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_383 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_384 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_385 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_386 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_387 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_388 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_389 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_390 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_391 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_392 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_393 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_394 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_395 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_396 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_397 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_398 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_399 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_400 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_401 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_402 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_403 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_404 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_405 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_406 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_407 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_408 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_409 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_410 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_411 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_412 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_413 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_414 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_415 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_1 _252_ (.A(\l_fifo.genblk1[46].entry.empty ),
    .B(net27),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_089_));
 sky130_fd_sc_hd__clkbuf_1 _253_ (.A(_089_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.ready ));
 sky130_fd_sc_hd__or2_1 _254_ (.A(net1),
    .B(net2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_090_));
 sky130_fd_sc_hd__clkbuf_1 _255_ (.A(_090_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(reset_n_in));
 sky130_fd_sc_hd__and4b_1 _256_ (.A_N(\l_fifo.genblk1[47].entry.write_in ),
    .B(\l_fifo.genblk1[47].entry.empty ),
    .C(\l_fifo.genblk1[46].entry.empty ),
    .D(\l_fifo.genblk1[45].entry.empty ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_091_));
 sky130_fd_sc_hd__and4_1 _257_ (.A(\l_fifo.genblk1[44].entry.empty ),
    .B(\l_fifo.genblk1[43].entry.empty ),
    .C(\l_fifo.genblk1[42].entry.empty ),
    .D(_091_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_092_));
 sky130_fd_sc_hd__and4_1 _258_ (.A(\l_fifo.genblk1[41].entry.empty ),
    .B(\l_fifo.genblk1[40].entry.empty ),
    .C(\l_fifo.genblk1[39].entry.empty ),
    .D(_092_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_093_));
 sky130_fd_sc_hd__and4_1 _259_ (.A(\l_fifo.genblk1[38].entry.empty ),
    .B(\l_fifo.genblk1[37].entry.empty ),
    .C(\l_fifo.genblk1[36].entry.empty ),
    .D(_093_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_094_));
 sky130_fd_sc_hd__and4_1 _260_ (.A(\l_fifo.genblk1[35].entry.empty ),
    .B(\l_fifo.genblk1[34].entry.empty ),
    .C(\l_fifo.genblk1[33].entry.empty ),
    .D(_094_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_095_));
 sky130_fd_sc_hd__and4_1 _261_ (.A(\l_fifo.genblk1[32].entry.empty ),
    .B(\l_fifo.genblk1[31].entry.empty ),
    .C(\l_fifo.genblk1[30].entry.empty ),
    .D(_095_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_096_));
 sky130_fd_sc_hd__and4_1 _262_ (.A(\l_fifo.genblk1[29].entry.empty ),
    .B(\l_fifo.genblk1[28].entry.empty ),
    .C(\l_fifo.genblk1[27].entry.empty ),
    .D(_096_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_097_));
 sky130_fd_sc_hd__and4_1 _263_ (.A(\l_fifo.genblk1[26].entry.empty ),
    .B(\l_fifo.genblk1[25].entry.empty ),
    .C(\l_fifo.genblk1[24].entry.empty ),
    .D(_097_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_098_));
 sky130_fd_sc_hd__and4_1 _264_ (.A(\l_fifo.genblk1[23].entry.empty ),
    .B(\l_fifo.genblk1[22].entry.empty ),
    .C(\l_fifo.genblk1[21].entry.empty ),
    .D(_098_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_099_));
 sky130_fd_sc_hd__and4_1 _265_ (.A(\l_fifo.genblk1[20].entry.empty ),
    .B(\l_fifo.genblk1[19].entry.empty ),
    .C(\l_fifo.genblk1[18].entry.empty ),
    .D(_099_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_100_));
 sky130_fd_sc_hd__and4_1 _266_ (.A(\l_fifo.genblk1[17].entry.empty ),
    .B(\l_fifo.genblk1[16].entry.empty ),
    .C(\l_fifo.genblk1[15].entry.empty ),
    .D(_100_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_101_));
 sky130_fd_sc_hd__inv_2 _267_ (.A(net25),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_102_));
 sky130_fd_sc_hd__clkbuf_4 _268_ (.A(_102_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_103_));
 sky130_fd_sc_hd__a311o_1 _269_ (.A1(\l_fifo.genblk1[14].entry.empty ),
    .A2(\l_fifo.genblk1[13].entry.empty ),
    .A3(_101_),
    .B1(_103_),
    .C1(\l_fifo.genblk1[12].entry.empty ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_000_));
 sky130_fd_sc_hd__buf_2 _270_ (.A(_102_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_104_));
 sky130_fd_sc_hd__and4_1 _271_ (.A(\l_fifo.genblk1[14].entry.empty ),
    .B(\l_fifo.genblk1[13].entry.empty ),
    .C(\l_fifo.genblk1[12].entry.empty ),
    .D(_101_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_105_));
 sky130_fd_sc_hd__or3_1 _272_ (.A(\l_fifo.genblk1[11].entry.empty ),
    .B(_104_),
    .C(_105_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_106_));
 sky130_fd_sc_hd__clkbuf_1 _273_ (.A(_106_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_001_));
 sky130_fd_sc_hd__clkbuf_4 _274_ (.A(_104_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_107_));
 sky130_fd_sc_hd__a211o_1 _275_ (.A1(\l_fifo.genblk1[11].entry.empty ),
    .A2(_105_),
    .B1(_107_),
    .C1(\l_fifo.genblk1[10].entry.empty ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_002_));
 sky130_fd_sc_hd__a311o_1 _276_ (.A1(\l_fifo.genblk1[11].entry.empty ),
    .A2(\l_fifo.genblk1[10].entry.empty ),
    .A3(_105_),
    .B1(_103_),
    .C1(\l_fifo.genblk1[10].entry.next_is_empty ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_003_));
 sky130_fd_sc_hd__and4_1 _277_ (.A(\l_fifo.genblk1[11].entry.empty ),
    .B(\l_fifo.genblk1[10].entry.empty ),
    .C(\l_fifo.genblk1[10].entry.next_is_empty ),
    .D(_105_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_108_));
 sky130_fd_sc_hd__and4_1 _278_ (.A(\l_fifo.genblk1[8].entry.empty ),
    .B(\l_fifo.genblk1[7].entry.empty ),
    .C(\l_fifo.genblk1[6].entry.empty ),
    .D(_108_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_109_));
 sky130_fd_sc_hd__and4_1 _279_ (.A(\l_fifo.genblk1[5].entry.empty ),
    .B(\l_fifo.genblk1[4].entry.empty ),
    .C(\l_fifo.genblk1[3].entry.empty ),
    .D(_109_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_110_));
 sky130_fd_sc_hd__and3_1 _280_ (.A(\l_fifo.genblk1[2].entry.empty ),
    .B(\l_fifo.genblk1[1].entry.empty ),
    .C(_110_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_111_));
 sky130_fd_sc_hd__buf_2 _281_ (.A(net22),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_112_));
 sky130_fd_sc_hd__inv_2 _282_ (.A(\f_fifo.write_addr[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_113_));
 sky130_fd_sc_hd__and2_1 _283_ (.A(_113_),
    .B(\f_fifo.read_addr[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_114_));
 sky130_fd_sc_hd__nor2_1 _284_ (.A(_113_),
    .B(\f_fifo.read_addr[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_115_));
 sky130_fd_sc_hd__xnor2_1 _285_ (.A(\f_fifo.write_addr[1] ),
    .B(\f_fifo.read_addr[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_116_));
 sky130_fd_sc_hd__and4bb_1 _286_ (.A_N(_114_),
    .B_N(_115_),
    .C(\f_fifo.empty_n ),
    .D(_116_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_117_));
 sky130_fd_sc_hd__nand2_1 _287_ (.A(_112_),
    .B(_117_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_118_));
 sky130_fd_sc_hd__a21o_1 _288_ (.A1(\l_fifo.genblk1[0].entry.empty ),
    .A2(_111_),
    .B1(_118_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_004_));
 sky130_fd_sc_hd__a211o_1 _289_ (.A1(\l_fifo.genblk1[8].entry.empty ),
    .A2(_108_),
    .B1(_107_),
    .C1(\l_fifo.genblk1[7].entry.empty ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_005_));
 sky130_fd_sc_hd__a311o_1 _290_ (.A1(\l_fifo.genblk1[8].entry.empty ),
    .A2(\l_fifo.genblk1[7].entry.empty ),
    .A3(_108_),
    .B1(_103_),
    .C1(\l_fifo.genblk1[6].entry.empty ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_006_));
 sky130_fd_sc_hd__or3_1 _291_ (.A(\l_fifo.genblk1[5].entry.empty ),
    .B(_104_),
    .C(_109_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_119_));
 sky130_fd_sc_hd__clkbuf_1 _292_ (.A(_119_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_007_));
 sky130_fd_sc_hd__a211o_1 _293_ (.A1(\l_fifo.genblk1[5].entry.empty ),
    .A2(_109_),
    .B1(_107_),
    .C1(\l_fifo.genblk1[4].entry.empty ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_008_));
 sky130_fd_sc_hd__clkbuf_4 _294_ (.A(_102_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_120_));
 sky130_fd_sc_hd__a311o_1 _295_ (.A1(\l_fifo.genblk1[5].entry.empty ),
    .A2(\l_fifo.genblk1[4].entry.empty ),
    .A3(_109_),
    .B1(_120_),
    .C1(\l_fifo.genblk1[3].entry.empty ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_009_));
 sky130_fd_sc_hd__and2b_1 _296_ (.A_N(\l_fifo.genblk1[47].entry.write_in ),
    .B(\l_fifo.genblk1[47].entry.empty ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_121_));
 sky130_fd_sc_hd__or3_1 _297_ (.A(\l_fifo.genblk1[46].entry.empty ),
    .B(_104_),
    .C(_121_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_122_));
 sky130_fd_sc_hd__clkbuf_1 _298_ (.A(_122_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_010_));
 sky130_fd_sc_hd__or3_1 _299_ (.A(\l_fifo.genblk1[38].entry.empty ),
    .B(_104_),
    .C(_093_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_123_));
 sky130_fd_sc_hd__clkbuf_1 _300_ (.A(_123_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_011_));
 sky130_fd_sc_hd__a211o_1 _301_ (.A1(\l_fifo.genblk1[29].entry.empty ),
    .A2(_096_),
    .B1(_107_),
    .C1(\l_fifo.genblk1[28].entry.empty ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_012_));
 sky130_fd_sc_hd__a311o_1 _302_ (.A1(\l_fifo.genblk1[20].entry.empty ),
    .A2(\l_fifo.genblk1[19].entry.empty ),
    .A3(_099_),
    .B1(_120_),
    .C1(\l_fifo.genblk1[18].entry.empty ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_013_));
 sky130_fd_sc_hd__and2_1 _303_ (.A(net1),
    .B(net2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_124_));
 sky130_fd_sc_hd__clkbuf_1 _304_ (.A(_124_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_014_));
 sky130_fd_sc_hd__and2_1 _305_ (.A(net3),
    .B(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_125_));
 sky130_fd_sc_hd__clkbuf_1 _306_ (.A(_125_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_015_));
 sky130_fd_sc_hd__and2_1 _307_ (.A(net1),
    .B(net4),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_126_));
 sky130_fd_sc_hd__clkbuf_1 _308_ (.A(_126_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_016_));
 sky130_fd_sc_hd__and2_1 _309_ (.A(net1),
    .B(net5),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_127_));
 sky130_fd_sc_hd__clkbuf_1 _310_ (.A(_127_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_017_));
 sky130_fd_sc_hd__and2_1 _311_ (.A(net1),
    .B(net6),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_128_));
 sky130_fd_sc_hd__clkbuf_1 _312_ (.A(_128_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_018_));
 sky130_fd_sc_hd__and2_1 _313_ (.A(net1),
    .B(net7),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_129_));
 sky130_fd_sc_hd__clkbuf_1 _314_ (.A(_129_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_019_));
 sky130_fd_sc_hd__inv_2 _315_ (.A(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_130_));
 sky130_fd_sc_hd__and3_1 _316_ (.A(\f_fifo.empty_n ),
    .B(net3),
    .C(_130_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_131_));
 sky130_fd_sc_hd__and2_1 _317_ (.A(\f_fifo.read_addr[0] ),
    .B(_131_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_132_));
 sky130_fd_sc_hd__o21ai_1 _318_ (.A1(\f_fifo.read_addr[0] ),
    .A2(_131_),
    .B1(_112_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_133_));
 sky130_fd_sc_hd__nor2_1 _319_ (.A(_132_),
    .B(_133_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_020_));
 sky130_fd_sc_hd__a31o_1 _320_ (.A1(\f_fifo.read_addr[1] ),
    .A2(\f_fifo.read_addr[0] ),
    .A3(_131_),
    .B1(_104_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_134_));
 sky130_fd_sc_hd__o21ba_1 _321_ (.A1(\f_fifo.read_addr[1] ),
    .A2(_132_),
    .B1_N(_134_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_021_));
 sky130_fd_sc_hd__a41o_1 _322_ (.A1(\l_fifo.genblk1[2].entry.empty ),
    .A2(\l_fifo.genblk1[1].entry.empty ),
    .A3(\l_fifo.genblk1[0].entry.empty ),
    .A4(_110_),
    .B1(_117_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_135_));
 sky130_fd_sc_hd__clkbuf_4 _323_ (.A(_135_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_136_));
 sky130_fd_sc_hd__o21ai_1 _324_ (.A1(_113_),
    .A2(_136_),
    .B1(_112_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_137_));
 sky130_fd_sc_hd__a21oi_1 _325_ (.A1(_113_),
    .A2(_136_),
    .B1(_137_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_022_));
 sky130_fd_sc_hd__nor2_2 _326_ (.A(\f_fifo.write_addr[1] ),
    .B(\f_fifo.write_addr[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_138_));
 sky130_fd_sc_hd__and2_2 _327_ (.A(\f_fifo.write_addr[1] ),
    .B(\f_fifo.write_addr[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_139_));
 sky130_fd_sc_hd__nor2_1 _328_ (.A(_138_),
    .B(_139_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_140_));
 sky130_fd_sc_hd__mux2_1 _329_ (.A0(_140_),
    .A1(\f_fifo.write_addr[1] ),
    .S(_136_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_141_));
 sky130_fd_sc_hd__and2_1 _330_ (.A(_112_),
    .B(_141_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_142_));
 sky130_fd_sc_hd__clkbuf_1 _331_ (.A(_142_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_023_));
 sky130_fd_sc_hd__mux2_1 _332_ (.A0(_114_),
    .A1(_115_),
    .S(_116_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_143_));
 sky130_fd_sc_hd__nand2_2 _333_ (.A(_131_),
    .B(_143_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_144_));
 sky130_fd_sc_hd__nand2_1 _334_ (.A(\f_fifo.empty_n ),
    .B(_144_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_145_));
 sky130_fd_sc_hd__a21oi_1 _335_ (.A1(_136_),
    .A2(_145_),
    .B1(_107_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_024_));
 sky130_fd_sc_hd__clkbuf_2 _336_ (.A(net22),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_146_));
 sky130_fd_sc_hd__a21bo_1 _337_ (.A1(_135_),
    .A2(_144_),
    .B1_N(_138_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_147_));
 sky130_fd_sc_hd__inv_2 _338_ (.A(\f_fifo.data_in[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_148_));
 sky130_fd_sc_hd__nor2_2 _339_ (.A(_148_),
    .B(_136_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_149_));
 sky130_fd_sc_hd__a22o_1 _340_ (.A1(\f_fifo.fifo_data[0][0] ),
    .A2(_147_),
    .B1(_149_),
    .B2(_138_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_150_));
 sky130_fd_sc_hd__and2_1 _341_ (.A(_146_),
    .B(_150_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_151_));
 sky130_fd_sc_hd__clkbuf_1 _342_ (.A(_151_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_025_));
 sky130_fd_sc_hd__inv_2 _343_ (.A(\f_fifo.data_in[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_152_));
 sky130_fd_sc_hd__nor2_1 _344_ (.A(_152_),
    .B(_136_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_153_));
 sky130_fd_sc_hd__a22o_1 _345_ (.A1(\f_fifo.fifo_data[0][1] ),
    .A2(_147_),
    .B1(_153_),
    .B2(_138_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_154_));
 sky130_fd_sc_hd__and2_1 _346_ (.A(_146_),
    .B(_154_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_155_));
 sky130_fd_sc_hd__clkbuf_1 _347_ (.A(_155_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_026_));
 sky130_fd_sc_hd__inv_2 _348_ (.A(\f_fifo.data_in[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_156_));
 sky130_fd_sc_hd__nor2_2 _349_ (.A(_156_),
    .B(_136_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_157_));
 sky130_fd_sc_hd__a22o_1 _350_ (.A1(\f_fifo.fifo_data[0][2] ),
    .A2(_147_),
    .B1(_157_),
    .B2(_138_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_158_));
 sky130_fd_sc_hd__and2_1 _351_ (.A(_146_),
    .B(_158_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_159_));
 sky130_fd_sc_hd__clkbuf_1 _352_ (.A(_159_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_027_));
 sky130_fd_sc_hd__inv_2 _353_ (.A(\f_fifo.data_in[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_160_));
 sky130_fd_sc_hd__nor2_1 _354_ (.A(_160_),
    .B(_136_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_161_));
 sky130_fd_sc_hd__a22o_1 _355_ (.A1(\f_fifo.fifo_data[0][3] ),
    .A2(_147_),
    .B1(_161_),
    .B2(_138_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_162_));
 sky130_fd_sc_hd__and2_1 _356_ (.A(_146_),
    .B(_162_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_163_));
 sky130_fd_sc_hd__clkbuf_1 _357_ (.A(_163_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_028_));
 sky130_fd_sc_hd__inv_2 _358_ (.A(\f_fifo.data_in[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_164_));
 sky130_fd_sc_hd__nor2_1 _359_ (.A(_164_),
    .B(_136_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_165_));
 sky130_fd_sc_hd__a22o_1 _360_ (.A1(\f_fifo.fifo_data[0][4] ),
    .A2(_147_),
    .B1(_165_),
    .B2(_138_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_166_));
 sky130_fd_sc_hd__and2_1 _361_ (.A(_146_),
    .B(_166_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_167_));
 sky130_fd_sc_hd__clkbuf_1 _362_ (.A(_167_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_029_));
 sky130_fd_sc_hd__inv_2 _363_ (.A(\f_fifo.data_in[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_168_));
 sky130_fd_sc_hd__nor2_2 _364_ (.A(_168_),
    .B(_136_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_169_));
 sky130_fd_sc_hd__a22o_1 _365_ (.A1(\f_fifo.fifo_data[0][5] ),
    .A2(_147_),
    .B1(_169_),
    .B2(_138_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_170_));
 sky130_fd_sc_hd__and2_1 _366_ (.A(_146_),
    .B(_170_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_171_));
 sky130_fd_sc_hd__clkbuf_1 _367_ (.A(_171_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_030_));
 sky130_fd_sc_hd__nor2_2 _368_ (.A(\f_fifo.write_addr[1] ),
    .B(_113_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_172_));
 sky130_fd_sc_hd__a21bo_1 _369_ (.A1(_135_),
    .A2(_144_),
    .B1_N(_172_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_173_));
 sky130_fd_sc_hd__a22o_1 _370_ (.A1(_149_),
    .A2(_172_),
    .B1(_173_),
    .B2(\f_fifo.fifo_data[1][0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_174_));
 sky130_fd_sc_hd__and2_1 _371_ (.A(_146_),
    .B(_174_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_175_));
 sky130_fd_sc_hd__clkbuf_1 _372_ (.A(_175_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_031_));
 sky130_fd_sc_hd__a22o_1 _373_ (.A1(_153_),
    .A2(_172_),
    .B1(_173_),
    .B2(\f_fifo.fifo_data[1][1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_176_));
 sky130_fd_sc_hd__and2_1 _374_ (.A(_146_),
    .B(_176_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_177_));
 sky130_fd_sc_hd__clkbuf_1 _375_ (.A(_177_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_032_));
 sky130_fd_sc_hd__a22o_1 _376_ (.A1(_157_),
    .A2(_172_),
    .B1(_173_),
    .B2(\f_fifo.fifo_data[1][2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_178_));
 sky130_fd_sc_hd__and2_1 _377_ (.A(_146_),
    .B(_178_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_179_));
 sky130_fd_sc_hd__clkbuf_1 _378_ (.A(_179_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_033_));
 sky130_fd_sc_hd__a22o_1 _379_ (.A1(_161_),
    .A2(_172_),
    .B1(_173_),
    .B2(\f_fifo.fifo_data[1][3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_180_));
 sky130_fd_sc_hd__and2_1 _380_ (.A(_146_),
    .B(_180_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_181_));
 sky130_fd_sc_hd__clkbuf_1 _381_ (.A(_181_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_034_));
 sky130_fd_sc_hd__clkbuf_2 _382_ (.A(net10),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_182_));
 sky130_fd_sc_hd__a22o_1 _383_ (.A1(_165_),
    .A2(_172_),
    .B1(_173_),
    .B2(\f_fifo.fifo_data[1][4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_183_));
 sky130_fd_sc_hd__and2_1 _384_ (.A(_182_),
    .B(_183_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_184_));
 sky130_fd_sc_hd__clkbuf_1 _385_ (.A(_184_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_035_));
 sky130_fd_sc_hd__a22o_1 _386_ (.A1(_169_),
    .A2(_172_),
    .B1(_173_),
    .B2(\f_fifo.fifo_data[1][5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_185_));
 sky130_fd_sc_hd__and2_1 _387_ (.A(_182_),
    .B(_185_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_186_));
 sky130_fd_sc_hd__clkbuf_1 _388_ (.A(_186_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_036_));
 sky130_fd_sc_hd__and2_2 _389_ (.A(\f_fifo.write_addr[1] ),
    .B(_113_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_187_));
 sky130_fd_sc_hd__a21bo_1 _390_ (.A1(_135_),
    .A2(_144_),
    .B1_N(_187_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_188_));
 sky130_fd_sc_hd__a22o_1 _391_ (.A1(_149_),
    .A2(_187_),
    .B1(_188_),
    .B2(\f_fifo.fifo_data[2][0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_189_));
 sky130_fd_sc_hd__and2_1 _392_ (.A(_182_),
    .B(_189_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_190_));
 sky130_fd_sc_hd__clkbuf_1 _393_ (.A(_190_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_037_));
 sky130_fd_sc_hd__a22o_1 _394_ (.A1(_153_),
    .A2(_187_),
    .B1(_188_),
    .B2(\f_fifo.fifo_data[2][1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_191_));
 sky130_fd_sc_hd__and2_1 _395_ (.A(_182_),
    .B(_191_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_192_));
 sky130_fd_sc_hd__clkbuf_1 _396_ (.A(_192_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_038_));
 sky130_fd_sc_hd__a22o_1 _397_ (.A1(_157_),
    .A2(_187_),
    .B1(_188_),
    .B2(\f_fifo.fifo_data[2][2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_193_));
 sky130_fd_sc_hd__and2_1 _398_ (.A(_182_),
    .B(_193_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_194_));
 sky130_fd_sc_hd__clkbuf_1 _399_ (.A(_194_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_039_));
 sky130_fd_sc_hd__a22o_1 _400_ (.A1(_161_),
    .A2(_187_),
    .B1(_188_),
    .B2(\f_fifo.fifo_data[2][3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_195_));
 sky130_fd_sc_hd__and2_1 _401_ (.A(_182_),
    .B(_195_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_196_));
 sky130_fd_sc_hd__clkbuf_1 _402_ (.A(_196_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_040_));
 sky130_fd_sc_hd__a22o_1 _403_ (.A1(_165_),
    .A2(_187_),
    .B1(_188_),
    .B2(\f_fifo.fifo_data[2][4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_197_));
 sky130_fd_sc_hd__and2_1 _404_ (.A(_182_),
    .B(_197_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_198_));
 sky130_fd_sc_hd__clkbuf_1 _405_ (.A(_198_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_041_));
 sky130_fd_sc_hd__a22o_1 _406_ (.A1(_169_),
    .A2(_187_),
    .B1(_188_),
    .B2(\f_fifo.fifo_data[2][5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_199_));
 sky130_fd_sc_hd__and2_1 _407_ (.A(_182_),
    .B(_199_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_200_));
 sky130_fd_sc_hd__clkbuf_1 _408_ (.A(_200_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_042_));
 sky130_fd_sc_hd__a21bo_1 _409_ (.A1(_135_),
    .A2(_144_),
    .B1_N(_139_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_201_));
 sky130_fd_sc_hd__a22o_1 _410_ (.A1(_139_),
    .A2(_149_),
    .B1(_201_),
    .B2(\f_fifo.fifo_data[3][0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_202_));
 sky130_fd_sc_hd__and2_1 _411_ (.A(_182_),
    .B(_202_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_203_));
 sky130_fd_sc_hd__clkbuf_1 _412_ (.A(_203_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_043_));
 sky130_fd_sc_hd__a22o_1 _413_ (.A1(_139_),
    .A2(_153_),
    .B1(_201_),
    .B2(\f_fifo.fifo_data[3][1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_204_));
 sky130_fd_sc_hd__and2_1 _414_ (.A(_182_),
    .B(_204_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_205_));
 sky130_fd_sc_hd__clkbuf_1 _415_ (.A(_205_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_044_));
 sky130_fd_sc_hd__a22o_1 _416_ (.A1(_139_),
    .A2(_157_),
    .B1(_201_),
    .B2(\f_fifo.fifo_data[3][2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_206_));
 sky130_fd_sc_hd__and2_1 _417_ (.A(net22),
    .B(_206_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_207_));
 sky130_fd_sc_hd__clkbuf_1 _418_ (.A(_207_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_045_));
 sky130_fd_sc_hd__a22o_1 _419_ (.A1(_139_),
    .A2(_161_),
    .B1(_201_),
    .B2(\f_fifo.fifo_data[3][3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_208_));
 sky130_fd_sc_hd__and2_1 _420_ (.A(net22),
    .B(_208_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_209_));
 sky130_fd_sc_hd__clkbuf_1 _421_ (.A(_209_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_046_));
 sky130_fd_sc_hd__a22o_1 _422_ (.A1(_139_),
    .A2(_165_),
    .B1(_201_),
    .B2(\f_fifo.fifo_data[3][4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_210_));
 sky130_fd_sc_hd__and2_1 _423_ (.A(net9),
    .B(_210_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_211_));
 sky130_fd_sc_hd__clkbuf_1 _424_ (.A(_211_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_047_));
 sky130_fd_sc_hd__a22o_1 _425_ (.A1(_139_),
    .A2(_169_),
    .B1(_201_),
    .B2(\f_fifo.fifo_data[3][5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_212_));
 sky130_fd_sc_hd__and2_1 _426_ (.A(net22),
    .B(_212_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_213_));
 sky130_fd_sc_hd__clkbuf_1 _427_ (.A(_213_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_048_));
 sky130_fd_sc_hd__and2_1 _428_ (.A(_130_),
    .B(net5),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_214_));
 sky130_fd_sc_hd__xnor2_2 _429_ (.A(\f_fifo.read_addr[1] ),
    .B(_214_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_215_));
 sky130_fd_sc_hd__inv_2 _430_ (.A(_215_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_216_));
 sky130_fd_sc_hd__a21oi_1 _431_ (.A1(_130_),
    .A2(net4),
    .B1(\f_fifo.read_addr[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_217_));
 sky130_fd_sc_hd__and3_1 _432_ (.A(\f_fifo.read_addr[0] ),
    .B(_130_),
    .C(net4),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_218_));
 sky130_fd_sc_hd__or2_1 _433_ (.A(_215_),
    .B(_218_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_219_));
 sky130_fd_sc_hd__o21ai_2 _434_ (.A1(_216_),
    .A2(_217_),
    .B1(_219_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_220_));
 sky130_fd_sc_hd__or2_1 _435_ (.A(_217_),
    .B(_218_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_221_));
 sky130_fd_sc_hd__buf_2 _436_ (.A(_221_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_222_));
 sky130_fd_sc_hd__o21a_1 _437_ (.A1(_216_),
    .A2(_217_),
    .B1(_219_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_223_));
 sky130_fd_sc_hd__a21o_1 _438_ (.A1(\f_fifo.fifo_data[2][0] ),
    .A2(_222_),
    .B1(_223_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_224_));
 sky130_fd_sc_hd__nor2_2 _439_ (.A(_215_),
    .B(_222_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_225_));
 sky130_fd_sc_hd__nor2_2 _440_ (.A(_216_),
    .B(_222_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_226_));
 sky130_fd_sc_hd__a22o_1 _441_ (.A1(\f_fifo.fifo_data[3][0] ),
    .A2(_225_),
    .B1(_226_),
    .B2(\f_fifo.fifo_data[1][0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_227_));
 sky130_fd_sc_hd__o221a_1 _442_ (.A1(\f_fifo.fifo_data[0][0] ),
    .A2(_220_),
    .B1(_224_),
    .B2(_227_),
    .C1(_112_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_049_));
 sky130_fd_sc_hd__a22o_1 _443_ (.A1(\f_fifo.fifo_data[3][1] ),
    .A2(_225_),
    .B1(_226_),
    .B2(\f_fifo.fifo_data[1][1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_228_));
 sky130_fd_sc_hd__a21o_1 _444_ (.A1(\f_fifo.fifo_data[2][1] ),
    .A2(_222_),
    .B1(_223_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_229_));
 sky130_fd_sc_hd__o221a_1 _445_ (.A1(\f_fifo.fifo_data[0][1] ),
    .A2(_220_),
    .B1(_228_),
    .B2(_229_),
    .C1(_112_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_050_));
 sky130_fd_sc_hd__a22o_1 _446_ (.A1(\f_fifo.fifo_data[3][2] ),
    .A2(_225_),
    .B1(_226_),
    .B2(\f_fifo.fifo_data[1][2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_230_));
 sky130_fd_sc_hd__a21o_1 _447_ (.A1(\f_fifo.fifo_data[2][2] ),
    .A2(_222_),
    .B1(_223_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_231_));
 sky130_fd_sc_hd__o221a_1 _448_ (.A1(\f_fifo.fifo_data[0][2] ),
    .A2(_220_),
    .B1(_230_),
    .B2(_231_),
    .C1(_112_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_051_));
 sky130_fd_sc_hd__a22o_1 _449_ (.A1(\f_fifo.fifo_data[3][3] ),
    .A2(_225_),
    .B1(_226_),
    .B2(\f_fifo.fifo_data[1][3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_232_));
 sky130_fd_sc_hd__a21o_1 _450_ (.A1(\f_fifo.fifo_data[2][3] ),
    .A2(_222_),
    .B1(_223_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_233_));
 sky130_fd_sc_hd__o221a_1 _451_ (.A1(\f_fifo.fifo_data[0][3] ),
    .A2(_220_),
    .B1(_232_),
    .B2(_233_),
    .C1(_112_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_052_));
 sky130_fd_sc_hd__a22o_1 _452_ (.A1(\f_fifo.fifo_data[3][4] ),
    .A2(_225_),
    .B1(_226_),
    .B2(\f_fifo.fifo_data[1][4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_234_));
 sky130_fd_sc_hd__a21o_1 _453_ (.A1(\f_fifo.fifo_data[2][4] ),
    .A2(_222_),
    .B1(_223_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_235_));
 sky130_fd_sc_hd__o221a_1 _454_ (.A1(\f_fifo.fifo_data[0][4] ),
    .A2(_220_),
    .B1(_234_),
    .B2(_235_),
    .C1(_112_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_053_));
 sky130_fd_sc_hd__a221o_1 _455_ (.A1(\f_fifo.fifo_data[2][5] ),
    .A2(_222_),
    .B1(_225_),
    .B2(\f_fifo.fifo_data[3][5] ),
    .C1(_223_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_236_));
 sky130_fd_sc_hd__a21o_1 _456_ (.A1(\f_fifo.fifo_data[1][5] ),
    .A2(_226_),
    .B1(_236_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_237_));
 sky130_fd_sc_hd__o211a_1 _457_ (.A1(\f_fifo.fifo_data[0][5] ),
    .A2(_220_),
    .B1(_237_),
    .C1(_112_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_054_));
 sky130_fd_sc_hd__or3_1 _458_ (.A(\l_fifo.genblk1[8].entry.empty ),
    .B(_104_),
    .C(_108_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_238_));
 sky130_fd_sc_hd__clkbuf_1 _459_ (.A(_238_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_055_));
 sky130_fd_sc_hd__a211o_1 _460_ (.A1(\l_fifo.genblk1[46].entry.empty ),
    .A2(_121_),
    .B1(_107_),
    .C1(\l_fifo.genblk1[45].entry.empty ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_056_));
 sky130_fd_sc_hd__or3_1 _461_ (.A(\l_fifo.genblk1[44].entry.empty ),
    .B(_104_),
    .C(_091_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_239_));
 sky130_fd_sc_hd__clkbuf_1 _462_ (.A(_239_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_057_));
 sky130_fd_sc_hd__a211o_1 _463_ (.A1(\l_fifo.genblk1[44].entry.empty ),
    .A2(_091_),
    .B1(_107_),
    .C1(\l_fifo.genblk1[43].entry.empty ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_058_));
 sky130_fd_sc_hd__a311o_1 _464_ (.A1(\l_fifo.genblk1[44].entry.empty ),
    .A2(\l_fifo.genblk1[43].entry.empty ),
    .A3(_091_),
    .B1(_120_),
    .C1(\l_fifo.genblk1[42].entry.empty ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_059_));
 sky130_fd_sc_hd__or3_1 _465_ (.A(\l_fifo.genblk1[41].entry.empty ),
    .B(_104_),
    .C(_092_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_240_));
 sky130_fd_sc_hd__clkbuf_1 _466_ (.A(_240_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_060_));
 sky130_fd_sc_hd__a211o_1 _467_ (.A1(\l_fifo.genblk1[41].entry.empty ),
    .A2(_092_),
    .B1(_107_),
    .C1(\l_fifo.genblk1[40].entry.empty ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_061_));
 sky130_fd_sc_hd__a311o_1 _468_ (.A1(\l_fifo.genblk1[41].entry.empty ),
    .A2(\l_fifo.genblk1[40].entry.empty ),
    .A3(_092_),
    .B1(_120_),
    .C1(\l_fifo.genblk1[39].entry.empty ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_062_));
 sky130_fd_sc_hd__clkbuf_4 _469_ (.A(_102_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_241_));
 sky130_fd_sc_hd__or3_1 _470_ (.A(\l_fifo.genblk1[2].entry.empty ),
    .B(_241_),
    .C(_110_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_242_));
 sky130_fd_sc_hd__clkbuf_1 _471_ (.A(_242_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_063_));
 sky130_fd_sc_hd__a211o_1 _472_ (.A1(\l_fifo.genblk1[38].entry.empty ),
    .A2(_093_),
    .B1(_107_),
    .C1(\l_fifo.genblk1[37].entry.empty ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_064_));
 sky130_fd_sc_hd__a311o_1 _473_ (.A1(\l_fifo.genblk1[38].entry.empty ),
    .A2(\l_fifo.genblk1[37].entry.empty ),
    .A3(_093_),
    .B1(_120_),
    .C1(\l_fifo.genblk1[36].entry.empty ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_065_));
 sky130_fd_sc_hd__or3_1 _474_ (.A(\l_fifo.genblk1[35].entry.empty ),
    .B(_241_),
    .C(_094_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_243_));
 sky130_fd_sc_hd__clkbuf_1 _475_ (.A(_243_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_066_));
 sky130_fd_sc_hd__a211o_1 _476_ (.A1(\l_fifo.genblk1[35].entry.empty ),
    .A2(_094_),
    .B1(_107_),
    .C1(\l_fifo.genblk1[34].entry.empty ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_067_));
 sky130_fd_sc_hd__a311o_1 _477_ (.A1(\l_fifo.genblk1[35].entry.empty ),
    .A2(\l_fifo.genblk1[34].entry.empty ),
    .A3(_094_),
    .B1(_120_),
    .C1(\l_fifo.genblk1[33].entry.empty ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_068_));
 sky130_fd_sc_hd__or3_1 _478_ (.A(\l_fifo.genblk1[32].entry.empty ),
    .B(_241_),
    .C(_095_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_244_));
 sky130_fd_sc_hd__clkbuf_1 _479_ (.A(_244_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_069_));
 sky130_fd_sc_hd__a211o_1 _480_ (.A1(\l_fifo.genblk1[32].entry.empty ),
    .A2(_095_),
    .B1(_103_),
    .C1(\l_fifo.genblk1[31].entry.empty ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_070_));
 sky130_fd_sc_hd__a311o_1 _481_ (.A1(\l_fifo.genblk1[32].entry.empty ),
    .A2(\l_fifo.genblk1[31].entry.empty ),
    .A3(_095_),
    .B1(_120_),
    .C1(\l_fifo.genblk1[30].entry.empty ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_071_));
 sky130_fd_sc_hd__or3_1 _482_ (.A(\l_fifo.genblk1[29].entry.empty ),
    .B(_241_),
    .C(_096_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_245_));
 sky130_fd_sc_hd__clkbuf_1 _483_ (.A(_245_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_072_));
 sky130_fd_sc_hd__a211o_1 _484_ (.A1(\l_fifo.genblk1[2].entry.empty ),
    .A2(_110_),
    .B1(_103_),
    .C1(\l_fifo.genblk1[1].entry.empty ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_073_));
 sky130_fd_sc_hd__a311o_1 _485_ (.A1(\l_fifo.genblk1[29].entry.empty ),
    .A2(\l_fifo.genblk1[28].entry.empty ),
    .A3(_096_),
    .B1(_120_),
    .C1(\l_fifo.genblk1[27].entry.empty ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_074_));
 sky130_fd_sc_hd__or3_1 _486_ (.A(\l_fifo.genblk1[26].entry.empty ),
    .B(_241_),
    .C(_097_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_246_));
 sky130_fd_sc_hd__clkbuf_1 _487_ (.A(_246_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_075_));
 sky130_fd_sc_hd__a211o_1 _488_ (.A1(\l_fifo.genblk1[26].entry.empty ),
    .A2(_097_),
    .B1(_103_),
    .C1(\l_fifo.genblk1[25].entry.empty ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_076_));
 sky130_fd_sc_hd__a311o_1 _489_ (.A1(\l_fifo.genblk1[26].entry.empty ),
    .A2(\l_fifo.genblk1[25].entry.empty ),
    .A3(_097_),
    .B1(_120_),
    .C1(\l_fifo.genblk1[24].entry.empty ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_077_));
 sky130_fd_sc_hd__or3_1 _490_ (.A(\l_fifo.genblk1[23].entry.empty ),
    .B(_241_),
    .C(_098_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_247_));
 sky130_fd_sc_hd__clkbuf_1 _491_ (.A(_247_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_078_));
 sky130_fd_sc_hd__a211o_1 _492_ (.A1(\l_fifo.genblk1[23].entry.empty ),
    .A2(_098_),
    .B1(_103_),
    .C1(\l_fifo.genblk1[22].entry.empty ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_079_));
 sky130_fd_sc_hd__a311o_1 _493_ (.A1(\l_fifo.genblk1[23].entry.empty ),
    .A2(\l_fifo.genblk1[22].entry.empty ),
    .A3(_098_),
    .B1(_120_),
    .C1(\l_fifo.genblk1[21].entry.empty ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_080_));
 sky130_fd_sc_hd__or3_1 _494_ (.A(\l_fifo.genblk1[20].entry.empty ),
    .B(_241_),
    .C(_099_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_248_));
 sky130_fd_sc_hd__clkbuf_1 _495_ (.A(_248_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_081_));
 sky130_fd_sc_hd__a211o_1 _496_ (.A1(\l_fifo.genblk1[20].entry.empty ),
    .A2(_099_),
    .B1(_103_),
    .C1(\l_fifo.genblk1[19].entry.empty ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_082_));
 sky130_fd_sc_hd__or3_1 _497_ (.A(\l_fifo.genblk1[0].entry.empty ),
    .B(_241_),
    .C(_111_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_249_));
 sky130_fd_sc_hd__clkbuf_1 _498_ (.A(_249_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_083_));
 sky130_fd_sc_hd__or3_1 _499_ (.A(\l_fifo.genblk1[17].entry.empty ),
    .B(_241_),
    .C(_100_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_250_));
 sky130_fd_sc_hd__clkbuf_1 _500_ (.A(_250_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_084_));
 sky130_fd_sc_hd__a211o_1 _501_ (.A1(\l_fifo.genblk1[17].entry.empty ),
    .A2(_100_),
    .B1(_103_),
    .C1(\l_fifo.genblk1[16].entry.empty ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_085_));
 sky130_fd_sc_hd__a311o_1 _502_ (.A1(\l_fifo.genblk1[17].entry.empty ),
    .A2(\l_fifo.genblk1[16].entry.empty ),
    .A3(_100_),
    .B1(_104_),
    .C1(\l_fifo.genblk1[15].entry.empty ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_086_));
 sky130_fd_sc_hd__or3_1 _503_ (.A(\l_fifo.genblk1[14].entry.empty ),
    .B(_241_),
    .C(_101_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_251_));
 sky130_fd_sc_hd__clkbuf_1 _504_ (.A(_251_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_087_));
 sky130_fd_sc_hd__a211o_1 _505_ (.A1(\l_fifo.genblk1[14].entry.empty ),
    .A2(_101_),
    .B1(_103_),
    .C1(\l_fifo.genblk1[13].entry.empty ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_088_));
 sky130_fd_sc_hd__dfxtp_2 _506_ (.CLK(clknet_3_2__leaf_io_in[0]),
    .D(_000_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[13].entry.empty ));
 sky130_fd_sc_hd__dfxtp_2 _507_ (.CLK(clknet_3_7__leaf_io_in[0]),
    .D(_001_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[12].entry.empty ));
 sky130_fd_sc_hd__dfxtp_2 _508_ (.CLK(clknet_3_0__leaf_io_in[0]),
    .D(_002_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[11].entry.empty ));
 sky130_fd_sc_hd__dfxtp_2 _509_ (.CLK(clknet_3_7__leaf_io_in[0]),
    .D(_003_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[10].entry.empty ));
 sky130_fd_sc_hd__dfxtp_2 _510_ (.CLK(clknet_3_4__leaf_io_in[0]),
    .D(_004_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[0].entry.empty ));
 sky130_fd_sc_hd__dfxtp_2 _511_ (.CLK(clknet_3_0__leaf_io_in[0]),
    .D(_005_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[8].entry.empty ));
 sky130_fd_sc_hd__dfxtp_2 _512_ (.CLK(clknet_3_7__leaf_io_in[0]),
    .D(_006_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[7].entry.empty ));
 sky130_fd_sc_hd__dfxtp_2 _513_ (.CLK(clknet_3_5__leaf_io_in[0]),
    .D(_007_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[6].entry.empty ));
 sky130_fd_sc_hd__dfxtp_2 _514_ (.CLK(clknet_3_2__leaf_io_in[0]),
    .D(_008_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[5].entry.empty ));
 sky130_fd_sc_hd__dfxtp_2 _515_ (.CLK(clknet_3_5__leaf_io_in[0]),
    .D(_009_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[4].entry.empty ));
 sky130_fd_sc_hd__dfxtp_2 _516_ (.CLK(clknet_3_5__leaf_io_in[0]),
    .D(_010_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[47].entry.empty ));
 sky130_fd_sc_hd__dfxtp_2 _517_ (.CLK(clknet_3_1__leaf_io_in[0]),
    .D(_011_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[39].entry.empty ));
 sky130_fd_sc_hd__dfxtp_2 _518_ (.CLK(clknet_3_3__leaf_io_in[0]),
    .D(_012_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[29].entry.empty ));
 sky130_fd_sc_hd__dfxtp_2 _519_ (.CLK(clknet_3_5__leaf_io_in[0]),
    .D(_013_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[19].entry.empty ));
 sky130_fd_sc_hd__dfxtp_1 _520_ (.CLK(clknet_3_0__leaf_io_in[0]),
    .D(_014_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\data_in_buffer[0].A ));
 sky130_fd_sc_hd__dfxtp_1 _521_ (.CLK(clknet_3_1__leaf_io_in[0]),
    .D(_015_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\data_in_buffer[1].A ));
 sky130_fd_sc_hd__dfxtp_1 _522_ (.CLK(clknet_3_4__leaf_io_in[0]),
    .D(_016_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\data_in_buffer[2].A ));
 sky130_fd_sc_hd__dfxtp_1 _523_ (.CLK(clknet_3_7__leaf_io_in[0]),
    .D(_017_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\data_in_buffer[3].A ));
 sky130_fd_sc_hd__dfxtp_1 _524_ (.CLK(clknet_3_3__leaf_io_in[0]),
    .D(_018_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\data_in_buffer[4].A ));
 sky130_fd_sc_hd__dfxtp_1 _525_ (.CLK(clknet_3_1__leaf_io_in[0]),
    .D(_019_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\data_in_buffer[5].A ));
 sky130_fd_sc_hd__dfxtp_1 _526_ (.CLK(clknet_3_2__leaf_io_in[0]),
    .D(_020_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\f_fifo.read_addr[0] ));
 sky130_fd_sc_hd__dfxtp_2 _527_ (.CLK(clknet_3_5__leaf_io_in[0]),
    .D(_021_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\f_fifo.read_addr[1] ));
 sky130_fd_sc_hd__dfxtp_1 _528_ (.CLK(clknet_3_2__leaf_io_in[0]),
    .D(_022_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\f_fifo.write_addr[0] ));
 sky130_fd_sc_hd__dfxtp_2 _529_ (.CLK(clknet_3_3__leaf_io_in[0]),
    .D(_023_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\f_fifo.write_addr[1] ));
 sky130_fd_sc_hd__dfxtp_1 _530_ (.CLK(clknet_3_4__leaf_io_in[0]),
    .D(_024_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\f_fifo.empty_n ));
 sky130_fd_sc_hd__dfxtp_1 _531_ (.CLK(clknet_3_3__leaf_io_in[0]),
    .D(_025_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\f_fifo.fifo_data[0][0] ));
 sky130_fd_sc_hd__dfxtp_1 _532_ (.CLK(clknet_3_2__leaf_io_in[0]),
    .D(_026_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\f_fifo.fifo_data[0][1] ));
 sky130_fd_sc_hd__dfxtp_1 _533_ (.CLK(clknet_3_2__leaf_io_in[0]),
    .D(_027_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\f_fifo.fifo_data[0][2] ));
 sky130_fd_sc_hd__dfxtp_1 _534_ (.CLK(clknet_3_4__leaf_io_in[0]),
    .D(_028_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\f_fifo.fifo_data[0][3] ));
 sky130_fd_sc_hd__dfxtp_1 _535_ (.CLK(clknet_3_1__leaf_io_in[0]),
    .D(_029_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\f_fifo.fifo_data[0][4] ));
 sky130_fd_sc_hd__dfxtp_1 _536_ (.CLK(clknet_3_3__leaf_io_in[0]),
    .D(_030_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\f_fifo.fifo_data[0][5] ));
 sky130_fd_sc_hd__dfxtp_1 _537_ (.CLK(clknet_3_2__leaf_io_in[0]),
    .D(_031_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\f_fifo.fifo_data[1][0] ));
 sky130_fd_sc_hd__dfxtp_1 _538_ (.CLK(clknet_3_0__leaf_io_in[0]),
    .D(_032_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\f_fifo.fifo_data[1][1] ));
 sky130_fd_sc_hd__dfxtp_1 _539_ (.CLK(clknet_3_0__leaf_io_in[0]),
    .D(_033_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\f_fifo.fifo_data[1][2] ));
 sky130_fd_sc_hd__dfxtp_1 _540_ (.CLK(clknet_3_6__leaf_io_in[0]),
    .D(_034_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\f_fifo.fifo_data[1][3] ));
 sky130_fd_sc_hd__dfxtp_1 _541_ (.CLK(clknet_3_5__leaf_io_in[0]),
    .D(_035_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\f_fifo.fifo_data[1][4] ));
 sky130_fd_sc_hd__dfxtp_1 _542_ (.CLK(clknet_3_3__leaf_io_in[0]),
    .D(_036_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\f_fifo.fifo_data[1][5] ));
 sky130_fd_sc_hd__dfxtp_1 _543_ (.CLK(clknet_3_0__leaf_io_in[0]),
    .D(_037_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\f_fifo.fifo_data[2][0] ));
 sky130_fd_sc_hd__dfxtp_1 _544_ (.CLK(clknet_3_2__leaf_io_in[0]),
    .D(_038_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\f_fifo.fifo_data[2][1] ));
 sky130_fd_sc_hd__dfxtp_1 _545_ (.CLK(clknet_3_0__leaf_io_in[0]),
    .D(_039_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\f_fifo.fifo_data[2][2] ));
 sky130_fd_sc_hd__dfxtp_1 _546_ (.CLK(clknet_3_7__leaf_io_in[0]),
    .D(_040_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\f_fifo.fifo_data[2][3] ));
 sky130_fd_sc_hd__dfxtp_1 _547_ (.CLK(clknet_3_5__leaf_io_in[0]),
    .D(_041_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\f_fifo.fifo_data[2][4] ));
 sky130_fd_sc_hd__dfxtp_1 _548_ (.CLK(clknet_3_4__leaf_io_in[0]),
    .D(_042_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\f_fifo.fifo_data[2][5] ));
 sky130_fd_sc_hd__dfxtp_1 _549_ (.CLK(clknet_3_6__leaf_io_in[0]),
    .D(_043_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\f_fifo.fifo_data[3][0] ));
 sky130_fd_sc_hd__dfxtp_1 _550_ (.CLK(clknet_3_6__leaf_io_in[0]),
    .D(_044_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\f_fifo.fifo_data[3][1] ));
 sky130_fd_sc_hd__dfxtp_1 _551_ (.CLK(clknet_3_0__leaf_io_in[0]),
    .D(_045_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\f_fifo.fifo_data[3][2] ));
 sky130_fd_sc_hd__dfxtp_1 _552_ (.CLK(clknet_3_4__leaf_io_in[0]),
    .D(_046_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\f_fifo.fifo_data[3][3] ));
 sky130_fd_sc_hd__dfxtp_1 _553_ (.CLK(clknet_3_3__leaf_io_in[0]),
    .D(_047_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\f_fifo.fifo_data[3][4] ));
 sky130_fd_sc_hd__dfxtp_1 _554_ (.CLK(clknet_3_6__leaf_io_in[0]),
    .D(_048_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\f_fifo.fifo_data[3][5] ));
 sky130_fd_sc_hd__dfxtp_1 _555_ (.CLK(clknet_3_5__leaf_io_in[0]),
    .D(reset_n_in),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\f_fifo.reset_n ));
 sky130_fd_sc_hd__dfxtp_1 _556_ (.CLK(clknet_3_4__leaf_io_in[0]),
    .D(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[47].entry.write_in ));
 sky130_fd_sc_hd__dfxtp_2 _557_ (.CLK(clknet_3_3__leaf_io_in[0]),
    .D(_049_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(io_out[2]));
 sky130_fd_sc_hd__dfxtp_2 _558_ (.CLK(clknet_3_1__leaf_io_in[0]),
    .D(_050_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(io_out[3]));
 sky130_fd_sc_hd__dfxtp_2 _559_ (.CLK(clknet_3_5__leaf_io_in[0]),
    .D(_051_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(io_out[4]));
 sky130_fd_sc_hd__dfxtp_2 _560_ (.CLK(clknet_3_7__leaf_io_in[0]),
    .D(_052_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(io_out[5]));
 sky130_fd_sc_hd__dfxtp_2 _561_ (.CLK(clknet_3_3__leaf_io_in[0]),
    .D(_053_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(io_out[6]));
 sky130_fd_sc_hd__dfxtp_2 _562_ (.CLK(clknet_3_1__leaf_io_in[0]),
    .D(_054_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(io_out[7]));
 sky130_fd_sc_hd__dfxtp_2 _563_ (.CLK(clknet_3_3__leaf_io_in[0]),
    .D(_055_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[10].entry.next_is_empty ));
 sky130_fd_sc_hd__dfxtp_2 _564_ (.CLK(clknet_3_4__leaf_io_in[0]),
    .D(_056_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[46].entry.empty ));
 sky130_fd_sc_hd__dfxtp_2 _565_ (.CLK(clknet_3_3__leaf_io_in[0]),
    .D(_057_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[45].entry.empty ));
 sky130_fd_sc_hd__dfxtp_2 _566_ (.CLK(clknet_3_3__leaf_io_in[0]),
    .D(_058_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[44].entry.empty ));
 sky130_fd_sc_hd__dfxtp_2 _567_ (.CLK(clknet_3_0__leaf_io_in[0]),
    .D(_059_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[43].entry.empty ));
 sky130_fd_sc_hd__dfxtp_2 _568_ (.CLK(clknet_3_0__leaf_io_in[0]),
    .D(_060_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[42].entry.empty ));
 sky130_fd_sc_hd__dfxtp_2 _569_ (.CLK(clknet_3_0__leaf_io_in[0]),
    .D(_061_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[41].entry.empty ));
 sky130_fd_sc_hd__dfxtp_2 _570_ (.CLK(clknet_3_1__leaf_io_in[0]),
    .D(_062_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[40].entry.empty ));
 sky130_fd_sc_hd__dfxtp_2 _571_ (.CLK(clknet_3_7__leaf_io_in[0]),
    .D(_063_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[3].entry.empty ));
 sky130_fd_sc_hd__dfxtp_2 _572_ (.CLK(clknet_3_2__leaf_io_in[0]),
    .D(_064_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[38].entry.empty ));
 sky130_fd_sc_hd__dfxtp_2 _573_ (.CLK(clknet_3_0__leaf_io_in[0]),
    .D(_065_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[37].entry.empty ));
 sky130_fd_sc_hd__dfxtp_2 _574_ (.CLK(clknet_3_1__leaf_io_in[0]),
    .D(_066_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[36].entry.empty ));
 sky130_fd_sc_hd__dfxtp_2 _575_ (.CLK(clknet_3_2__leaf_io_in[0]),
    .D(_067_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[35].entry.empty ));
 sky130_fd_sc_hd__dfxtp_2 _576_ (.CLK(clknet_3_4__leaf_io_in[0]),
    .D(_068_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[34].entry.empty ));
 sky130_fd_sc_hd__dfxtp_2 _577_ (.CLK(clknet_3_2__leaf_io_in[0]),
    .D(_069_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[33].entry.empty ));
 sky130_fd_sc_hd__dfxtp_2 _578_ (.CLK(clknet_3_6__leaf_io_in[0]),
    .D(_070_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[32].entry.empty ));
 sky130_fd_sc_hd__dfxtp_2 _579_ (.CLK(clknet_3_2__leaf_io_in[0]),
    .D(_071_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[31].entry.empty ));
 sky130_fd_sc_hd__dfxtp_2 _580_ (.CLK(clknet_3_2__leaf_io_in[0]),
    .D(_072_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[30].entry.empty ));
 sky130_fd_sc_hd__dfxtp_2 _581_ (.CLK(clknet_3_5__leaf_io_in[0]),
    .D(_073_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[2].entry.empty ));
 sky130_fd_sc_hd__dfxtp_2 _582_ (.CLK(clknet_3_6__leaf_io_in[0]),
    .D(_074_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[28].entry.empty ));
 sky130_fd_sc_hd__dfxtp_2 _583_ (.CLK(clknet_3_3__leaf_io_in[0]),
    .D(_075_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[27].entry.empty ));
 sky130_fd_sc_hd__dfxtp_2 _584_ (.CLK(clknet_3_6__leaf_io_in[0]),
    .D(_076_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[26].entry.empty ));
 sky130_fd_sc_hd__dfxtp_2 _585_ (.CLK(clknet_3_2__leaf_io_in[0]),
    .D(_077_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[25].entry.empty ));
 sky130_fd_sc_hd__dfxtp_2 _586_ (.CLK(clknet_3_0__leaf_io_in[0]),
    .D(_078_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[24].entry.empty ));
 sky130_fd_sc_hd__dfxtp_2 _587_ (.CLK(clknet_3_1__leaf_io_in[0]),
    .D(_079_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[23].entry.empty ));
 sky130_fd_sc_hd__dfxtp_2 _588_ (.CLK(clknet_3_1__leaf_io_in[0]),
    .D(_080_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[22].entry.empty ));
 sky130_fd_sc_hd__dfxtp_2 _589_ (.CLK(clknet_3_0__leaf_io_in[0]),
    .D(_081_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[21].entry.empty ));
 sky130_fd_sc_hd__dfxtp_4 _590_ (.CLK(clknet_3_0__leaf_io_in[0]),
    .D(_082_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[20].entry.empty ));
 sky130_fd_sc_hd__dfxtp_2 _591_ (.CLK(clknet_3_0__leaf_io_in[0]),
    .D(_083_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[1].entry.empty ));
 sky130_fd_sc_hd__dfxtp_2 _592_ (.CLK(clknet_3_2__leaf_io_in[0]),
    .D(_084_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[18].entry.empty ));
 sky130_fd_sc_hd__dfxtp_2 _593_ (.CLK(clknet_3_7__leaf_io_in[0]),
    .D(_085_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[17].entry.empty ));
 sky130_fd_sc_hd__dfxtp_4 _594_ (.CLK(clknet_3_0__leaf_io_in[0]),
    .D(_086_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[16].entry.empty ));
 sky130_fd_sc_hd__dfxtp_2 _595_ (.CLK(clknet_3_7__leaf_io_in[0]),
    .D(_087_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[15].entry.empty ));
 sky130_fd_sc_hd__dfxtp_2 _596_ (.CLK(clknet_3_5__leaf_io_in[0]),
    .D(_088_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[14].entry.empty ));
 sky130_fd_sc_hd__buf_2 _597_ (.A(\l_fifo.ready ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(io_out[0]));
 sky130_fd_sc_hd__buf_2 _598_ (.A(\f_fifo.empty_n ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(io_out[1]));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_io_in[0]  (.A(io_in[0]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(clknet_0_io_in[0]));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_3_0__f_io_in[0]  (.A(clknet_0_io_in[0]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(clknet_3_0__leaf_io_in[0]));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_3_1__f_io_in[0]  (.A(clknet_0_io_in[0]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(clknet_3_1__leaf_io_in[0]));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_3_2__f_io_in[0]  (.A(clknet_0_io_in[0]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(clknet_3_2__leaf_io_in[0]));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_3_3__f_io_in[0]  (.A(clknet_0_io_in[0]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(clknet_3_3__leaf_io_in[0]));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_3_4__f_io_in[0]  (.A(clknet_0_io_in[0]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(clknet_3_4__leaf_io_in[0]));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_3_5__f_io_in[0]  (.A(clknet_0_io_in[0]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(clknet_3_5__leaf_io_in[0]));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_3_6__f_io_in[0]  (.A(clknet_0_io_in[0]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(clknet_3_6__leaf_io_in[0]));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_3_7__f_io_in[0]  (.A(clknet_0_io_in[0]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(clknet_3_7__leaf_io_in[0]));
 sky130_fd_sc_hd__inv_1 \data_in_buffer[0].genblk1[0].genblk1.inv_first  (.A(\data_in_buffer[0].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\data_in_buffer[0].genblk1[0].mid ));
 sky130_fd_sc_hd__inv_1 \data_in_buffer[0].genblk1[0].genblk2.inv2  (.A(\data_in_buffer[0].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\data_in_buffer[0].b[0] ));
 sky130_fd_sc_hd__inv_1 \data_in_buffer[0].genblk1[1].genblk1.inv1  (.A(\data_in_buffer[0].b[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\data_in_buffer[0].genblk1[1].mid ));
 sky130_fd_sc_hd__inv_2 \data_in_buffer[0].genblk1[1].genblk2.inv_last  (.A(\data_in_buffer[0].genblk1[1].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\data_in_buffer[0].X ));
 sky130_fd_sc_hd__inv_1 \data_in_buffer[1].genblk1[0].genblk1.inv_first  (.A(\data_in_buffer[1].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\data_in_buffer[1].genblk1[0].mid ));
 sky130_fd_sc_hd__inv_1 \data_in_buffer[1].genblk1[0].genblk2.inv2  (.A(\data_in_buffer[1].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\data_in_buffer[1].b[0] ));
 sky130_fd_sc_hd__inv_1 \data_in_buffer[1].genblk1[1].genblk1.inv1  (.A(\data_in_buffer[1].b[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\data_in_buffer[1].genblk1[1].mid ));
 sky130_fd_sc_hd__inv_2 \data_in_buffer[1].genblk1[1].genblk2.inv_last  (.A(\data_in_buffer[1].genblk1[1].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\data_in_buffer[1].X ));
 sky130_fd_sc_hd__inv_1 \data_in_buffer[2].genblk1[0].genblk1.inv_first  (.A(\data_in_buffer[2].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\data_in_buffer[2].genblk1[0].mid ));
 sky130_fd_sc_hd__inv_1 \data_in_buffer[2].genblk1[0].genblk2.inv2  (.A(\data_in_buffer[2].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\data_in_buffer[2].b[0] ));
 sky130_fd_sc_hd__inv_1 \data_in_buffer[2].genblk1[1].genblk1.inv1  (.A(\data_in_buffer[2].b[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\data_in_buffer[2].genblk1[1].mid ));
 sky130_fd_sc_hd__inv_2 \data_in_buffer[2].genblk1[1].genblk2.inv_last  (.A(\data_in_buffer[2].genblk1[1].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\data_in_buffer[2].X ));
 sky130_fd_sc_hd__inv_1 \data_in_buffer[3].genblk1[0].genblk1.inv_first  (.A(\data_in_buffer[3].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\data_in_buffer[3].genblk1[0].mid ));
 sky130_fd_sc_hd__inv_1 \data_in_buffer[3].genblk1[0].genblk2.inv2  (.A(\data_in_buffer[3].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\data_in_buffer[3].b[0] ));
 sky130_fd_sc_hd__inv_1 \data_in_buffer[3].genblk1[1].genblk1.inv1  (.A(\data_in_buffer[3].b[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\data_in_buffer[3].genblk1[1].mid ));
 sky130_fd_sc_hd__inv_2 \data_in_buffer[3].genblk1[1].genblk2.inv_last  (.A(\data_in_buffer[3].genblk1[1].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\data_in_buffer[3].X ));
 sky130_fd_sc_hd__inv_1 \data_in_buffer[4].genblk1[0].genblk1.inv_first  (.A(\data_in_buffer[4].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\data_in_buffer[4].genblk1[0].mid ));
 sky130_fd_sc_hd__inv_1 \data_in_buffer[4].genblk1[0].genblk2.inv2  (.A(\data_in_buffer[4].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\data_in_buffer[4].b[0] ));
 sky130_fd_sc_hd__inv_1 \data_in_buffer[4].genblk1[1].genblk1.inv1  (.A(\data_in_buffer[4].b[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\data_in_buffer[4].genblk1[1].mid ));
 sky130_fd_sc_hd__inv_2 \data_in_buffer[4].genblk1[1].genblk2.inv_last  (.A(\data_in_buffer[4].genblk1[1].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\data_in_buffer[4].X ));
 sky130_fd_sc_hd__inv_1 \data_in_buffer[5].genblk1[0].genblk1.inv_first  (.A(\data_in_buffer[5].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\data_in_buffer[5].genblk1[0].mid ));
 sky130_fd_sc_hd__inv_1 \data_in_buffer[5].genblk1[0].genblk2.inv2  (.A(\data_in_buffer[5].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\data_in_buffer[5].b[0] ));
 sky130_fd_sc_hd__inv_1 \data_in_buffer[5].genblk1[1].genblk1.inv1  (.A(\data_in_buffer[5].b[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\data_in_buffer[5].genblk1[1].mid ));
 sky130_fd_sc_hd__inv_2 \data_in_buffer[5].genblk1[1].genblk2.inv_last  (.A(\data_in_buffer[5].genblk1[1].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\data_in_buffer[5].X ));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout10 (.A(net11),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net10));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout11 (.A(net21),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net11));
 sky130_fd_sc_hd__buf_2 fanout12 (.A(net21),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net12));
 sky130_fd_sc_hd__buf_2 fanout13 (.A(net16),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net13));
 sky130_fd_sc_hd__buf_2 fanout14 (.A(net16),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net14));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout15 (.A(net16),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net15));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout16 (.A(net21),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net16));
 sky130_fd_sc_hd__buf_2 fanout17 (.A(net20),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net17));
 sky130_fd_sc_hd__buf_2 fanout18 (.A(net20),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net18));
 sky130_fd_sc_hd__clkbuf_2 fanout19 (.A(net20),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net19));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout20 (.A(net21),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net20));
 sky130_fd_sc_hd__clkbuf_2 fanout21 (.A(net22),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net21));
 sky130_fd_sc_hd__buf_2 fanout22 (.A(net49),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net22));
 sky130_fd_sc_hd__buf_2 fanout23 (.A(net24),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net23));
 sky130_fd_sc_hd__buf_2 fanout24 (.A(net25),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net24));
 sky130_fd_sc_hd__clkbuf_2 fanout25 (.A(net49),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net25));
 sky130_fd_sc_hd__buf_2 fanout26 (.A(net32),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net26));
 sky130_fd_sc_hd__buf_2 fanout27 (.A(net32),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net27));
 sky130_fd_sc_hd__buf_2 fanout28 (.A(net32),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net28));
 sky130_fd_sc_hd__clkbuf_2 fanout29 (.A(net32),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net29));
 sky130_fd_sc_hd__buf_2 fanout30 (.A(net32),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net30));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout31 (.A(net32),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net31));
 sky130_fd_sc_hd__buf_2 fanout32 (.A(net49),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net32));
 sky130_fd_sc_hd__buf_2 fanout33 (.A(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net33));
 sky130_fd_sc_hd__buf_2 fanout34 (.A(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net34));
 sky130_fd_sc_hd__clkbuf_2 fanout35 (.A(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net35));
 sky130_fd_sc_hd__clkbuf_2 fanout36 (.A(net41),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net36));
 sky130_fd_sc_hd__buf_2 fanout37 (.A(net41),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net37));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout38 (.A(net41),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net38));
 sky130_fd_sc_hd__buf_2 fanout39 (.A(net41),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net39));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout40 (.A(net41),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net40));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout41 (.A(net49),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net41));
 sky130_fd_sc_hd__buf_2 fanout42 (.A(net48),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net42));
 sky130_fd_sc_hd__buf_2 fanout43 (.A(net48),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net43));
 sky130_fd_sc_hd__buf_2 fanout44 (.A(net48),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net44));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout45 (.A(net48),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net45));
 sky130_fd_sc_hd__buf_2 fanout46 (.A(net48),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net46));
 sky130_fd_sc_hd__buf_2 fanout47 (.A(net48),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net47));
 sky130_fd_sc_hd__buf_2 fanout48 (.A(net49),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net48));
 sky130_fd_sc_hd__clkbuf_2 fanout49 (.A(\f_fifo.reset_n ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net49));
 sky130_fd_sc_hd__buf_2 fanout8 (.A(net11),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net8));
 sky130_fd_sc_hd__buf_2 fanout9 (.A(net11),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net9));
 sky130_fd_sc_hd__buf_2 input1 (.A(io_in[1]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_1 input2 (.A(io_in[2]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_1 input3 (.A(io_in[3]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net3));
 sky130_fd_sc_hd__dlymetal6s2s_1 input4 (.A(io_in[4]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_1 input5 (.A(io_in[5]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_1 input6 (.A(io_in[6]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_1 input7 (.A(io_in[7]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net7));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[0].entry.input_buf[0].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[0].entry.input_buf[0].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[0].entry.input_buf[0].genblk1[0].mid ));
 sky130_fd_sc_hd__inv_2 \l_fifo.genblk1[0].entry.input_buf[0].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[0].entry.input_buf[0].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[0].entry.input_buf[0].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[0].entry.input_buf[1].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[0].entry.input_buf[1].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[0].entry.input_buf[1].genblk1[0].mid ));
 sky130_fd_sc_hd__inv_2 \l_fifo.genblk1[0].entry.input_buf[1].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[0].entry.input_buf[1].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[0].entry.input_buf[1].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[0].entry.input_buf[2].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[0].entry.input_buf[2].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[0].entry.input_buf[2].genblk1[0].mid ));
 sky130_fd_sc_hd__clkinv_2 \l_fifo.genblk1[0].entry.input_buf[2].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[0].entry.input_buf[2].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[0].entry.input_buf[2].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[0].entry.input_buf[3].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[0].entry.input_buf[3].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[0].entry.input_buf[3].genblk1[0].mid ));
 sky130_fd_sc_hd__clkinv_2 \l_fifo.genblk1[0].entry.input_buf[3].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[0].entry.input_buf[3].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[0].entry.input_buf[3].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[0].entry.input_buf[4].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[0].entry.input_buf[4].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[0].entry.input_buf[4].genblk1[0].mid ));
 sky130_fd_sc_hd__clkinv_2 \l_fifo.genblk1[0].entry.input_buf[4].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[0].entry.input_buf[4].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[0].entry.input_buf[4].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[0].entry.input_buf[5].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[0].entry.input_buf[5].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[0].entry.input_buf[5].genblk1[0].mid ));
 sky130_fd_sc_hd__inv_2 \l_fifo.genblk1[0].entry.input_buf[5].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[0].entry.input_buf[5].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[0].entry.input_buf[5].X ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[0].entry.latch[0]  (.D(\l_fifo.genblk1[0].entry.input_buf[0].X ),
    .GATE(\l_fifo.genblk1[0].entry.empty ),
    .RESET_B(net22),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\f_fifo.data_in[0] ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[0].entry.latch[1]  (.D(\l_fifo.genblk1[0].entry.input_buf[1].X ),
    .GATE(\l_fifo.genblk1[0].entry.empty ),
    .RESET_B(net24),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\f_fifo.data_in[1] ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[0].entry.latch[2]  (.D(\l_fifo.genblk1[0].entry.input_buf[2].X ),
    .GATE(\l_fifo.genblk1[0].entry.empty ),
    .RESET_B(net23),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\f_fifo.data_in[2] ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[0].entry.latch[3]  (.D(\l_fifo.genblk1[0].entry.input_buf[3].X ),
    .GATE(\l_fifo.genblk1[0].entry.empty ),
    .RESET_B(net22),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\f_fifo.data_in[3] ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[0].entry.latch[4]  (.D(\l_fifo.genblk1[0].entry.input_buf[4].X ),
    .GATE(\l_fifo.genblk1[0].entry.empty ),
    .RESET_B(net23),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\f_fifo.data_in[4] ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[0].entry.latch[5]  (.D(\l_fifo.genblk1[0].entry.input_buf[5].X ),
    .GATE(\l_fifo.genblk1[0].entry.empty ),
    .RESET_B(net23),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\f_fifo.data_in[5] ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[10].entry.input_buf[0].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[10].entry.input_buf[0].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[10].entry.input_buf[0].genblk1[0].mid ));
 sky130_fd_sc_hd__clkinv_2 \l_fifo.genblk1[10].entry.input_buf[0].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[10].entry.input_buf[0].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[10].entry.input_buf[0].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[10].entry.input_buf[1].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[10].entry.input_buf[1].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[10].entry.input_buf[1].genblk1[0].mid ));
 sky130_fd_sc_hd__inv_2 \l_fifo.genblk1[10].entry.input_buf[1].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[10].entry.input_buf[1].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[10].entry.input_buf[1].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[10].entry.input_buf[2].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[10].entry.input_buf[2].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[10].entry.input_buf[2].genblk1[0].mid ));
 sky130_fd_sc_hd__inv_2 \l_fifo.genblk1[10].entry.input_buf[2].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[10].entry.input_buf[2].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[10].entry.input_buf[2].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[10].entry.input_buf[3].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[10].entry.input_buf[3].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[10].entry.input_buf[3].genblk1[0].mid ));
 sky130_fd_sc_hd__clkinv_2 \l_fifo.genblk1[10].entry.input_buf[3].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[10].entry.input_buf[3].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[10].entry.input_buf[3].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[10].entry.input_buf[4].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[10].entry.input_buf[4].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[10].entry.input_buf[4].genblk1[0].mid ));
 sky130_fd_sc_hd__clkinv_2 \l_fifo.genblk1[10].entry.input_buf[4].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[10].entry.input_buf[4].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[10].entry.input_buf[4].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[10].entry.input_buf[5].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[10].entry.input_buf[5].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[10].entry.input_buf[5].genblk1[0].mid ));
 sky130_fd_sc_hd__clkinv_2 \l_fifo.genblk1[10].entry.input_buf[5].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[10].entry.input_buf[5].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[10].entry.input_buf[5].X ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[10].entry.latch[0]  (.D(\l_fifo.genblk1[10].entry.input_buf[0].X ),
    .GATE(\l_fifo.genblk1[10].entry.empty ),
    .RESET_B(net42),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[9].entry.input_buf[0].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[10].entry.latch[1]  (.D(\l_fifo.genblk1[10].entry.input_buf[1].X ),
    .GATE(\l_fifo.genblk1[10].entry.empty ),
    .RESET_B(net42),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[9].entry.input_buf[1].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[10].entry.latch[2]  (.D(\l_fifo.genblk1[10].entry.input_buf[2].X ),
    .GATE(\l_fifo.genblk1[10].entry.empty ),
    .RESET_B(net42),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[9].entry.input_buf[2].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[10].entry.latch[3]  (.D(\l_fifo.genblk1[10].entry.input_buf[3].X ),
    .GATE(\l_fifo.genblk1[10].entry.empty ),
    .RESET_B(net44),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[9].entry.input_buf[3].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[10].entry.latch[4]  (.D(\l_fifo.genblk1[10].entry.input_buf[4].X ),
    .GATE(\l_fifo.genblk1[10].entry.empty ),
    .RESET_B(net42),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[9].entry.input_buf[4].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[10].entry.latch[5]  (.D(\l_fifo.genblk1[10].entry.input_buf[5].X ),
    .GATE(\l_fifo.genblk1[10].entry.empty ),
    .RESET_B(net30),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[9].entry.input_buf[5].A ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[11].entry.input_buf[0].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[11].entry.input_buf[0].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[11].entry.input_buf[0].genblk1[0].mid ));
 sky130_fd_sc_hd__inv_2 \l_fifo.genblk1[11].entry.input_buf[0].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[11].entry.input_buf[0].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[11].entry.input_buf[0].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[11].entry.input_buf[1].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[11].entry.input_buf[1].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[11].entry.input_buf[1].genblk1[0].mid ));
 sky130_fd_sc_hd__clkinv_2 \l_fifo.genblk1[11].entry.input_buf[1].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[11].entry.input_buf[1].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[11].entry.input_buf[1].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[11].entry.input_buf[2].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[11].entry.input_buf[2].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[11].entry.input_buf[2].genblk1[0].mid ));
 sky130_fd_sc_hd__clkinv_2 \l_fifo.genblk1[11].entry.input_buf[2].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[11].entry.input_buf[2].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[11].entry.input_buf[2].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[11].entry.input_buf[3].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[11].entry.input_buf[3].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[11].entry.input_buf[3].genblk1[0].mid ));
 sky130_fd_sc_hd__clkinv_2 \l_fifo.genblk1[11].entry.input_buf[3].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[11].entry.input_buf[3].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[11].entry.input_buf[3].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[11].entry.input_buf[4].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[11].entry.input_buf[4].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[11].entry.input_buf[4].genblk1[0].mid ));
 sky130_fd_sc_hd__inv_2 \l_fifo.genblk1[11].entry.input_buf[4].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[11].entry.input_buf[4].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[11].entry.input_buf[4].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[11].entry.input_buf[5].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[11].entry.input_buf[5].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[11].entry.input_buf[5].genblk1[0].mid ));
 sky130_fd_sc_hd__clkinv_2 \l_fifo.genblk1[11].entry.input_buf[5].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[11].entry.input_buf[5].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[11].entry.input_buf[5].X ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[11].entry.latch[0]  (.D(\l_fifo.genblk1[11].entry.input_buf[0].X ),
    .GATE(\l_fifo.genblk1[11].entry.empty ),
    .RESET_B(net42),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[10].entry.input_buf[0].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[11].entry.latch[1]  (.D(\l_fifo.genblk1[11].entry.input_buf[1].X ),
    .GATE(\l_fifo.genblk1[11].entry.empty ),
    .RESET_B(net44),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[10].entry.input_buf[1].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[11].entry.latch[2]  (.D(\l_fifo.genblk1[11].entry.input_buf[2].X ),
    .GATE(\l_fifo.genblk1[11].entry.empty ),
    .RESET_B(net44),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[10].entry.input_buf[2].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[11].entry.latch[3]  (.D(\l_fifo.genblk1[11].entry.input_buf[3].X ),
    .GATE(\l_fifo.genblk1[11].entry.empty ),
    .RESET_B(net44),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[10].entry.input_buf[3].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[11].entry.latch[4]  (.D(\l_fifo.genblk1[11].entry.input_buf[4].X ),
    .GATE(\l_fifo.genblk1[11].entry.empty ),
    .RESET_B(net31),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[10].entry.input_buf[4].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[11].entry.latch[5]  (.D(\l_fifo.genblk1[11].entry.input_buf[5].X ),
    .GATE(\l_fifo.genblk1[11].entry.empty ),
    .RESET_B(net29),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[10].entry.input_buf[5].A ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[12].entry.input_buf[0].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[12].entry.input_buf[0].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[12].entry.input_buf[0].genblk1[0].mid ));
 sky130_fd_sc_hd__inv_2 \l_fifo.genblk1[12].entry.input_buf[0].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[12].entry.input_buf[0].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[12].entry.input_buf[0].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[12].entry.input_buf[1].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[12].entry.input_buf[1].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[12].entry.input_buf[1].genblk1[0].mid ));
 sky130_fd_sc_hd__inv_2 \l_fifo.genblk1[12].entry.input_buf[1].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[12].entry.input_buf[1].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[12].entry.input_buf[1].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[12].entry.input_buf[2].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[12].entry.input_buf[2].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[12].entry.input_buf[2].genblk1[0].mid ));
 sky130_fd_sc_hd__clkinv_2 \l_fifo.genblk1[12].entry.input_buf[2].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[12].entry.input_buf[2].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[12].entry.input_buf[2].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[12].entry.input_buf[3].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[12].entry.input_buf[3].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[12].entry.input_buf[3].genblk1[0].mid ));
 sky130_fd_sc_hd__clkinv_2 \l_fifo.genblk1[12].entry.input_buf[3].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[12].entry.input_buf[3].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[12].entry.input_buf[3].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[12].entry.input_buf[4].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[12].entry.input_buf[4].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[12].entry.input_buf[4].genblk1[0].mid ));
 sky130_fd_sc_hd__clkinv_2 \l_fifo.genblk1[12].entry.input_buf[4].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[12].entry.input_buf[4].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[12].entry.input_buf[4].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[12].entry.input_buf[5].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[12].entry.input_buf[5].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[12].entry.input_buf[5].genblk1[0].mid ));
 sky130_fd_sc_hd__inv_2 \l_fifo.genblk1[12].entry.input_buf[5].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[12].entry.input_buf[5].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[12].entry.input_buf[5].X ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[12].entry.latch[0]  (.D(\l_fifo.genblk1[12].entry.input_buf[0].X ),
    .GATE(\l_fifo.genblk1[12].entry.empty ),
    .RESET_B(net44),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[11].entry.input_buf[0].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[12].entry.latch[1]  (.D(\l_fifo.genblk1[12].entry.input_buf[1].X ),
    .GATE(\l_fifo.genblk1[12].entry.empty ),
    .RESET_B(net30),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[11].entry.input_buf[1].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[12].entry.latch[2]  (.D(\l_fifo.genblk1[12].entry.input_buf[2].X ),
    .GATE(\l_fifo.genblk1[12].entry.empty ),
    .RESET_B(net43),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[11].entry.input_buf[2].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[12].entry.latch[3]  (.D(\l_fifo.genblk1[12].entry.input_buf[3].X ),
    .GATE(\l_fifo.genblk1[12].entry.empty ),
    .RESET_B(net44),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[11].entry.input_buf[3].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[12].entry.latch[4]  (.D(\l_fifo.genblk1[12].entry.input_buf[4].X ),
    .GATE(\l_fifo.genblk1[12].entry.empty ),
    .RESET_B(net31),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[11].entry.input_buf[4].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[12].entry.latch[5]  (.D(\l_fifo.genblk1[12].entry.input_buf[5].X ),
    .GATE(\l_fifo.genblk1[12].entry.empty ),
    .RESET_B(net44),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[11].entry.input_buf[5].A ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[13].entry.input_buf[0].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[13].entry.input_buf[0].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[13].entry.input_buf[0].genblk1[0].mid ));
 sky130_fd_sc_hd__inv_2 \l_fifo.genblk1[13].entry.input_buf[0].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[13].entry.input_buf[0].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[13].entry.input_buf[0].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[13].entry.input_buf[1].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[13].entry.input_buf[1].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[13].entry.input_buf[1].genblk1[0].mid ));
 sky130_fd_sc_hd__inv_2 \l_fifo.genblk1[13].entry.input_buf[1].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[13].entry.input_buf[1].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[13].entry.input_buf[1].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[13].entry.input_buf[2].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[13].entry.input_buf[2].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[13].entry.input_buf[2].genblk1[0].mid ));
 sky130_fd_sc_hd__inv_2 \l_fifo.genblk1[13].entry.input_buf[2].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[13].entry.input_buf[2].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[13].entry.input_buf[2].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[13].entry.input_buf[3].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[13].entry.input_buf[3].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[13].entry.input_buf[3].genblk1[0].mid ));
 sky130_fd_sc_hd__clkinv_2 \l_fifo.genblk1[13].entry.input_buf[3].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[13].entry.input_buf[3].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[13].entry.input_buf[3].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[13].entry.input_buf[4].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[13].entry.input_buf[4].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[13].entry.input_buf[4].genblk1[0].mid ));
 sky130_fd_sc_hd__inv_2 \l_fifo.genblk1[13].entry.input_buf[4].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[13].entry.input_buf[4].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[13].entry.input_buf[4].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[13].entry.input_buf[5].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[13].entry.input_buf[5].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[13].entry.input_buf[5].genblk1[0].mid ));
 sky130_fd_sc_hd__clkinv_2 \l_fifo.genblk1[13].entry.input_buf[5].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[13].entry.input_buf[5].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[13].entry.input_buf[5].X ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[13].entry.latch[0]  (.D(\l_fifo.genblk1[13].entry.input_buf[0].X ),
    .GATE(\l_fifo.genblk1[13].entry.empty ),
    .RESET_B(net44),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[12].entry.input_buf[0].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[13].entry.latch[1]  (.D(\l_fifo.genblk1[13].entry.input_buf[1].X ),
    .GATE(\l_fifo.genblk1[13].entry.empty ),
    .RESET_B(net44),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[12].entry.input_buf[1].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[13].entry.latch[2]  (.D(\l_fifo.genblk1[13].entry.input_buf[2].X ),
    .GATE(\l_fifo.genblk1[13].entry.empty ),
    .RESET_B(net43),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[12].entry.input_buf[2].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[13].entry.latch[3]  (.D(\l_fifo.genblk1[13].entry.input_buf[3].X ),
    .GATE(\l_fifo.genblk1[13].entry.empty ),
    .RESET_B(net44),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[12].entry.input_buf[3].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[13].entry.latch[4]  (.D(\l_fifo.genblk1[13].entry.input_buf[4].X ),
    .GATE(\l_fifo.genblk1[13].entry.empty ),
    .RESET_B(net43),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[12].entry.input_buf[4].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[13].entry.latch[5]  (.D(\l_fifo.genblk1[13].entry.input_buf[5].X ),
    .GATE(\l_fifo.genblk1[13].entry.empty ),
    .RESET_B(net45),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[12].entry.input_buf[5].A ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[14].entry.input_buf[0].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[14].entry.input_buf[0].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[14].entry.input_buf[0].genblk1[0].mid ));
 sky130_fd_sc_hd__inv_2 \l_fifo.genblk1[14].entry.input_buf[0].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[14].entry.input_buf[0].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[14].entry.input_buf[0].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[14].entry.input_buf[1].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[14].entry.input_buf[1].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[14].entry.input_buf[1].genblk1[0].mid ));
 sky130_fd_sc_hd__clkinv_2 \l_fifo.genblk1[14].entry.input_buf[1].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[14].entry.input_buf[1].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[14].entry.input_buf[1].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[14].entry.input_buf[2].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[14].entry.input_buf[2].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[14].entry.input_buf[2].genblk1[0].mid ));
 sky130_fd_sc_hd__clkinv_2 \l_fifo.genblk1[14].entry.input_buf[2].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[14].entry.input_buf[2].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[14].entry.input_buf[2].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[14].entry.input_buf[3].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[14].entry.input_buf[3].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[14].entry.input_buf[3].genblk1[0].mid ));
 sky130_fd_sc_hd__inv_2 \l_fifo.genblk1[14].entry.input_buf[3].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[14].entry.input_buf[3].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[14].entry.input_buf[3].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[14].entry.input_buf[4].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[14].entry.input_buf[4].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[14].entry.input_buf[4].genblk1[0].mid ));
 sky130_fd_sc_hd__inv_2 \l_fifo.genblk1[14].entry.input_buf[4].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[14].entry.input_buf[4].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[14].entry.input_buf[4].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[14].entry.input_buf[5].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[14].entry.input_buf[5].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[14].entry.input_buf[5].genblk1[0].mid ));
 sky130_fd_sc_hd__inv_2 \l_fifo.genblk1[14].entry.input_buf[5].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[14].entry.input_buf[5].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[14].entry.input_buf[5].X ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[14].entry.latch[0]  (.D(\l_fifo.genblk1[14].entry.input_buf[0].X ),
    .GATE(\l_fifo.genblk1[14].entry.empty ),
    .RESET_B(net45),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[13].entry.input_buf[0].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[14].entry.latch[1]  (.D(\l_fifo.genblk1[14].entry.input_buf[1].X ),
    .GATE(\l_fifo.genblk1[14].entry.empty ),
    .RESET_B(net45),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[13].entry.input_buf[1].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[14].entry.latch[2]  (.D(\l_fifo.genblk1[14].entry.input_buf[2].X ),
    .GATE(\l_fifo.genblk1[14].entry.empty ),
    .RESET_B(net43),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[13].entry.input_buf[2].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[14].entry.latch[3]  (.D(\l_fifo.genblk1[14].entry.input_buf[3].X ),
    .GATE(\l_fifo.genblk1[14].entry.empty ),
    .RESET_B(net45),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[13].entry.input_buf[3].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[14].entry.latch[4]  (.D(\l_fifo.genblk1[14].entry.input_buf[4].X ),
    .GATE(\l_fifo.genblk1[14].entry.empty ),
    .RESET_B(net39),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[13].entry.input_buf[4].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[14].entry.latch[5]  (.D(\l_fifo.genblk1[14].entry.input_buf[5].X ),
    .GATE(\l_fifo.genblk1[14].entry.empty ),
    .RESET_B(net47),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[13].entry.input_buf[5].A ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[15].entry.input_buf[0].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[15].entry.input_buf[0].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[15].entry.input_buf[0].genblk1[0].mid ));
 sky130_fd_sc_hd__clkinv_2 \l_fifo.genblk1[15].entry.input_buf[0].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[15].entry.input_buf[0].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[15].entry.input_buf[0].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[15].entry.input_buf[1].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[15].entry.input_buf[1].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[15].entry.input_buf[1].genblk1[0].mid ));
 sky130_fd_sc_hd__inv_2 \l_fifo.genblk1[15].entry.input_buf[1].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[15].entry.input_buf[1].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[15].entry.input_buf[1].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[15].entry.input_buf[2].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[15].entry.input_buf[2].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[15].entry.input_buf[2].genblk1[0].mid ));
 sky130_fd_sc_hd__inv_2 \l_fifo.genblk1[15].entry.input_buf[2].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[15].entry.input_buf[2].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[15].entry.input_buf[2].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[15].entry.input_buf[3].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[15].entry.input_buf[3].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[15].entry.input_buf[3].genblk1[0].mid ));
 sky130_fd_sc_hd__inv_2 \l_fifo.genblk1[15].entry.input_buf[3].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[15].entry.input_buf[3].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[15].entry.input_buf[3].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[15].entry.input_buf[4].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[15].entry.input_buf[4].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[15].entry.input_buf[4].genblk1[0].mid ));
 sky130_fd_sc_hd__inv_2 \l_fifo.genblk1[15].entry.input_buf[4].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[15].entry.input_buf[4].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[15].entry.input_buf[4].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[15].entry.input_buf[5].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[15].entry.input_buf[5].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[15].entry.input_buf[5].genblk1[0].mid ));
 sky130_fd_sc_hd__inv_2 \l_fifo.genblk1[15].entry.input_buf[5].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[15].entry.input_buf[5].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[15].entry.input_buf[5].X ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[15].entry.latch[0]  (.D(\l_fifo.genblk1[15].entry.input_buf[0].X ),
    .GATE(\l_fifo.genblk1[15].entry.empty ),
    .RESET_B(net47),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[14].entry.input_buf[0].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[15].entry.latch[1]  (.D(\l_fifo.genblk1[15].entry.input_buf[1].X ),
    .GATE(\l_fifo.genblk1[15].entry.empty ),
    .RESET_B(net45),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[14].entry.input_buf[1].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[15].entry.latch[2]  (.D(\l_fifo.genblk1[15].entry.input_buf[2].X ),
    .GATE(\l_fifo.genblk1[15].entry.empty ),
    .RESET_B(net43),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[14].entry.input_buf[2].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[15].entry.latch[3]  (.D(\l_fifo.genblk1[15].entry.input_buf[3].X ),
    .GATE(\l_fifo.genblk1[15].entry.empty ),
    .RESET_B(net47),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[14].entry.input_buf[3].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[15].entry.latch[4]  (.D(\l_fifo.genblk1[15].entry.input_buf[4].X ),
    .GATE(\l_fifo.genblk1[15].entry.empty ),
    .RESET_B(net39),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[14].entry.input_buf[4].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[15].entry.latch[5]  (.D(\l_fifo.genblk1[15].entry.input_buf[5].X ),
    .GATE(\l_fifo.genblk1[15].entry.empty ),
    .RESET_B(net47),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[14].entry.input_buf[5].A ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[16].entry.input_buf[0].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[16].entry.input_buf[0].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[16].entry.input_buf[0].genblk1[0].mid ));
 sky130_fd_sc_hd__inv_2 \l_fifo.genblk1[16].entry.input_buf[0].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[16].entry.input_buf[0].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[16].entry.input_buf[0].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[16].entry.input_buf[1].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[16].entry.input_buf[1].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[16].entry.input_buf[1].genblk1[0].mid ));
 sky130_fd_sc_hd__clkinv_2 \l_fifo.genblk1[16].entry.input_buf[1].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[16].entry.input_buf[1].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[16].entry.input_buf[1].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[16].entry.input_buf[2].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[16].entry.input_buf[2].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[16].entry.input_buf[2].genblk1[0].mid ));
 sky130_fd_sc_hd__clkinv_2 \l_fifo.genblk1[16].entry.input_buf[2].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[16].entry.input_buf[2].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[16].entry.input_buf[2].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[16].entry.input_buf[3].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[16].entry.input_buf[3].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[16].entry.input_buf[3].genblk1[0].mid ));
 sky130_fd_sc_hd__clkinv_2 \l_fifo.genblk1[16].entry.input_buf[3].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[16].entry.input_buf[3].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[16].entry.input_buf[3].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[16].entry.input_buf[4].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[16].entry.input_buf[4].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[16].entry.input_buf[4].genblk1[0].mid ));
 sky130_fd_sc_hd__clkinv_2 \l_fifo.genblk1[16].entry.input_buf[4].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[16].entry.input_buf[4].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[16].entry.input_buf[4].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[16].entry.input_buf[5].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[16].entry.input_buf[5].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[16].entry.input_buf[5].genblk1[0].mid ));
 sky130_fd_sc_hd__inv_2 \l_fifo.genblk1[16].entry.input_buf[5].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[16].entry.input_buf[5].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[16].entry.input_buf[5].X ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[16].entry.latch[0]  (.D(\l_fifo.genblk1[16].entry.input_buf[0].X ),
    .GATE(\l_fifo.genblk1[16].entry.empty ),
    .RESET_B(net47),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[15].entry.input_buf[0].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[16].entry.latch[1]  (.D(\l_fifo.genblk1[16].entry.input_buf[1].X ),
    .GATE(\l_fifo.genblk1[16].entry.empty ),
    .RESET_B(net46),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[15].entry.input_buf[1].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[16].entry.latch[2]  (.D(\l_fifo.genblk1[16].entry.input_buf[2].X ),
    .GATE(\l_fifo.genblk1[16].entry.empty ),
    .RESET_B(net46),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[15].entry.input_buf[2].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[16].entry.latch[3]  (.D(\l_fifo.genblk1[16].entry.input_buf[3].X ),
    .GATE(\l_fifo.genblk1[16].entry.empty ),
    .RESET_B(net48),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[15].entry.input_buf[3].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[16].entry.latch[4]  (.D(\l_fifo.genblk1[16].entry.input_buf[4].X ),
    .GATE(\l_fifo.genblk1[16].entry.empty ),
    .RESET_B(net46),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[15].entry.input_buf[4].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[16].entry.latch[5]  (.D(\l_fifo.genblk1[16].entry.input_buf[5].X ),
    .GATE(\l_fifo.genblk1[16].entry.empty ),
    .RESET_B(net47),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[15].entry.input_buf[5].A ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[17].entry.input_buf[0].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[17].entry.input_buf[0].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[17].entry.input_buf[0].genblk1[0].mid ));
 sky130_fd_sc_hd__inv_2 \l_fifo.genblk1[17].entry.input_buf[0].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[17].entry.input_buf[0].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[17].entry.input_buf[0].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[17].entry.input_buf[1].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[17].entry.input_buf[1].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[17].entry.input_buf[1].genblk1[0].mid ));
 sky130_fd_sc_hd__inv_2 \l_fifo.genblk1[17].entry.input_buf[1].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[17].entry.input_buf[1].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[17].entry.input_buf[1].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[17].entry.input_buf[2].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[17].entry.input_buf[2].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[17].entry.input_buf[2].genblk1[0].mid ));
 sky130_fd_sc_hd__inv_2 \l_fifo.genblk1[17].entry.input_buf[2].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[17].entry.input_buf[2].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[17].entry.input_buf[2].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[17].entry.input_buf[3].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[17].entry.input_buf[3].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[17].entry.input_buf[3].genblk1[0].mid ));
 sky130_fd_sc_hd__inv_2 \l_fifo.genblk1[17].entry.input_buf[3].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[17].entry.input_buf[3].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[17].entry.input_buf[3].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[17].entry.input_buf[4].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[17].entry.input_buf[4].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[17].entry.input_buf[4].genblk1[0].mid ));
 sky130_fd_sc_hd__inv_2 \l_fifo.genblk1[17].entry.input_buf[4].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[17].entry.input_buf[4].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[17].entry.input_buf[4].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[17].entry.input_buf[5].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[17].entry.input_buf[5].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[17].entry.input_buf[5].genblk1[0].mid ));
 sky130_fd_sc_hd__inv_2 \l_fifo.genblk1[17].entry.input_buf[5].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[17].entry.input_buf[5].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[17].entry.input_buf[5].X ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[17].entry.latch[0]  (.D(\l_fifo.genblk1[17].entry.input_buf[0].X ),
    .GATE(\l_fifo.genblk1[17].entry.empty ),
    .RESET_B(net47),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[16].entry.input_buf[0].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[17].entry.latch[1]  (.D(\l_fifo.genblk1[17].entry.input_buf[1].X ),
    .GATE(\l_fifo.genblk1[17].entry.empty ),
    .RESET_B(net46),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[16].entry.input_buf[1].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[17].entry.latch[2]  (.D(\l_fifo.genblk1[17].entry.input_buf[2].X ),
    .GATE(\l_fifo.genblk1[17].entry.empty ),
    .RESET_B(net47),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[16].entry.input_buf[2].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[17].entry.latch[3]  (.D(\l_fifo.genblk1[17].entry.input_buf[3].X ),
    .GATE(\l_fifo.genblk1[17].entry.empty ),
    .RESET_B(net47),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[16].entry.input_buf[3].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[17].entry.latch[4]  (.D(\l_fifo.genblk1[17].entry.input_buf[4].X ),
    .GATE(\l_fifo.genblk1[17].entry.empty ),
    .RESET_B(net47),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[16].entry.input_buf[4].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[17].entry.latch[5]  (.D(\l_fifo.genblk1[17].entry.input_buf[5].X ),
    .GATE(\l_fifo.genblk1[17].entry.empty ),
    .RESET_B(net46),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[16].entry.input_buf[5].A ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[18].entry.input_buf[0].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[18].entry.input_buf[0].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[18].entry.input_buf[0].genblk1[0].mid ));
 sky130_fd_sc_hd__clkinv_2 \l_fifo.genblk1[18].entry.input_buf[0].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[18].entry.input_buf[0].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[18].entry.input_buf[0].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[18].entry.input_buf[1].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[18].entry.input_buf[1].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[18].entry.input_buf[1].genblk1[0].mid ));
 sky130_fd_sc_hd__clkinv_2 \l_fifo.genblk1[18].entry.input_buf[1].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[18].entry.input_buf[1].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[18].entry.input_buf[1].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[18].entry.input_buf[2].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[18].entry.input_buf[2].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[18].entry.input_buf[2].genblk1[0].mid ));
 sky130_fd_sc_hd__clkinv_2 \l_fifo.genblk1[18].entry.input_buf[2].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[18].entry.input_buf[2].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[18].entry.input_buf[2].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[18].entry.input_buf[3].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[18].entry.input_buf[3].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[18].entry.input_buf[3].genblk1[0].mid ));
 sky130_fd_sc_hd__clkinv_2 \l_fifo.genblk1[18].entry.input_buf[3].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[18].entry.input_buf[3].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[18].entry.input_buf[3].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[18].entry.input_buf[4].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[18].entry.input_buf[4].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[18].entry.input_buf[4].genblk1[0].mid ));
 sky130_fd_sc_hd__inv_2 \l_fifo.genblk1[18].entry.input_buf[4].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[18].entry.input_buf[4].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[18].entry.input_buf[4].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[18].entry.input_buf[5].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[18].entry.input_buf[5].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[18].entry.input_buf[5].genblk1[0].mid ));
 sky130_fd_sc_hd__clkinv_2 \l_fifo.genblk1[18].entry.input_buf[5].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[18].entry.input_buf[5].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[18].entry.input_buf[5].X ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[18].entry.latch[0]  (.D(\l_fifo.genblk1[18].entry.input_buf[0].X ),
    .GATE(\l_fifo.genblk1[18].entry.empty ),
    .RESET_B(net39),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[17].entry.input_buf[0].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[18].entry.latch[1]  (.D(\l_fifo.genblk1[18].entry.input_buf[1].X ),
    .GATE(\l_fifo.genblk1[18].entry.empty ),
    .RESET_B(net39),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[17].entry.input_buf[1].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[18].entry.latch[2]  (.D(\l_fifo.genblk1[18].entry.input_buf[2].X ),
    .GATE(\l_fifo.genblk1[18].entry.empty ),
    .RESET_B(net46),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[17].entry.input_buf[2].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[18].entry.latch[3]  (.D(\l_fifo.genblk1[18].entry.input_buf[3].X ),
    .GATE(\l_fifo.genblk1[18].entry.empty ),
    .RESET_B(net46),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[17].entry.input_buf[3].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[18].entry.latch[4]  (.D(\l_fifo.genblk1[18].entry.input_buf[4].X ),
    .GATE(\l_fifo.genblk1[18].entry.empty ),
    .RESET_B(net46),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[17].entry.input_buf[4].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[18].entry.latch[5]  (.D(\l_fifo.genblk1[18].entry.input_buf[5].X ),
    .GATE(\l_fifo.genblk1[18].entry.empty ),
    .RESET_B(net43),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[17].entry.input_buf[5].A ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[19].entry.input_buf[0].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[19].entry.input_buf[0].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[19].entry.input_buf[0].genblk1[0].mid ));
 sky130_fd_sc_hd__inv_2 \l_fifo.genblk1[19].entry.input_buf[0].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[19].entry.input_buf[0].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[19].entry.input_buf[0].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[19].entry.input_buf[1].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[19].entry.input_buf[1].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[19].entry.input_buf[1].genblk1[0].mid ));
 sky130_fd_sc_hd__clkinv_2 \l_fifo.genblk1[19].entry.input_buf[1].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[19].entry.input_buf[1].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[19].entry.input_buf[1].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[19].entry.input_buf[2].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[19].entry.input_buf[2].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[19].entry.input_buf[2].genblk1[0].mid ));
 sky130_fd_sc_hd__inv_2 \l_fifo.genblk1[19].entry.input_buf[2].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[19].entry.input_buf[2].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[19].entry.input_buf[2].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[19].entry.input_buf[3].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[19].entry.input_buf[3].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[19].entry.input_buf[3].genblk1[0].mid ));
 sky130_fd_sc_hd__inv_2 \l_fifo.genblk1[19].entry.input_buf[3].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[19].entry.input_buf[3].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[19].entry.input_buf[3].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[19].entry.input_buf[4].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[19].entry.input_buf[4].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[19].entry.input_buf[4].genblk1[0].mid ));
 sky130_fd_sc_hd__clkinv_2 \l_fifo.genblk1[19].entry.input_buf[4].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[19].entry.input_buf[4].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[19].entry.input_buf[4].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[19].entry.input_buf[5].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[19].entry.input_buf[5].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[19].entry.input_buf[5].genblk1[0].mid ));
 sky130_fd_sc_hd__inv_2 \l_fifo.genblk1[19].entry.input_buf[5].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[19].entry.input_buf[5].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[19].entry.input_buf[5].X ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[19].entry.latch[0]  (.D(\l_fifo.genblk1[19].entry.input_buf[0].X ),
    .GATE(\l_fifo.genblk1[19].entry.empty ),
    .RESET_B(net39),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[18].entry.input_buf[0].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[19].entry.latch[1]  (.D(\l_fifo.genblk1[19].entry.input_buf[1].X ),
    .GATE(\l_fifo.genblk1[19].entry.empty ),
    .RESET_B(net39),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[18].entry.input_buf[1].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[19].entry.latch[2]  (.D(\l_fifo.genblk1[19].entry.input_buf[2].X ),
    .GATE(\l_fifo.genblk1[19].entry.empty ),
    .RESET_B(net40),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[18].entry.input_buf[2].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[19].entry.latch[3]  (.D(\l_fifo.genblk1[19].entry.input_buf[3].X ),
    .GATE(\l_fifo.genblk1[19].entry.empty ),
    .RESET_B(net46),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[18].entry.input_buf[3].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[19].entry.latch[4]  (.D(\l_fifo.genblk1[19].entry.input_buf[4].X ),
    .GATE(\l_fifo.genblk1[19].entry.empty ),
    .RESET_B(net46),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[18].entry.input_buf[4].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[19].entry.latch[5]  (.D(\l_fifo.genblk1[19].entry.input_buf[5].X ),
    .GATE(\l_fifo.genblk1[19].entry.empty ),
    .RESET_B(net35),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[18].entry.input_buf[5].A ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[1].entry.input_buf[0].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[1].entry.input_buf[0].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[1].entry.input_buf[0].genblk1[0].mid ));
 sky130_fd_sc_hd__inv_2 \l_fifo.genblk1[1].entry.input_buf[0].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[1].entry.input_buf[0].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[1].entry.input_buf[0].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[1].entry.input_buf[1].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[1].entry.input_buf[1].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[1].entry.input_buf[1].genblk1[0].mid ));
 sky130_fd_sc_hd__inv_2 \l_fifo.genblk1[1].entry.input_buf[1].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[1].entry.input_buf[1].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[1].entry.input_buf[1].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[1].entry.input_buf[2].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[1].entry.input_buf[2].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[1].entry.input_buf[2].genblk1[0].mid ));
 sky130_fd_sc_hd__inv_2 \l_fifo.genblk1[1].entry.input_buf[2].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[1].entry.input_buf[2].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[1].entry.input_buf[2].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[1].entry.input_buf[3].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[1].entry.input_buf[3].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[1].entry.input_buf[3].genblk1[0].mid ));
 sky130_fd_sc_hd__clkinv_2 \l_fifo.genblk1[1].entry.input_buf[3].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[1].entry.input_buf[3].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[1].entry.input_buf[3].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[1].entry.input_buf[4].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[1].entry.input_buf[4].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[1].entry.input_buf[4].genblk1[0].mid ));
 sky130_fd_sc_hd__inv_2 \l_fifo.genblk1[1].entry.input_buf[4].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[1].entry.input_buf[4].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[1].entry.input_buf[4].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[1].entry.input_buf[5].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[1].entry.input_buf[5].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[1].entry.input_buf[5].genblk1[0].mid ));
 sky130_fd_sc_hd__inv_2 \l_fifo.genblk1[1].entry.input_buf[5].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[1].entry.input_buf[5].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[1].entry.input_buf[5].X ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[1].entry.latch[0]  (.D(\l_fifo.genblk1[1].entry.input_buf[0].X ),
    .GATE(\l_fifo.genblk1[1].entry.empty ),
    .RESET_B(net27),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[0].entry.input_buf[0].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[1].entry.latch[1]  (.D(\l_fifo.genblk1[1].entry.input_buf[1].X ),
    .GATE(\l_fifo.genblk1[1].entry.empty ),
    .RESET_B(net23),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[0].entry.input_buf[1].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[1].entry.latch[2]  (.D(\l_fifo.genblk1[1].entry.input_buf[2].X ),
    .GATE(\l_fifo.genblk1[1].entry.empty ),
    .RESET_B(net28),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[0].entry.input_buf[2].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[1].entry.latch[3]  (.D(\l_fifo.genblk1[1].entry.input_buf[3].X ),
    .GATE(\l_fifo.genblk1[1].entry.empty ),
    .RESET_B(net28),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[0].entry.input_buf[3].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[1].entry.latch[4]  (.D(\l_fifo.genblk1[1].entry.input_buf[4].X ),
    .GATE(\l_fifo.genblk1[1].entry.empty ),
    .RESET_B(net28),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[0].entry.input_buf[4].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[1].entry.latch[5]  (.D(\l_fifo.genblk1[1].entry.input_buf[5].X ),
    .GATE(\l_fifo.genblk1[1].entry.empty ),
    .RESET_B(net27),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[0].entry.input_buf[5].A ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[20].entry.input_buf[0].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[20].entry.input_buf[0].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[20].entry.input_buf[0].genblk1[0].mid ));
 sky130_fd_sc_hd__clkinv_2 \l_fifo.genblk1[20].entry.input_buf[0].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[20].entry.input_buf[0].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[20].entry.input_buf[0].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[20].entry.input_buf[1].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[20].entry.input_buf[1].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[20].entry.input_buf[1].genblk1[0].mid ));
 sky130_fd_sc_hd__clkinv_2 \l_fifo.genblk1[20].entry.input_buf[1].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[20].entry.input_buf[1].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[20].entry.input_buf[1].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[20].entry.input_buf[2].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[20].entry.input_buf[2].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[20].entry.input_buf[2].genblk1[0].mid ));
 sky130_fd_sc_hd__inv_2 \l_fifo.genblk1[20].entry.input_buf[2].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[20].entry.input_buf[2].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[20].entry.input_buf[2].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[20].entry.input_buf[3].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[20].entry.input_buf[3].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[20].entry.input_buf[3].genblk1[0].mid ));
 sky130_fd_sc_hd__inv_2 \l_fifo.genblk1[20].entry.input_buf[3].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[20].entry.input_buf[3].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[20].entry.input_buf[3].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[20].entry.input_buf[4].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[20].entry.input_buf[4].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[20].entry.input_buf[4].genblk1[0].mid ));
 sky130_fd_sc_hd__clkinv_2 \l_fifo.genblk1[20].entry.input_buf[4].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[20].entry.input_buf[4].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[20].entry.input_buf[4].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[20].entry.input_buf[5].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[20].entry.input_buf[5].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[20].entry.input_buf[5].genblk1[0].mid ));
 sky130_fd_sc_hd__clkinv_2 \l_fifo.genblk1[20].entry.input_buf[5].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[20].entry.input_buf[5].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[20].entry.input_buf[5].X ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[20].entry.latch[0]  (.D(\l_fifo.genblk1[20].entry.input_buf[0].X ),
    .GATE(\l_fifo.genblk1[20].entry.empty ),
    .RESET_B(net35),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[19].entry.input_buf[0].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[20].entry.latch[1]  (.D(\l_fifo.genblk1[20].entry.input_buf[1].X ),
    .GATE(\l_fifo.genblk1[20].entry.empty ),
    .RESET_B(net39),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[19].entry.input_buf[1].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[20].entry.latch[2]  (.D(\l_fifo.genblk1[20].entry.input_buf[2].X ),
    .GATE(\l_fifo.genblk1[20].entry.empty ),
    .RESET_B(net48),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[19].entry.input_buf[2].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[20].entry.latch[3]  (.D(\l_fifo.genblk1[20].entry.input_buf[3].X ),
    .GATE(\l_fifo.genblk1[20].entry.empty ),
    .RESET_B(net35),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[19].entry.input_buf[3].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[20].entry.latch[4]  (.D(\l_fifo.genblk1[20].entry.input_buf[4].X ),
    .GATE(\l_fifo.genblk1[20].entry.empty ),
    .RESET_B(net39),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[19].entry.input_buf[4].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[20].entry.latch[5]  (.D(\l_fifo.genblk1[20].entry.input_buf[5].X ),
    .GATE(\l_fifo.genblk1[20].entry.empty ),
    .RESET_B(net40),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[19].entry.input_buf[5].A ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[21].entry.input_buf[0].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[21].entry.input_buf[0].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[21].entry.input_buf[0].genblk1[0].mid ));
 sky130_fd_sc_hd__inv_2 \l_fifo.genblk1[21].entry.input_buf[0].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[21].entry.input_buf[0].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[21].entry.input_buf[0].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[21].entry.input_buf[1].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[21].entry.input_buf[1].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[21].entry.input_buf[1].genblk1[0].mid ));
 sky130_fd_sc_hd__inv_2 \l_fifo.genblk1[21].entry.input_buf[1].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[21].entry.input_buf[1].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[21].entry.input_buf[1].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[21].entry.input_buf[2].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[21].entry.input_buf[2].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[21].entry.input_buf[2].genblk1[0].mid ));
 sky130_fd_sc_hd__inv_2 \l_fifo.genblk1[21].entry.input_buf[2].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[21].entry.input_buf[2].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[21].entry.input_buf[2].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[21].entry.input_buf[3].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[21].entry.input_buf[3].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[21].entry.input_buf[3].genblk1[0].mid ));
 sky130_fd_sc_hd__clkinv_2 \l_fifo.genblk1[21].entry.input_buf[3].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[21].entry.input_buf[3].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[21].entry.input_buf[3].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[21].entry.input_buf[4].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[21].entry.input_buf[4].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[21].entry.input_buf[4].genblk1[0].mid ));
 sky130_fd_sc_hd__clkinv_2 \l_fifo.genblk1[21].entry.input_buf[4].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[21].entry.input_buf[4].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[21].entry.input_buf[4].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[21].entry.input_buf[5].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[21].entry.input_buf[5].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[21].entry.input_buf[5].genblk1[0].mid ));
 sky130_fd_sc_hd__clkinv_2 \l_fifo.genblk1[21].entry.input_buf[5].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[21].entry.input_buf[5].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[21].entry.input_buf[5].X ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[21].entry.latch[0]  (.D(\l_fifo.genblk1[21].entry.input_buf[0].X ),
    .GATE(\l_fifo.genblk1[21].entry.empty ),
    .RESET_B(net35),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[20].entry.input_buf[0].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[21].entry.latch[1]  (.D(\l_fifo.genblk1[21].entry.input_buf[1].X ),
    .GATE(\l_fifo.genblk1[21].entry.empty ),
    .RESET_B(net37),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[20].entry.input_buf[1].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[21].entry.latch[2]  (.D(\l_fifo.genblk1[21].entry.input_buf[2].X ),
    .GATE(\l_fifo.genblk1[21].entry.empty ),
    .RESET_B(net40),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[20].entry.input_buf[2].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[21].entry.latch[3]  (.D(\l_fifo.genblk1[21].entry.input_buf[3].X ),
    .GATE(\l_fifo.genblk1[21].entry.empty ),
    .RESET_B(net35),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[20].entry.input_buf[3].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[21].entry.latch[4]  (.D(\l_fifo.genblk1[21].entry.input_buf[4].X ),
    .GATE(\l_fifo.genblk1[21].entry.empty ),
    .RESET_B(net38),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[20].entry.input_buf[4].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[21].entry.latch[5]  (.D(\l_fifo.genblk1[21].entry.input_buf[5].X ),
    .GATE(\l_fifo.genblk1[21].entry.empty ),
    .RESET_B(net40),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[20].entry.input_buf[5].A ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[22].entry.input_buf[0].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[22].entry.input_buf[0].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[22].entry.input_buf[0].genblk1[0].mid ));
 sky130_fd_sc_hd__inv_2 \l_fifo.genblk1[22].entry.input_buf[0].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[22].entry.input_buf[0].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[22].entry.input_buf[0].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[22].entry.input_buf[1].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[22].entry.input_buf[1].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[22].entry.input_buf[1].genblk1[0].mid ));
 sky130_fd_sc_hd__inv_2 \l_fifo.genblk1[22].entry.input_buf[1].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[22].entry.input_buf[1].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[22].entry.input_buf[1].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[22].entry.input_buf[2].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[22].entry.input_buf[2].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[22].entry.input_buf[2].genblk1[0].mid ));
 sky130_fd_sc_hd__clkinv_2 \l_fifo.genblk1[22].entry.input_buf[2].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[22].entry.input_buf[2].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[22].entry.input_buf[2].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[22].entry.input_buf[3].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[22].entry.input_buf[3].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[22].entry.input_buf[3].genblk1[0].mid ));
 sky130_fd_sc_hd__inv_2 \l_fifo.genblk1[22].entry.input_buf[3].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[22].entry.input_buf[3].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[22].entry.input_buf[3].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[22].entry.input_buf[4].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[22].entry.input_buf[4].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[22].entry.input_buf[4].genblk1[0].mid ));
 sky130_fd_sc_hd__clkinv_2 \l_fifo.genblk1[22].entry.input_buf[4].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[22].entry.input_buf[4].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[22].entry.input_buf[4].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[22].entry.input_buf[5].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[22].entry.input_buf[5].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[22].entry.input_buf[5].genblk1[0].mid ));
 sky130_fd_sc_hd__inv_2 \l_fifo.genblk1[22].entry.input_buf[5].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[22].entry.input_buf[5].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[22].entry.input_buf[5].X ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[22].entry.latch[0]  (.D(\l_fifo.genblk1[22].entry.input_buf[0].X ),
    .GATE(\l_fifo.genblk1[22].entry.empty ),
    .RESET_B(net37),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[21].entry.input_buf[0].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[22].entry.latch[1]  (.D(\l_fifo.genblk1[22].entry.input_buf[1].X ),
    .GATE(\l_fifo.genblk1[22].entry.empty ),
    .RESET_B(net38),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[21].entry.input_buf[1].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[22].entry.latch[2]  (.D(\l_fifo.genblk1[22].entry.input_buf[2].X ),
    .GATE(\l_fifo.genblk1[22].entry.empty ),
    .RESET_B(net40),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[21].entry.input_buf[2].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[22].entry.latch[3]  (.D(\l_fifo.genblk1[22].entry.input_buf[3].X ),
    .GATE(\l_fifo.genblk1[22].entry.empty ),
    .RESET_B(net14),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[21].entry.input_buf[3].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[22].entry.latch[4]  (.D(\l_fifo.genblk1[22].entry.input_buf[4].X ),
    .GATE(\l_fifo.genblk1[22].entry.empty ),
    .RESET_B(net37),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[21].entry.input_buf[4].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[22].entry.latch[5]  (.D(\l_fifo.genblk1[22].entry.input_buf[5].X ),
    .GATE(\l_fifo.genblk1[22].entry.empty ),
    .RESET_B(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[21].entry.input_buf[5].A ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[23].entry.input_buf[0].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[23].entry.input_buf[0].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[23].entry.input_buf[0].genblk1[0].mid ));
 sky130_fd_sc_hd__clkinv_2 \l_fifo.genblk1[23].entry.input_buf[0].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[23].entry.input_buf[0].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[23].entry.input_buf[0].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[23].entry.input_buf[1].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[23].entry.input_buf[1].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[23].entry.input_buf[1].genblk1[0].mid ));
 sky130_fd_sc_hd__clkinv_2 \l_fifo.genblk1[23].entry.input_buf[1].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[23].entry.input_buf[1].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[23].entry.input_buf[1].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[23].entry.input_buf[2].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[23].entry.input_buf[2].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[23].entry.input_buf[2].genblk1[0].mid ));
 sky130_fd_sc_hd__inv_2 \l_fifo.genblk1[23].entry.input_buf[2].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[23].entry.input_buf[2].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[23].entry.input_buf[2].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[23].entry.input_buf[3].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[23].entry.input_buf[3].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[23].entry.input_buf[3].genblk1[0].mid ));
 sky130_fd_sc_hd__inv_2 \l_fifo.genblk1[23].entry.input_buf[3].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[23].entry.input_buf[3].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[23].entry.input_buf[3].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[23].entry.input_buf[4].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[23].entry.input_buf[4].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[23].entry.input_buf[4].genblk1[0].mid ));
 sky130_fd_sc_hd__inv_2 \l_fifo.genblk1[23].entry.input_buf[4].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[23].entry.input_buf[4].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[23].entry.input_buf[4].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[23].entry.input_buf[5].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[23].entry.input_buf[5].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[23].entry.input_buf[5].genblk1[0].mid ));
 sky130_fd_sc_hd__inv_2 \l_fifo.genblk1[23].entry.input_buf[5].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[23].entry.input_buf[5].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[23].entry.input_buf[5].X ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[23].entry.latch[0]  (.D(\l_fifo.genblk1[23].entry.input_buf[0].X ),
    .GATE(\l_fifo.genblk1[23].entry.empty ),
    .RESET_B(net37),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[22].entry.input_buf[0].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[23].entry.latch[1]  (.D(\l_fifo.genblk1[23].entry.input_buf[1].X ),
    .GATE(\l_fifo.genblk1[23].entry.empty ),
    .RESET_B(net37),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[22].entry.input_buf[1].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[23].entry.latch[2]  (.D(\l_fifo.genblk1[23].entry.input_buf[2].X ),
    .GATE(\l_fifo.genblk1[23].entry.empty ),
    .RESET_B(net39),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[22].entry.input_buf[2].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[23].entry.latch[3]  (.D(\l_fifo.genblk1[23].entry.input_buf[3].X ),
    .GATE(\l_fifo.genblk1[23].entry.empty ),
    .RESET_B(net38),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[22].entry.input_buf[3].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[23].entry.latch[4]  (.D(\l_fifo.genblk1[23].entry.input_buf[4].X ),
    .GATE(\l_fifo.genblk1[23].entry.empty ),
    .RESET_B(net39),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[22].entry.input_buf[4].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[23].entry.latch[5]  (.D(\l_fifo.genblk1[23].entry.input_buf[5].X ),
    .GATE(\l_fifo.genblk1[23].entry.empty ),
    .RESET_B(net34),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[22].entry.input_buf[5].A ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[24].entry.input_buf[0].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[24].entry.input_buf[0].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[24].entry.input_buf[0].genblk1[0].mid ));
 sky130_fd_sc_hd__clkinv_2 \l_fifo.genblk1[24].entry.input_buf[0].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[24].entry.input_buf[0].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[24].entry.input_buf[0].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[24].entry.input_buf[1].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[24].entry.input_buf[1].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[24].entry.input_buf[1].genblk1[0].mid ));
 sky130_fd_sc_hd__clkinv_2 \l_fifo.genblk1[24].entry.input_buf[1].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[24].entry.input_buf[1].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[24].entry.input_buf[1].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[24].entry.input_buf[2].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[24].entry.input_buf[2].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[24].entry.input_buf[2].genblk1[0].mid ));
 sky130_fd_sc_hd__clkinv_2 \l_fifo.genblk1[24].entry.input_buf[2].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[24].entry.input_buf[2].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[24].entry.input_buf[2].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[24].entry.input_buf[3].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[24].entry.input_buf[3].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[24].entry.input_buf[3].genblk1[0].mid ));
 sky130_fd_sc_hd__clkinv_2 \l_fifo.genblk1[24].entry.input_buf[3].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[24].entry.input_buf[3].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[24].entry.input_buf[3].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[24].entry.input_buf[4].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[24].entry.input_buf[4].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[24].entry.input_buf[4].genblk1[0].mid ));
 sky130_fd_sc_hd__clkinv_2 \l_fifo.genblk1[24].entry.input_buf[4].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[24].entry.input_buf[4].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[24].entry.input_buf[4].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[24].entry.input_buf[5].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[24].entry.input_buf[5].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[24].entry.input_buf[5].genblk1[0].mid ));
 sky130_fd_sc_hd__inv_2 \l_fifo.genblk1[24].entry.input_buf[5].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[24].entry.input_buf[5].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[24].entry.input_buf[5].X ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[24].entry.latch[0]  (.D(\l_fifo.genblk1[24].entry.input_buf[0].X ),
    .GATE(\l_fifo.genblk1[24].entry.empty ),
    .RESET_B(net38),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[23].entry.input_buf[0].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[24].entry.latch[1]  (.D(\l_fifo.genblk1[24].entry.input_buf[1].X ),
    .GATE(\l_fifo.genblk1[24].entry.empty ),
    .RESET_B(net19),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[23].entry.input_buf[1].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[24].entry.latch[2]  (.D(\l_fifo.genblk1[24].entry.input_buf[2].X ),
    .GATE(\l_fifo.genblk1[24].entry.empty ),
    .RESET_B(net18),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[23].entry.input_buf[2].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[24].entry.latch[3]  (.D(\l_fifo.genblk1[24].entry.input_buf[3].X ),
    .GATE(\l_fifo.genblk1[24].entry.empty ),
    .RESET_B(net38),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[23].entry.input_buf[3].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[24].entry.latch[4]  (.D(\l_fifo.genblk1[24].entry.input_buf[4].X ),
    .GATE(\l_fifo.genblk1[24].entry.empty ),
    .RESET_B(net37),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[23].entry.input_buf[4].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[24].entry.latch[5]  (.D(\l_fifo.genblk1[24].entry.input_buf[5].X ),
    .GATE(\l_fifo.genblk1[24].entry.empty ),
    .RESET_B(net37),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[23].entry.input_buf[5].A ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[25].entry.input_buf[0].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[25].entry.input_buf[0].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[25].entry.input_buf[0].genblk1[0].mid ));
 sky130_fd_sc_hd__inv_2 \l_fifo.genblk1[25].entry.input_buf[0].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[25].entry.input_buf[0].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[25].entry.input_buf[0].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[25].entry.input_buf[1].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[25].entry.input_buf[1].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[25].entry.input_buf[1].genblk1[0].mid ));
 sky130_fd_sc_hd__inv_2 \l_fifo.genblk1[25].entry.input_buf[1].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[25].entry.input_buf[1].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[25].entry.input_buf[1].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[25].entry.input_buf[2].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[25].entry.input_buf[2].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[25].entry.input_buf[2].genblk1[0].mid ));
 sky130_fd_sc_hd__inv_2 \l_fifo.genblk1[25].entry.input_buf[2].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[25].entry.input_buf[2].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[25].entry.input_buf[2].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[25].entry.input_buf[3].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[25].entry.input_buf[3].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[25].entry.input_buf[3].genblk1[0].mid ));
 sky130_fd_sc_hd__clkinv_2 \l_fifo.genblk1[25].entry.input_buf[3].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[25].entry.input_buf[3].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[25].entry.input_buf[3].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[25].entry.input_buf[4].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[25].entry.input_buf[4].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[25].entry.input_buf[4].genblk1[0].mid ));
 sky130_fd_sc_hd__clkinv_2 \l_fifo.genblk1[25].entry.input_buf[4].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[25].entry.input_buf[4].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[25].entry.input_buf[4].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[25].entry.input_buf[5].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[25].entry.input_buf[5].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[25].entry.input_buf[5].genblk1[0].mid ));
 sky130_fd_sc_hd__clkinv_2 \l_fifo.genblk1[25].entry.input_buf[5].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[25].entry.input_buf[5].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[25].entry.input_buf[5].X ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[25].entry.latch[0]  (.D(\l_fifo.genblk1[25].entry.input_buf[0].X ),
    .GATE(\l_fifo.genblk1[25].entry.empty ),
    .RESET_B(net37),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[24].entry.input_buf[0].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[25].entry.latch[1]  (.D(\l_fifo.genblk1[25].entry.input_buf[1].X ),
    .GATE(\l_fifo.genblk1[25].entry.empty ),
    .RESET_B(net19),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[24].entry.input_buf[1].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[25].entry.latch[2]  (.D(\l_fifo.genblk1[25].entry.input_buf[2].X ),
    .GATE(\l_fifo.genblk1[25].entry.empty ),
    .RESET_B(net18),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[24].entry.input_buf[2].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[25].entry.latch[3]  (.D(\l_fifo.genblk1[25].entry.input_buf[3].X ),
    .GATE(\l_fifo.genblk1[25].entry.empty ),
    .RESET_B(net37),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[24].entry.input_buf[3].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[25].entry.latch[4]  (.D(\l_fifo.genblk1[25].entry.input_buf[4].X ),
    .GATE(\l_fifo.genblk1[25].entry.empty ),
    .RESET_B(net18),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[24].entry.input_buf[4].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[25].entry.latch[5]  (.D(\l_fifo.genblk1[25].entry.input_buf[5].X ),
    .GATE(\l_fifo.genblk1[25].entry.empty ),
    .RESET_B(net18),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[24].entry.input_buf[5].A ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[26].entry.input_buf[0].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[26].entry.input_buf[0].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[26].entry.input_buf[0].genblk1[0].mid ));
 sky130_fd_sc_hd__inv_2 \l_fifo.genblk1[26].entry.input_buf[0].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[26].entry.input_buf[0].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[26].entry.input_buf[0].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[26].entry.input_buf[1].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[26].entry.input_buf[1].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[26].entry.input_buf[1].genblk1[0].mid ));
 sky130_fd_sc_hd__clkinv_2 \l_fifo.genblk1[26].entry.input_buf[1].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[26].entry.input_buf[1].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[26].entry.input_buf[1].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[26].entry.input_buf[2].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[26].entry.input_buf[2].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[26].entry.input_buf[2].genblk1[0].mid ));
 sky130_fd_sc_hd__clkinv_2 \l_fifo.genblk1[26].entry.input_buf[2].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[26].entry.input_buf[2].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[26].entry.input_buf[2].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[26].entry.input_buf[3].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[26].entry.input_buf[3].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[26].entry.input_buf[3].genblk1[0].mid ));
 sky130_fd_sc_hd__clkinv_2 \l_fifo.genblk1[26].entry.input_buf[3].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[26].entry.input_buf[3].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[26].entry.input_buf[3].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[26].entry.input_buf[4].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[26].entry.input_buf[4].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[26].entry.input_buf[4].genblk1[0].mid ));
 sky130_fd_sc_hd__inv_2 \l_fifo.genblk1[26].entry.input_buf[4].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[26].entry.input_buf[4].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[26].entry.input_buf[4].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[26].entry.input_buf[5].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[26].entry.input_buf[5].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[26].entry.input_buf[5].genblk1[0].mid ));
 sky130_fd_sc_hd__inv_2 \l_fifo.genblk1[26].entry.input_buf[5].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[26].entry.input_buf[5].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[26].entry.input_buf[5].X ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[26].entry.latch[0]  (.D(\l_fifo.genblk1[26].entry.input_buf[0].X ),
    .GATE(\l_fifo.genblk1[26].entry.empty ),
    .RESET_B(net18),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[25].entry.input_buf[0].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[26].entry.latch[1]  (.D(\l_fifo.genblk1[26].entry.input_buf[1].X ),
    .GATE(\l_fifo.genblk1[26].entry.empty ),
    .RESET_B(net19),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[25].entry.input_buf[1].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[26].entry.latch[2]  (.D(\l_fifo.genblk1[26].entry.input_buf[2].X ),
    .GATE(\l_fifo.genblk1[26].entry.empty ),
    .RESET_B(net14),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[25].entry.input_buf[2].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[26].entry.latch[3]  (.D(\l_fifo.genblk1[26].entry.input_buf[3].X ),
    .GATE(\l_fifo.genblk1[26].entry.empty ),
    .RESET_B(net13),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[25].entry.input_buf[3].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[26].entry.latch[4]  (.D(\l_fifo.genblk1[26].entry.input_buf[4].X ),
    .GATE(\l_fifo.genblk1[26].entry.empty ),
    .RESET_B(net18),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[25].entry.input_buf[4].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[26].entry.latch[5]  (.D(\l_fifo.genblk1[26].entry.input_buf[5].X ),
    .GATE(\l_fifo.genblk1[26].entry.empty ),
    .RESET_B(net15),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[25].entry.input_buf[5].A ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[27].entry.input_buf[0].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[27].entry.input_buf[0].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[27].entry.input_buf[0].genblk1[0].mid ));
 sky130_fd_sc_hd__inv_2 \l_fifo.genblk1[27].entry.input_buf[0].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[27].entry.input_buf[0].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[27].entry.input_buf[0].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[27].entry.input_buf[1].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[27].entry.input_buf[1].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[27].entry.input_buf[1].genblk1[0].mid ));
 sky130_fd_sc_hd__inv_2 \l_fifo.genblk1[27].entry.input_buf[1].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[27].entry.input_buf[1].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[27].entry.input_buf[1].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[27].entry.input_buf[2].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[27].entry.input_buf[2].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[27].entry.input_buf[2].genblk1[0].mid ));
 sky130_fd_sc_hd__inv_2 \l_fifo.genblk1[27].entry.input_buf[2].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[27].entry.input_buf[2].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[27].entry.input_buf[2].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[27].entry.input_buf[3].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[27].entry.input_buf[3].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[27].entry.input_buf[3].genblk1[0].mid ));
 sky130_fd_sc_hd__clkinv_2 \l_fifo.genblk1[27].entry.input_buf[3].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[27].entry.input_buf[3].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[27].entry.input_buf[3].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[27].entry.input_buf[4].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[27].entry.input_buf[4].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[27].entry.input_buf[4].genblk1[0].mid ));
 sky130_fd_sc_hd__inv_2 \l_fifo.genblk1[27].entry.input_buf[4].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[27].entry.input_buf[4].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[27].entry.input_buf[4].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[27].entry.input_buf[5].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[27].entry.input_buf[5].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[27].entry.input_buf[5].genblk1[0].mid ));
 sky130_fd_sc_hd__inv_2 \l_fifo.genblk1[27].entry.input_buf[5].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[27].entry.input_buf[5].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[27].entry.input_buf[5].X ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[27].entry.latch[0]  (.D(\l_fifo.genblk1[27].entry.input_buf[0].X ),
    .GATE(\l_fifo.genblk1[27].entry.empty ),
    .RESET_B(net19),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[26].entry.input_buf[0].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[27].entry.latch[1]  (.D(\l_fifo.genblk1[27].entry.input_buf[1].X ),
    .GATE(\l_fifo.genblk1[27].entry.empty ),
    .RESET_B(net18),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[26].entry.input_buf[1].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[27].entry.latch[2]  (.D(\l_fifo.genblk1[27].entry.input_buf[2].X ),
    .GATE(\l_fifo.genblk1[27].entry.empty ),
    .RESET_B(net16),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[26].entry.input_buf[2].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[27].entry.latch[3]  (.D(\l_fifo.genblk1[27].entry.input_buf[3].X ),
    .GATE(\l_fifo.genblk1[27].entry.empty ),
    .RESET_B(net18),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[26].entry.input_buf[3].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[27].entry.latch[4]  (.D(\l_fifo.genblk1[27].entry.input_buf[4].X ),
    .GATE(\l_fifo.genblk1[27].entry.empty ),
    .RESET_B(net19),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[26].entry.input_buf[4].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[27].entry.latch[5]  (.D(\l_fifo.genblk1[27].entry.input_buf[5].X ),
    .GATE(\l_fifo.genblk1[27].entry.empty ),
    .RESET_B(net37),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[26].entry.input_buf[5].A ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[28].entry.input_buf[0].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[28].entry.input_buf[0].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[28].entry.input_buf[0].genblk1[0].mid ));
 sky130_fd_sc_hd__clkinv_2 \l_fifo.genblk1[28].entry.input_buf[0].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[28].entry.input_buf[0].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[28].entry.input_buf[0].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[28].entry.input_buf[1].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[28].entry.input_buf[1].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[28].entry.input_buf[1].genblk1[0].mid ));
 sky130_fd_sc_hd__clkinv_2 \l_fifo.genblk1[28].entry.input_buf[1].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[28].entry.input_buf[1].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[28].entry.input_buf[1].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[28].entry.input_buf[2].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[28].entry.input_buf[2].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[28].entry.input_buf[2].genblk1[0].mid ));
 sky130_fd_sc_hd__inv_2 \l_fifo.genblk1[28].entry.input_buf[2].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[28].entry.input_buf[2].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[28].entry.input_buf[2].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[28].entry.input_buf[3].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[28].entry.input_buf[3].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[28].entry.input_buf[3].genblk1[0].mid ));
 sky130_fd_sc_hd__clkinv_2 \l_fifo.genblk1[28].entry.input_buf[3].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[28].entry.input_buf[3].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[28].entry.input_buf[3].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[28].entry.input_buf[4].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[28].entry.input_buf[4].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[28].entry.input_buf[4].genblk1[0].mid ));
 sky130_fd_sc_hd__clkinv_2 \l_fifo.genblk1[28].entry.input_buf[4].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[28].entry.input_buf[4].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[28].entry.input_buf[4].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[28].entry.input_buf[5].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[28].entry.input_buf[5].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[28].entry.input_buf[5].genblk1[0].mid ));
 sky130_fd_sc_hd__clkinv_2 \l_fifo.genblk1[28].entry.input_buf[5].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[28].entry.input_buf[5].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[28].entry.input_buf[5].X ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[28].entry.latch[0]  (.D(\l_fifo.genblk1[28].entry.input_buf[0].X ),
    .GATE(\l_fifo.genblk1[28].entry.empty ),
    .RESET_B(net17),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[27].entry.input_buf[0].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[28].entry.latch[1]  (.D(\l_fifo.genblk1[28].entry.input_buf[1].X ),
    .GATE(\l_fifo.genblk1[28].entry.empty ),
    .RESET_B(net20),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[27].entry.input_buf[1].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[28].entry.latch[2]  (.D(\l_fifo.genblk1[28].entry.input_buf[2].X ),
    .GATE(\l_fifo.genblk1[28].entry.empty ),
    .RESET_B(net19),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[27].entry.input_buf[2].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[28].entry.latch[3]  (.D(\l_fifo.genblk1[28].entry.input_buf[3].X ),
    .GATE(\l_fifo.genblk1[28].entry.empty ),
    .RESET_B(net18),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[27].entry.input_buf[3].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[28].entry.latch[4]  (.D(\l_fifo.genblk1[28].entry.input_buf[4].X ),
    .GATE(\l_fifo.genblk1[28].entry.empty ),
    .RESET_B(net17),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[27].entry.input_buf[4].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[28].entry.latch[5]  (.D(\l_fifo.genblk1[28].entry.input_buf[5].X ),
    .GATE(\l_fifo.genblk1[28].entry.empty ),
    .RESET_B(net18),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[27].entry.input_buf[5].A ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[29].entry.input_buf[0].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[29].entry.input_buf[0].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[29].entry.input_buf[0].genblk1[0].mid ));
 sky130_fd_sc_hd__inv_2 \l_fifo.genblk1[29].entry.input_buf[0].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[29].entry.input_buf[0].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[29].entry.input_buf[0].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[29].entry.input_buf[1].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[29].entry.input_buf[1].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[29].entry.input_buf[1].genblk1[0].mid ));
 sky130_fd_sc_hd__inv_2 \l_fifo.genblk1[29].entry.input_buf[1].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[29].entry.input_buf[1].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[29].entry.input_buf[1].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[29].entry.input_buf[2].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[29].entry.input_buf[2].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[29].entry.input_buf[2].genblk1[0].mid ));
 sky130_fd_sc_hd__clkinv_2 \l_fifo.genblk1[29].entry.input_buf[2].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[29].entry.input_buf[2].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[29].entry.input_buf[2].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[29].entry.input_buf[3].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[29].entry.input_buf[3].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[29].entry.input_buf[3].genblk1[0].mid ));
 sky130_fd_sc_hd__clkinv_2 \l_fifo.genblk1[29].entry.input_buf[3].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[29].entry.input_buf[3].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[29].entry.input_buf[3].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[29].entry.input_buf[4].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[29].entry.input_buf[4].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[29].entry.input_buf[4].genblk1[0].mid ));
 sky130_fd_sc_hd__inv_2 \l_fifo.genblk1[29].entry.input_buf[4].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[29].entry.input_buf[4].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[29].entry.input_buf[4].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[29].entry.input_buf[5].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[29].entry.input_buf[5].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[29].entry.input_buf[5].genblk1[0].mid ));
 sky130_fd_sc_hd__inv_2 \l_fifo.genblk1[29].entry.input_buf[5].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[29].entry.input_buf[5].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[29].entry.input_buf[5].X ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[29].entry.latch[0]  (.D(\l_fifo.genblk1[29].entry.input_buf[0].X ),
    .GATE(\l_fifo.genblk1[29].entry.empty ),
    .RESET_B(net12),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[28].entry.input_buf[0].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[29].entry.latch[1]  (.D(\l_fifo.genblk1[29].entry.input_buf[1].X ),
    .GATE(\l_fifo.genblk1[29].entry.empty ),
    .RESET_B(net17),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[28].entry.input_buf[1].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[29].entry.latch[2]  (.D(\l_fifo.genblk1[29].entry.input_buf[2].X ),
    .GATE(\l_fifo.genblk1[29].entry.empty ),
    .RESET_B(net17),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[28].entry.input_buf[2].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[29].entry.latch[3]  (.D(\l_fifo.genblk1[29].entry.input_buf[3].X ),
    .GATE(\l_fifo.genblk1[29].entry.empty ),
    .RESET_B(net17),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[28].entry.input_buf[3].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[29].entry.latch[4]  (.D(\l_fifo.genblk1[29].entry.input_buf[4].X ),
    .GATE(\l_fifo.genblk1[29].entry.empty ),
    .RESET_B(net13),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[28].entry.input_buf[4].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[29].entry.latch[5]  (.D(\l_fifo.genblk1[29].entry.input_buf[5].X ),
    .GATE(\l_fifo.genblk1[29].entry.empty ),
    .RESET_B(net17),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[28].entry.input_buf[5].A ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[2].entry.input_buf[0].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[2].entry.input_buf[0].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[2].entry.input_buf[0].genblk1[0].mid ));
 sky130_fd_sc_hd__inv_2 \l_fifo.genblk1[2].entry.input_buf[0].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[2].entry.input_buf[0].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[2].entry.input_buf[0].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[2].entry.input_buf[1].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[2].entry.input_buf[1].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[2].entry.input_buf[1].genblk1[0].mid ));
 sky130_fd_sc_hd__clkinv_2 \l_fifo.genblk1[2].entry.input_buf[1].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[2].entry.input_buf[1].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[2].entry.input_buf[1].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[2].entry.input_buf[2].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[2].entry.input_buf[2].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[2].entry.input_buf[2].genblk1[0].mid ));
 sky130_fd_sc_hd__clkinv_2 \l_fifo.genblk1[2].entry.input_buf[2].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[2].entry.input_buf[2].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[2].entry.input_buf[2].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[2].entry.input_buf[3].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[2].entry.input_buf[3].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[2].entry.input_buf[3].genblk1[0].mid ));
 sky130_fd_sc_hd__inv_2 \l_fifo.genblk1[2].entry.input_buf[3].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[2].entry.input_buf[3].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[2].entry.input_buf[3].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[2].entry.input_buf[4].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[2].entry.input_buf[4].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[2].entry.input_buf[4].genblk1[0].mid ));
 sky130_fd_sc_hd__inv_2 \l_fifo.genblk1[2].entry.input_buf[4].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[2].entry.input_buf[4].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[2].entry.input_buf[4].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[2].entry.input_buf[5].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[2].entry.input_buf[5].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[2].entry.input_buf[5].genblk1[0].mid ));
 sky130_fd_sc_hd__clkinv_2 \l_fifo.genblk1[2].entry.input_buf[5].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[2].entry.input_buf[5].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[2].entry.input_buf[5].X ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[2].entry.latch[0]  (.D(\l_fifo.genblk1[2].entry.input_buf[0].X ),
    .GATE(\l_fifo.genblk1[2].entry.empty ),
    .RESET_B(net27),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[1].entry.input_buf[0].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[2].entry.latch[1]  (.D(\l_fifo.genblk1[2].entry.input_buf[1].X ),
    .GATE(\l_fifo.genblk1[2].entry.empty ),
    .RESET_B(net27),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[1].entry.input_buf[1].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[2].entry.latch[2]  (.D(\l_fifo.genblk1[2].entry.input_buf[2].X ),
    .GATE(\l_fifo.genblk1[2].entry.empty ),
    .RESET_B(net26),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[1].entry.input_buf[2].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[2].entry.latch[3]  (.D(\l_fifo.genblk1[2].entry.input_buf[3].X ),
    .GATE(\l_fifo.genblk1[2].entry.empty ),
    .RESET_B(net26),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[1].entry.input_buf[3].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[2].entry.latch[4]  (.D(\l_fifo.genblk1[2].entry.input_buf[4].X ),
    .GATE(\l_fifo.genblk1[2].entry.empty ),
    .RESET_B(net26),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[1].entry.input_buf[4].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[2].entry.latch[5]  (.D(\l_fifo.genblk1[2].entry.input_buf[5].X ),
    .GATE(\l_fifo.genblk1[2].entry.empty ),
    .RESET_B(net26),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[1].entry.input_buf[5].A ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[30].entry.input_buf[0].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[30].entry.input_buf[0].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[30].entry.input_buf[0].genblk1[0].mid ));
 sky130_fd_sc_hd__clkinv_2 \l_fifo.genblk1[30].entry.input_buf[0].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[30].entry.input_buf[0].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[30].entry.input_buf[0].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[30].entry.input_buf[1].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[30].entry.input_buf[1].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[30].entry.input_buf[1].genblk1[0].mid ));
 sky130_fd_sc_hd__inv_2 \l_fifo.genblk1[30].entry.input_buf[1].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[30].entry.input_buf[1].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[30].entry.input_buf[1].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[30].entry.input_buf[2].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[30].entry.input_buf[2].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[30].entry.input_buf[2].genblk1[0].mid ));
 sky130_fd_sc_hd__inv_2 \l_fifo.genblk1[30].entry.input_buf[2].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[30].entry.input_buf[2].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[30].entry.input_buf[2].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[30].entry.input_buf[3].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[30].entry.input_buf[3].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[30].entry.input_buf[3].genblk1[0].mid ));
 sky130_fd_sc_hd__inv_2 \l_fifo.genblk1[30].entry.input_buf[3].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[30].entry.input_buf[3].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[30].entry.input_buf[3].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[30].entry.input_buf[4].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[30].entry.input_buf[4].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[30].entry.input_buf[4].genblk1[0].mid ));
 sky130_fd_sc_hd__inv_2 \l_fifo.genblk1[30].entry.input_buf[4].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[30].entry.input_buf[4].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[30].entry.input_buf[4].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[30].entry.input_buf[5].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[30].entry.input_buf[5].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[30].entry.input_buf[5].genblk1[0].mid ));
 sky130_fd_sc_hd__inv_2 \l_fifo.genblk1[30].entry.input_buf[5].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[30].entry.input_buf[5].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[30].entry.input_buf[5].X ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[30].entry.latch[0]  (.D(\l_fifo.genblk1[30].entry.input_buf[0].X ),
    .GATE(\l_fifo.genblk1[30].entry.empty ),
    .RESET_B(net12),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[29].entry.input_buf[0].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[30].entry.latch[1]  (.D(\l_fifo.genblk1[30].entry.input_buf[1].X ),
    .GATE(\l_fifo.genblk1[30].entry.empty ),
    .RESET_B(net17),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[29].entry.input_buf[1].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[30].entry.latch[2]  (.D(\l_fifo.genblk1[30].entry.input_buf[2].X ),
    .GATE(\l_fifo.genblk1[30].entry.empty ),
    .RESET_B(net20),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[29].entry.input_buf[2].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[30].entry.latch[3]  (.D(\l_fifo.genblk1[30].entry.input_buf[3].X ),
    .GATE(\l_fifo.genblk1[30].entry.empty ),
    .RESET_B(net9),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[29].entry.input_buf[3].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[30].entry.latch[4]  (.D(\l_fifo.genblk1[30].entry.input_buf[4].X ),
    .GATE(\l_fifo.genblk1[30].entry.empty ),
    .RESET_B(net17),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[29].entry.input_buf[4].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[30].entry.latch[5]  (.D(\l_fifo.genblk1[30].entry.input_buf[5].X ),
    .GATE(\l_fifo.genblk1[30].entry.empty ),
    .RESET_B(net17),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[29].entry.input_buf[5].A ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[31].entry.input_buf[0].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[31].entry.input_buf[0].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[31].entry.input_buf[0].genblk1[0].mid ));
 sky130_fd_sc_hd__inv_2 \l_fifo.genblk1[31].entry.input_buf[0].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[31].entry.input_buf[0].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[31].entry.input_buf[0].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[31].entry.input_buf[1].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[31].entry.input_buf[1].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[31].entry.input_buf[1].genblk1[0].mid ));
 sky130_fd_sc_hd__clkinv_2 \l_fifo.genblk1[31].entry.input_buf[1].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[31].entry.input_buf[1].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[31].entry.input_buf[1].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[31].entry.input_buf[2].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[31].entry.input_buf[2].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[31].entry.input_buf[2].genblk1[0].mid ));
 sky130_fd_sc_hd__clkinv_2 \l_fifo.genblk1[31].entry.input_buf[2].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[31].entry.input_buf[2].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[31].entry.input_buf[2].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[31].entry.input_buf[3].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[31].entry.input_buf[3].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[31].entry.input_buf[3].genblk1[0].mid ));
 sky130_fd_sc_hd__inv_2 \l_fifo.genblk1[31].entry.input_buf[3].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[31].entry.input_buf[3].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[31].entry.input_buf[3].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[31].entry.input_buf[4].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[31].entry.input_buf[4].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[31].entry.input_buf[4].genblk1[0].mid ));
 sky130_fd_sc_hd__inv_2 \l_fifo.genblk1[31].entry.input_buf[4].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[31].entry.input_buf[4].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[31].entry.input_buf[4].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[31].entry.input_buf[5].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[31].entry.input_buf[5].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[31].entry.input_buf[5].genblk1[0].mid ));
 sky130_fd_sc_hd__inv_2 \l_fifo.genblk1[31].entry.input_buf[5].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[31].entry.input_buf[5].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[31].entry.input_buf[5].X ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[31].entry.latch[0]  (.D(\l_fifo.genblk1[31].entry.input_buf[0].X ),
    .GATE(\l_fifo.genblk1[31].entry.empty ),
    .RESET_B(net12),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[30].entry.input_buf[0].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[31].entry.latch[1]  (.D(\l_fifo.genblk1[31].entry.input_buf[1].X ),
    .GATE(\l_fifo.genblk1[31].entry.empty ),
    .RESET_B(net21),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[30].entry.input_buf[1].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[31].entry.latch[2]  (.D(\l_fifo.genblk1[31].entry.input_buf[2].X ),
    .GATE(\l_fifo.genblk1[31].entry.empty ),
    .RESET_B(net12),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[30].entry.input_buf[2].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[31].entry.latch[3]  (.D(\l_fifo.genblk1[31].entry.input_buf[3].X ),
    .GATE(\l_fifo.genblk1[31].entry.empty ),
    .RESET_B(net16),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[30].entry.input_buf[3].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[31].entry.latch[4]  (.D(\l_fifo.genblk1[31].entry.input_buf[4].X ),
    .GATE(\l_fifo.genblk1[31].entry.empty ),
    .RESET_B(net13),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[30].entry.input_buf[4].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[31].entry.latch[5]  (.D(\l_fifo.genblk1[31].entry.input_buf[5].X ),
    .GATE(\l_fifo.genblk1[31].entry.empty ),
    .RESET_B(net17),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[30].entry.input_buf[5].A ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[32].entry.input_buf[0].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[32].entry.input_buf[0].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[32].entry.input_buf[0].genblk1[0].mid ));
 sky130_fd_sc_hd__clkinv_2 \l_fifo.genblk1[32].entry.input_buf[0].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[32].entry.input_buf[0].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[32].entry.input_buf[0].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[32].entry.input_buf[1].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[32].entry.input_buf[1].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[32].entry.input_buf[1].genblk1[0].mid ));
 sky130_fd_sc_hd__inv_2 \l_fifo.genblk1[32].entry.input_buf[1].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[32].entry.input_buf[1].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[32].entry.input_buf[1].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[32].entry.input_buf[2].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[32].entry.input_buf[2].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[32].entry.input_buf[2].genblk1[0].mid ));
 sky130_fd_sc_hd__inv_2 \l_fifo.genblk1[32].entry.input_buf[2].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[32].entry.input_buf[2].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[32].entry.input_buf[2].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[32].entry.input_buf[3].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[32].entry.input_buf[3].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[32].entry.input_buf[3].genblk1[0].mid ));
 sky130_fd_sc_hd__inv_2 \l_fifo.genblk1[32].entry.input_buf[3].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[32].entry.input_buf[3].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[32].entry.input_buf[3].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[32].entry.input_buf[4].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[32].entry.input_buf[4].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[32].entry.input_buf[4].genblk1[0].mid ));
 sky130_fd_sc_hd__inv_2 \l_fifo.genblk1[32].entry.input_buf[4].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[32].entry.input_buf[4].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[32].entry.input_buf[4].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[32].entry.input_buf[5].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[32].entry.input_buf[5].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[32].entry.input_buf[5].genblk1[0].mid ));
 sky130_fd_sc_hd__clkinv_2 \l_fifo.genblk1[32].entry.input_buf[5].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[32].entry.input_buf[5].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[32].entry.input_buf[5].X ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[32].entry.latch[0]  (.D(\l_fifo.genblk1[32].entry.input_buf[0].X ),
    .GATE(\l_fifo.genblk1[32].entry.empty ),
    .RESET_B(net12),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[31].entry.input_buf[0].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[32].entry.latch[1]  (.D(\l_fifo.genblk1[32].entry.input_buf[1].X ),
    .GATE(\l_fifo.genblk1[32].entry.empty ),
    .RESET_B(net10),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[31].entry.input_buf[1].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[32].entry.latch[2]  (.D(\l_fifo.genblk1[32].entry.input_buf[2].X ),
    .GATE(\l_fifo.genblk1[32].entry.empty ),
    .RESET_B(net12),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[31].entry.input_buf[2].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[32].entry.latch[3]  (.D(\l_fifo.genblk1[32].entry.input_buf[3].X ),
    .GATE(\l_fifo.genblk1[32].entry.empty ),
    .RESET_B(net9),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[31].entry.input_buf[3].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[32].entry.latch[4]  (.D(\l_fifo.genblk1[32].entry.input_buf[4].X ),
    .GATE(\l_fifo.genblk1[32].entry.empty ),
    .RESET_B(net9),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[31].entry.input_buf[4].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[32].entry.latch[5]  (.D(\l_fifo.genblk1[32].entry.input_buf[5].X ),
    .GATE(\l_fifo.genblk1[32].entry.empty ),
    .RESET_B(net21),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[31].entry.input_buf[5].A ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[33].entry.input_buf[0].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[33].entry.input_buf[0].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[33].entry.input_buf[0].genblk1[0].mid ));
 sky130_fd_sc_hd__inv_2 \l_fifo.genblk1[33].entry.input_buf[0].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[33].entry.input_buf[0].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[33].entry.input_buf[0].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[33].entry.input_buf[1].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[33].entry.input_buf[1].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[33].entry.input_buf[1].genblk1[0].mid ));
 sky130_fd_sc_hd__inv_2 \l_fifo.genblk1[33].entry.input_buf[1].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[33].entry.input_buf[1].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[33].entry.input_buf[1].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[33].entry.input_buf[2].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[33].entry.input_buf[2].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[33].entry.input_buf[2].genblk1[0].mid ));
 sky130_fd_sc_hd__inv_2 \l_fifo.genblk1[33].entry.input_buf[2].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[33].entry.input_buf[2].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[33].entry.input_buf[2].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[33].entry.input_buf[3].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[33].entry.input_buf[3].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[33].entry.input_buf[3].genblk1[0].mid ));
 sky130_fd_sc_hd__clkinv_2 \l_fifo.genblk1[33].entry.input_buf[3].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[33].entry.input_buf[3].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[33].entry.input_buf[3].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[33].entry.input_buf[4].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[33].entry.input_buf[4].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[33].entry.input_buf[4].genblk1[0].mid ));
 sky130_fd_sc_hd__inv_2 \l_fifo.genblk1[33].entry.input_buf[4].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[33].entry.input_buf[4].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[33].entry.input_buf[4].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[33].entry.input_buf[5].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[33].entry.input_buf[5].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[33].entry.input_buf[5].genblk1[0].mid ));
 sky130_fd_sc_hd__clkinv_2 \l_fifo.genblk1[33].entry.input_buf[5].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[33].entry.input_buf[5].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[33].entry.input_buf[5].X ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[33].entry.latch[0]  (.D(\l_fifo.genblk1[33].entry.input_buf[0].X ),
    .GATE(\l_fifo.genblk1[33].entry.empty ),
    .RESET_B(net8),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[32].entry.input_buf[0].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[33].entry.latch[1]  (.D(\l_fifo.genblk1[33].entry.input_buf[1].X ),
    .GATE(\l_fifo.genblk1[33].entry.empty ),
    .RESET_B(net9),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[32].entry.input_buf[1].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[33].entry.latch[2]  (.D(\l_fifo.genblk1[33].entry.input_buf[2].X ),
    .GATE(\l_fifo.genblk1[33].entry.empty ),
    .RESET_B(net12),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[32].entry.input_buf[2].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[33].entry.latch[3]  (.D(\l_fifo.genblk1[33].entry.input_buf[3].X ),
    .GATE(\l_fifo.genblk1[33].entry.empty ),
    .RESET_B(net9),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[32].entry.input_buf[3].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[33].entry.latch[4]  (.D(\l_fifo.genblk1[33].entry.input_buf[4].X ),
    .GATE(\l_fifo.genblk1[33].entry.empty ),
    .RESET_B(net8),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[32].entry.input_buf[4].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[33].entry.latch[5]  (.D(\l_fifo.genblk1[33].entry.input_buf[5].X ),
    .GATE(\l_fifo.genblk1[33].entry.empty ),
    .RESET_B(net8),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[32].entry.input_buf[5].A ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[34].entry.input_buf[0].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[34].entry.input_buf[0].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[34].entry.input_buf[0].genblk1[0].mid ));
 sky130_fd_sc_hd__inv_2 \l_fifo.genblk1[34].entry.input_buf[0].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[34].entry.input_buf[0].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[34].entry.input_buf[0].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[34].entry.input_buf[1].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[34].entry.input_buf[1].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[34].entry.input_buf[1].genblk1[0].mid ));
 sky130_fd_sc_hd__inv_2 \l_fifo.genblk1[34].entry.input_buf[1].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[34].entry.input_buf[1].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[34].entry.input_buf[1].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[34].entry.input_buf[2].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[34].entry.input_buf[2].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[34].entry.input_buf[2].genblk1[0].mid ));
 sky130_fd_sc_hd__inv_2 \l_fifo.genblk1[34].entry.input_buf[2].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[34].entry.input_buf[2].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[34].entry.input_buf[2].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[34].entry.input_buf[3].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[34].entry.input_buf[3].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[34].entry.input_buf[3].genblk1[0].mid ));
 sky130_fd_sc_hd__inv_2 \l_fifo.genblk1[34].entry.input_buf[3].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[34].entry.input_buf[3].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[34].entry.input_buf[3].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[34].entry.input_buf[4].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[34].entry.input_buf[4].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[34].entry.input_buf[4].genblk1[0].mid ));
 sky130_fd_sc_hd__clkinv_2 \l_fifo.genblk1[34].entry.input_buf[4].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[34].entry.input_buf[4].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[34].entry.input_buf[4].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[34].entry.input_buf[5].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[34].entry.input_buf[5].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[34].entry.input_buf[5].genblk1[0].mid ));
 sky130_fd_sc_hd__inv_2 \l_fifo.genblk1[34].entry.input_buf[5].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[34].entry.input_buf[5].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[34].entry.input_buf[5].X ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[34].entry.latch[0]  (.D(\l_fifo.genblk1[34].entry.input_buf[0].X ),
    .GATE(\l_fifo.genblk1[34].entry.empty ),
    .RESET_B(net12),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[33].entry.input_buf[0].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[34].entry.latch[1]  (.D(\l_fifo.genblk1[34].entry.input_buf[1].X ),
    .GATE(\l_fifo.genblk1[34].entry.empty ),
    .RESET_B(net10),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[33].entry.input_buf[1].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[34].entry.latch[2]  (.D(\l_fifo.genblk1[34].entry.input_buf[2].X ),
    .GATE(\l_fifo.genblk1[34].entry.empty ),
    .RESET_B(net10),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[33].entry.input_buf[2].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[34].entry.latch[3]  (.D(\l_fifo.genblk1[34].entry.input_buf[3].X ),
    .GATE(\l_fifo.genblk1[34].entry.empty ),
    .RESET_B(net8),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[33].entry.input_buf[3].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[34].entry.latch[4]  (.D(\l_fifo.genblk1[34].entry.input_buf[4].X ),
    .GATE(\l_fifo.genblk1[34].entry.empty ),
    .RESET_B(net12),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[33].entry.input_buf[4].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[34].entry.latch[5]  (.D(\l_fifo.genblk1[34].entry.input_buf[5].X ),
    .GATE(\l_fifo.genblk1[34].entry.empty ),
    .RESET_B(net12),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[33].entry.input_buf[5].A ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[35].entry.input_buf[0].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[35].entry.input_buf[0].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[35].entry.input_buf[0].genblk1[0].mid ));
 sky130_fd_sc_hd__inv_2 \l_fifo.genblk1[35].entry.input_buf[0].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[35].entry.input_buf[0].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[35].entry.input_buf[0].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[35].entry.input_buf[1].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[35].entry.input_buf[1].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[35].entry.input_buf[1].genblk1[0].mid ));
 sky130_fd_sc_hd__inv_2 \l_fifo.genblk1[35].entry.input_buf[1].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[35].entry.input_buf[1].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[35].entry.input_buf[1].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[35].entry.input_buf[2].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[35].entry.input_buf[2].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[35].entry.input_buf[2].genblk1[0].mid ));
 sky130_fd_sc_hd__clkinv_2 \l_fifo.genblk1[35].entry.input_buf[2].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[35].entry.input_buf[2].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[35].entry.input_buf[2].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[35].entry.input_buf[3].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[35].entry.input_buf[3].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[35].entry.input_buf[3].genblk1[0].mid ));
 sky130_fd_sc_hd__inv_2 \l_fifo.genblk1[35].entry.input_buf[3].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[35].entry.input_buf[3].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[35].entry.input_buf[3].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[35].entry.input_buf[4].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[35].entry.input_buf[4].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[35].entry.input_buf[4].genblk1[0].mid ));
 sky130_fd_sc_hd__inv_2 \l_fifo.genblk1[35].entry.input_buf[4].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[35].entry.input_buf[4].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[35].entry.input_buf[4].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[35].entry.input_buf[5].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[35].entry.input_buf[5].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[35].entry.input_buf[5].genblk1[0].mid ));
 sky130_fd_sc_hd__clkinv_2 \l_fifo.genblk1[35].entry.input_buf[5].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[35].entry.input_buf[5].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[35].entry.input_buf[5].X ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[35].entry.latch[0]  (.D(\l_fifo.genblk1[35].entry.input_buf[0].X ),
    .GATE(\l_fifo.genblk1[35].entry.empty ),
    .RESET_B(net11),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[34].entry.input_buf[0].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[35].entry.latch[1]  (.D(\l_fifo.genblk1[35].entry.input_buf[1].X ),
    .GATE(\l_fifo.genblk1[35].entry.empty ),
    .RESET_B(net8),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[34].entry.input_buf[1].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[35].entry.latch[2]  (.D(\l_fifo.genblk1[35].entry.input_buf[2].X ),
    .GATE(\l_fifo.genblk1[35].entry.empty ),
    .RESET_B(net11),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[34].entry.input_buf[2].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[35].entry.latch[3]  (.D(\l_fifo.genblk1[35].entry.input_buf[3].X ),
    .GATE(\l_fifo.genblk1[35].entry.empty ),
    .RESET_B(net8),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[34].entry.input_buf[3].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[35].entry.latch[4]  (.D(\l_fifo.genblk1[35].entry.input_buf[4].X ),
    .GATE(\l_fifo.genblk1[35].entry.empty ),
    .RESET_B(net8),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[34].entry.input_buf[4].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[35].entry.latch[5]  (.D(\l_fifo.genblk1[35].entry.input_buf[5].X ),
    .GATE(\l_fifo.genblk1[35].entry.empty ),
    .RESET_B(net8),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[34].entry.input_buf[5].A ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[36].entry.input_buf[0].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[36].entry.input_buf[0].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[36].entry.input_buf[0].genblk1[0].mid ));
 sky130_fd_sc_hd__clkinv_2 \l_fifo.genblk1[36].entry.input_buf[0].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[36].entry.input_buf[0].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[36].entry.input_buf[0].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[36].entry.input_buf[1].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[36].entry.input_buf[1].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[36].entry.input_buf[1].genblk1[0].mid ));
 sky130_fd_sc_hd__inv_2 \l_fifo.genblk1[36].entry.input_buf[1].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[36].entry.input_buf[1].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[36].entry.input_buf[1].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[36].entry.input_buf[2].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[36].entry.input_buf[2].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[36].entry.input_buf[2].genblk1[0].mid ));
 sky130_fd_sc_hd__inv_2 \l_fifo.genblk1[36].entry.input_buf[2].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[36].entry.input_buf[2].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[36].entry.input_buf[2].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[36].entry.input_buf[3].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[36].entry.input_buf[3].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[36].entry.input_buf[3].genblk1[0].mid ));
 sky130_fd_sc_hd__inv_2 \l_fifo.genblk1[36].entry.input_buf[3].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[36].entry.input_buf[3].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[36].entry.input_buf[3].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[36].entry.input_buf[4].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[36].entry.input_buf[4].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[36].entry.input_buf[4].genblk1[0].mid ));
 sky130_fd_sc_hd__inv_2 \l_fifo.genblk1[36].entry.input_buf[4].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[36].entry.input_buf[4].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[36].entry.input_buf[4].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[36].entry.input_buf[5].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[36].entry.input_buf[5].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[36].entry.input_buf[5].genblk1[0].mid ));
 sky130_fd_sc_hd__clkinv_2 \l_fifo.genblk1[36].entry.input_buf[5].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[36].entry.input_buf[5].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[36].entry.input_buf[5].X ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[36].entry.latch[0]  (.D(\l_fifo.genblk1[36].entry.input_buf[0].X ),
    .GATE(\l_fifo.genblk1[36].entry.empty ),
    .RESET_B(net13),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[35].entry.input_buf[0].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[36].entry.latch[1]  (.D(\l_fifo.genblk1[36].entry.input_buf[1].X ),
    .GATE(\l_fifo.genblk1[36].entry.empty ),
    .RESET_B(net9),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[35].entry.input_buf[1].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[36].entry.latch[2]  (.D(\l_fifo.genblk1[36].entry.input_buf[2].X ),
    .GATE(\l_fifo.genblk1[36].entry.empty ),
    .RESET_B(net8),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[35].entry.input_buf[2].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[36].entry.latch[3]  (.D(\l_fifo.genblk1[36].entry.input_buf[3].X ),
    .GATE(\l_fifo.genblk1[36].entry.empty ),
    .RESET_B(net9),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[35].entry.input_buf[3].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[36].entry.latch[4]  (.D(\l_fifo.genblk1[36].entry.input_buf[4].X ),
    .GATE(\l_fifo.genblk1[36].entry.empty ),
    .RESET_B(net9),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[35].entry.input_buf[4].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[36].entry.latch[5]  (.D(\l_fifo.genblk1[36].entry.input_buf[5].X ),
    .GATE(\l_fifo.genblk1[36].entry.empty ),
    .RESET_B(net9),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[35].entry.input_buf[5].A ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[37].entry.input_buf[0].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[37].entry.input_buf[0].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[37].entry.input_buf[0].genblk1[0].mid ));
 sky130_fd_sc_hd__inv_2 \l_fifo.genblk1[37].entry.input_buf[0].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[37].entry.input_buf[0].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[37].entry.input_buf[0].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[37].entry.input_buf[1].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[37].entry.input_buf[1].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[37].entry.input_buf[1].genblk1[0].mid ));
 sky130_fd_sc_hd__inv_2 \l_fifo.genblk1[37].entry.input_buf[1].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[37].entry.input_buf[1].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[37].entry.input_buf[1].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[37].entry.input_buf[2].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[37].entry.input_buf[2].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[37].entry.input_buf[2].genblk1[0].mid ));
 sky130_fd_sc_hd__clkinv_2 \l_fifo.genblk1[37].entry.input_buf[2].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[37].entry.input_buf[2].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[37].entry.input_buf[2].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[37].entry.input_buf[3].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[37].entry.input_buf[3].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[37].entry.input_buf[3].genblk1[0].mid ));
 sky130_fd_sc_hd__inv_2 \l_fifo.genblk1[37].entry.input_buf[3].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[37].entry.input_buf[3].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[37].entry.input_buf[3].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[37].entry.input_buf[4].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[37].entry.input_buf[4].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[37].entry.input_buf[4].genblk1[0].mid ));
 sky130_fd_sc_hd__inv_2 \l_fifo.genblk1[37].entry.input_buf[4].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[37].entry.input_buf[4].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[37].entry.input_buf[4].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[37].entry.input_buf[5].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[37].entry.input_buf[5].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[37].entry.input_buf[5].genblk1[0].mid ));
 sky130_fd_sc_hd__inv_2 \l_fifo.genblk1[37].entry.input_buf[5].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[37].entry.input_buf[5].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[37].entry.input_buf[5].X ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[37].entry.latch[0]  (.D(\l_fifo.genblk1[37].entry.input_buf[0].X ),
    .GATE(\l_fifo.genblk1[37].entry.empty ),
    .RESET_B(net13),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[36].entry.input_buf[0].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[37].entry.latch[1]  (.D(\l_fifo.genblk1[37].entry.input_buf[1].X ),
    .GATE(\l_fifo.genblk1[37].entry.empty ),
    .RESET_B(net13),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[36].entry.input_buf[1].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[37].entry.latch[2]  (.D(\l_fifo.genblk1[37].entry.input_buf[2].X ),
    .GATE(\l_fifo.genblk1[37].entry.empty ),
    .RESET_B(net8),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[36].entry.input_buf[2].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[37].entry.latch[3]  (.D(\l_fifo.genblk1[37].entry.input_buf[3].X ),
    .GATE(\l_fifo.genblk1[37].entry.empty ),
    .RESET_B(net14),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[36].entry.input_buf[3].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[37].entry.latch[4]  (.D(\l_fifo.genblk1[37].entry.input_buf[4].X ),
    .GATE(\l_fifo.genblk1[37].entry.empty ),
    .RESET_B(net13),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[36].entry.input_buf[4].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[37].entry.latch[5]  (.D(\l_fifo.genblk1[37].entry.input_buf[5].X ),
    .GATE(\l_fifo.genblk1[37].entry.empty ),
    .RESET_B(net10),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[36].entry.input_buf[5].A ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[38].entry.input_buf[0].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[38].entry.input_buf[0].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[38].entry.input_buf[0].genblk1[0].mid ));
 sky130_fd_sc_hd__inv_2 \l_fifo.genblk1[38].entry.input_buf[0].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[38].entry.input_buf[0].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[38].entry.input_buf[0].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[38].entry.input_buf[1].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[38].entry.input_buf[1].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[38].entry.input_buf[1].genblk1[0].mid ));
 sky130_fd_sc_hd__inv_2 \l_fifo.genblk1[38].entry.input_buf[1].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[38].entry.input_buf[1].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[38].entry.input_buf[1].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[38].entry.input_buf[2].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[38].entry.input_buf[2].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[38].entry.input_buf[2].genblk1[0].mid ));
 sky130_fd_sc_hd__clkinv_2 \l_fifo.genblk1[38].entry.input_buf[2].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[38].entry.input_buf[2].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[38].entry.input_buf[2].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[38].entry.input_buf[3].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[38].entry.input_buf[3].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[38].entry.input_buf[3].genblk1[0].mid ));
 sky130_fd_sc_hd__inv_2 \l_fifo.genblk1[38].entry.input_buf[3].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[38].entry.input_buf[3].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[38].entry.input_buf[3].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[38].entry.input_buf[4].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[38].entry.input_buf[4].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[38].entry.input_buf[4].genblk1[0].mid ));
 sky130_fd_sc_hd__inv_2 \l_fifo.genblk1[38].entry.input_buf[4].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[38].entry.input_buf[4].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[38].entry.input_buf[4].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[38].entry.input_buf[5].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[38].entry.input_buf[5].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[38].entry.input_buf[5].genblk1[0].mid ));
 sky130_fd_sc_hd__clkinv_2 \l_fifo.genblk1[38].entry.input_buf[5].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[38].entry.input_buf[5].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[38].entry.input_buf[5].X ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[38].entry.latch[0]  (.D(\l_fifo.genblk1[38].entry.input_buf[0].X ),
    .GATE(\l_fifo.genblk1[38].entry.empty ),
    .RESET_B(net13),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[37].entry.input_buf[0].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[38].entry.latch[1]  (.D(\l_fifo.genblk1[38].entry.input_buf[1].X ),
    .GATE(\l_fifo.genblk1[38].entry.empty ),
    .RESET_B(net14),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[37].entry.input_buf[1].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[38].entry.latch[2]  (.D(\l_fifo.genblk1[38].entry.input_buf[2].X ),
    .GATE(\l_fifo.genblk1[38].entry.empty ),
    .RESET_B(net13),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[37].entry.input_buf[2].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[38].entry.latch[3]  (.D(\l_fifo.genblk1[38].entry.input_buf[3].X ),
    .GATE(\l_fifo.genblk1[38].entry.empty ),
    .RESET_B(net14),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[37].entry.input_buf[3].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[38].entry.latch[4]  (.D(\l_fifo.genblk1[38].entry.input_buf[4].X ),
    .GATE(\l_fifo.genblk1[38].entry.empty ),
    .RESET_B(net13),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[37].entry.input_buf[4].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[38].entry.latch[5]  (.D(\l_fifo.genblk1[38].entry.input_buf[5].X ),
    .GATE(\l_fifo.genblk1[38].entry.empty ),
    .RESET_B(net14),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[37].entry.input_buf[5].A ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[39].entry.input_buf[0].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[39].entry.input_buf[0].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[39].entry.input_buf[0].genblk1[0].mid ));
 sky130_fd_sc_hd__inv_2 \l_fifo.genblk1[39].entry.input_buf[0].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[39].entry.input_buf[0].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[39].entry.input_buf[0].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[39].entry.input_buf[1].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[39].entry.input_buf[1].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[39].entry.input_buf[1].genblk1[0].mid ));
 sky130_fd_sc_hd__inv_2 \l_fifo.genblk1[39].entry.input_buf[1].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[39].entry.input_buf[1].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[39].entry.input_buf[1].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[39].entry.input_buf[2].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[39].entry.input_buf[2].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[39].entry.input_buf[2].genblk1[0].mid ));
 sky130_fd_sc_hd__inv_2 \l_fifo.genblk1[39].entry.input_buf[2].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[39].entry.input_buf[2].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[39].entry.input_buf[2].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[39].entry.input_buf[3].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[39].entry.input_buf[3].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[39].entry.input_buf[3].genblk1[0].mid ));
 sky130_fd_sc_hd__inv_2 \l_fifo.genblk1[39].entry.input_buf[3].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[39].entry.input_buf[3].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[39].entry.input_buf[3].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[39].entry.input_buf[4].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[39].entry.input_buf[4].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[39].entry.input_buf[4].genblk1[0].mid ));
 sky130_fd_sc_hd__inv_2 \l_fifo.genblk1[39].entry.input_buf[4].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[39].entry.input_buf[4].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[39].entry.input_buf[4].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[39].entry.input_buf[5].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[39].entry.input_buf[5].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[39].entry.input_buf[5].genblk1[0].mid ));
 sky130_fd_sc_hd__inv_2 \l_fifo.genblk1[39].entry.input_buf[5].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[39].entry.input_buf[5].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[39].entry.input_buf[5].X ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[39].entry.latch[0]  (.D(\l_fifo.genblk1[39].entry.input_buf[0].X ),
    .GATE(\l_fifo.genblk1[39].entry.empty ),
    .RESET_B(net15),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[38].entry.input_buf[0].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[39].entry.latch[1]  (.D(\l_fifo.genblk1[39].entry.input_buf[1].X ),
    .GATE(\l_fifo.genblk1[39].entry.empty ),
    .RESET_B(net14),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[38].entry.input_buf[1].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[39].entry.latch[2]  (.D(\l_fifo.genblk1[39].entry.input_buf[2].X ),
    .GATE(\l_fifo.genblk1[39].entry.empty ),
    .RESET_B(net15),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[38].entry.input_buf[2].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[39].entry.latch[3]  (.D(\l_fifo.genblk1[39].entry.input_buf[3].X ),
    .GATE(\l_fifo.genblk1[39].entry.empty ),
    .RESET_B(net14),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[38].entry.input_buf[3].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[39].entry.latch[4]  (.D(\l_fifo.genblk1[39].entry.input_buf[4].X ),
    .GATE(\l_fifo.genblk1[39].entry.empty ),
    .RESET_B(net33),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[38].entry.input_buf[4].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[39].entry.latch[5]  (.D(\l_fifo.genblk1[39].entry.input_buf[5].X ),
    .GATE(\l_fifo.genblk1[39].entry.empty ),
    .RESET_B(net15),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[38].entry.input_buf[5].A ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[3].entry.input_buf[0].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[3].entry.input_buf[0].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[3].entry.input_buf[0].genblk1[0].mid ));
 sky130_fd_sc_hd__clkinv_2 \l_fifo.genblk1[3].entry.input_buf[0].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[3].entry.input_buf[0].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[3].entry.input_buf[0].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[3].entry.input_buf[1].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[3].entry.input_buf[1].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[3].entry.input_buf[1].genblk1[0].mid ));
 sky130_fd_sc_hd__clkinv_2 \l_fifo.genblk1[3].entry.input_buf[1].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[3].entry.input_buf[1].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[3].entry.input_buf[1].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[3].entry.input_buf[2].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[3].entry.input_buf[2].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[3].entry.input_buf[2].genblk1[0].mid ));
 sky130_fd_sc_hd__clkinv_2 \l_fifo.genblk1[3].entry.input_buf[2].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[3].entry.input_buf[2].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[3].entry.input_buf[2].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[3].entry.input_buf[3].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[3].entry.input_buf[3].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[3].entry.input_buf[3].genblk1[0].mid ));
 sky130_fd_sc_hd__inv_2 \l_fifo.genblk1[3].entry.input_buf[3].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[3].entry.input_buf[3].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[3].entry.input_buf[3].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[3].entry.input_buf[4].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[3].entry.input_buf[4].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[3].entry.input_buf[4].genblk1[0].mid ));
 sky130_fd_sc_hd__clkinv_2 \l_fifo.genblk1[3].entry.input_buf[4].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[3].entry.input_buf[4].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[3].entry.input_buf[4].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[3].entry.input_buf[5].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[3].entry.input_buf[5].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[3].entry.input_buf[5].genblk1[0].mid ));
 sky130_fd_sc_hd__clkinv_2 \l_fifo.genblk1[3].entry.input_buf[5].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[3].entry.input_buf[5].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[3].entry.input_buf[5].X ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[3].entry.latch[0]  (.D(\l_fifo.genblk1[3].entry.input_buf[0].X ),
    .GATE(\l_fifo.genblk1[3].entry.empty ),
    .RESET_B(net26),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[2].entry.input_buf[0].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[3].entry.latch[1]  (.D(\l_fifo.genblk1[3].entry.input_buf[1].X ),
    .GATE(\l_fifo.genblk1[3].entry.empty ),
    .RESET_B(net26),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[2].entry.input_buf[1].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[3].entry.latch[2]  (.D(\l_fifo.genblk1[3].entry.input_buf[2].X ),
    .GATE(\l_fifo.genblk1[3].entry.empty ),
    .RESET_B(net26),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[2].entry.input_buf[2].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[3].entry.latch[3]  (.D(\l_fifo.genblk1[3].entry.input_buf[3].X ),
    .GATE(\l_fifo.genblk1[3].entry.empty ),
    .RESET_B(net26),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[2].entry.input_buf[3].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[3].entry.latch[4]  (.D(\l_fifo.genblk1[3].entry.input_buf[4].X ),
    .GATE(\l_fifo.genblk1[3].entry.empty ),
    .RESET_B(net27),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[2].entry.input_buf[4].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[3].entry.latch[5]  (.D(\l_fifo.genblk1[3].entry.input_buf[5].X ),
    .GATE(\l_fifo.genblk1[3].entry.empty ),
    .RESET_B(net32),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[2].entry.input_buf[5].A ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[40].entry.input_buf[0].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[40].entry.input_buf[0].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[40].entry.input_buf[0].genblk1[0].mid ));
 sky130_fd_sc_hd__clkinv_2 \l_fifo.genblk1[40].entry.input_buf[0].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[40].entry.input_buf[0].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[40].entry.input_buf[0].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[40].entry.input_buf[1].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[40].entry.input_buf[1].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[40].entry.input_buf[1].genblk1[0].mid ));
 sky130_fd_sc_hd__clkinv_2 \l_fifo.genblk1[40].entry.input_buf[1].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[40].entry.input_buf[1].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[40].entry.input_buf[1].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[40].entry.input_buf[2].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[40].entry.input_buf[2].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[40].entry.input_buf[2].genblk1[0].mid ));
 sky130_fd_sc_hd__clkinv_2 \l_fifo.genblk1[40].entry.input_buf[2].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[40].entry.input_buf[2].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[40].entry.input_buf[2].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[40].entry.input_buf[3].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[40].entry.input_buf[3].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[40].entry.input_buf[3].genblk1[0].mid ));
 sky130_fd_sc_hd__clkinv_2 \l_fifo.genblk1[40].entry.input_buf[3].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[40].entry.input_buf[3].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[40].entry.input_buf[3].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[40].entry.input_buf[4].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[40].entry.input_buf[4].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[40].entry.input_buf[4].genblk1[0].mid ));
 sky130_fd_sc_hd__clkinv_2 \l_fifo.genblk1[40].entry.input_buf[4].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[40].entry.input_buf[4].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[40].entry.input_buf[4].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[40].entry.input_buf[5].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[40].entry.input_buf[5].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[40].entry.input_buf[5].genblk1[0].mid ));
 sky130_fd_sc_hd__inv_2 \l_fifo.genblk1[40].entry.input_buf[5].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[40].entry.input_buf[5].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[40].entry.input_buf[5].X ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[40].entry.latch[0]  (.D(\l_fifo.genblk1[40].entry.input_buf[0].X ),
    .GATE(\l_fifo.genblk1[40].entry.empty ),
    .RESET_B(net33),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[39].entry.input_buf[0].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[40].entry.latch[1]  (.D(\l_fifo.genblk1[40].entry.input_buf[1].X ),
    .GATE(\l_fifo.genblk1[40].entry.empty ),
    .RESET_B(net33),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[39].entry.input_buf[1].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[40].entry.latch[2]  (.D(\l_fifo.genblk1[40].entry.input_buf[2].X ),
    .GATE(\l_fifo.genblk1[40].entry.empty ),
    .RESET_B(net33),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[39].entry.input_buf[2].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[40].entry.latch[3]  (.D(\l_fifo.genblk1[40].entry.input_buf[3].X ),
    .GATE(\l_fifo.genblk1[40].entry.empty ),
    .RESET_B(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[39].entry.input_buf[3].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[40].entry.latch[4]  (.D(\l_fifo.genblk1[40].entry.input_buf[4].X ),
    .GATE(\l_fifo.genblk1[40].entry.empty ),
    .RESET_B(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[39].entry.input_buf[4].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[40].entry.latch[5]  (.D(\l_fifo.genblk1[40].entry.input_buf[5].X ),
    .GATE(\l_fifo.genblk1[40].entry.empty ),
    .RESET_B(net15),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[39].entry.input_buf[5].A ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[41].entry.input_buf[0].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[41].entry.input_buf[0].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[41].entry.input_buf[0].genblk1[0].mid ));
 sky130_fd_sc_hd__clkinv_2 \l_fifo.genblk1[41].entry.input_buf[0].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[41].entry.input_buf[0].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[41].entry.input_buf[0].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[41].entry.input_buf[1].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[41].entry.input_buf[1].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[41].entry.input_buf[1].genblk1[0].mid ));
 sky130_fd_sc_hd__inv_2 \l_fifo.genblk1[41].entry.input_buf[1].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[41].entry.input_buf[1].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[41].entry.input_buf[1].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[41].entry.input_buf[2].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[41].entry.input_buf[2].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[41].entry.input_buf[2].genblk1[0].mid ));
 sky130_fd_sc_hd__inv_2 \l_fifo.genblk1[41].entry.input_buf[2].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[41].entry.input_buf[2].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[41].entry.input_buf[2].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[41].entry.input_buf[3].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[41].entry.input_buf[3].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[41].entry.input_buf[3].genblk1[0].mid ));
 sky130_fd_sc_hd__inv_2 \l_fifo.genblk1[41].entry.input_buf[3].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[41].entry.input_buf[3].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[41].entry.input_buf[3].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[41].entry.input_buf[4].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[41].entry.input_buf[4].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[41].entry.input_buf[4].genblk1[0].mid ));
 sky130_fd_sc_hd__clkinv_2 \l_fifo.genblk1[41].entry.input_buf[4].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[41].entry.input_buf[4].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[41].entry.input_buf[4].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[41].entry.input_buf[5].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[41].entry.input_buf[5].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[41].entry.input_buf[5].genblk1[0].mid ));
 sky130_fd_sc_hd__clkinv_2 \l_fifo.genblk1[41].entry.input_buf[5].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[41].entry.input_buf[5].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[41].entry.input_buf[5].X ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[41].entry.latch[0]  (.D(\l_fifo.genblk1[41].entry.input_buf[0].X ),
    .GATE(\l_fifo.genblk1[41].entry.empty ),
    .RESET_B(net14),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[40].entry.input_buf[0].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[41].entry.latch[1]  (.D(\l_fifo.genblk1[41].entry.input_buf[1].X ),
    .GATE(\l_fifo.genblk1[41].entry.empty ),
    .RESET_B(net33),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[40].entry.input_buf[1].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[41].entry.latch[2]  (.D(\l_fifo.genblk1[41].entry.input_buf[2].X ),
    .GATE(\l_fifo.genblk1[41].entry.empty ),
    .RESET_B(net33),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[40].entry.input_buf[2].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[41].entry.latch[3]  (.D(\l_fifo.genblk1[41].entry.input_buf[3].X ),
    .GATE(\l_fifo.genblk1[41].entry.empty ),
    .RESET_B(net33),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[40].entry.input_buf[3].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[41].entry.latch[4]  (.D(\l_fifo.genblk1[41].entry.input_buf[4].X ),
    .GATE(\l_fifo.genblk1[41].entry.empty ),
    .RESET_B(net33),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[40].entry.input_buf[4].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[41].entry.latch[5]  (.D(\l_fifo.genblk1[41].entry.input_buf[5].X ),
    .GATE(\l_fifo.genblk1[41].entry.empty ),
    .RESET_B(net33),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[40].entry.input_buf[5].A ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[42].entry.input_buf[0].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[42].entry.input_buf[0].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[42].entry.input_buf[0].genblk1[0].mid ));
 sky130_fd_sc_hd__clkinv_2 \l_fifo.genblk1[42].entry.input_buf[0].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[42].entry.input_buf[0].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[42].entry.input_buf[0].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[42].entry.input_buf[1].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[42].entry.input_buf[1].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[42].entry.input_buf[1].genblk1[0].mid ));
 sky130_fd_sc_hd__clkinv_2 \l_fifo.genblk1[42].entry.input_buf[1].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[42].entry.input_buf[1].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[42].entry.input_buf[1].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[42].entry.input_buf[2].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[42].entry.input_buf[2].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[42].entry.input_buf[2].genblk1[0].mid ));
 sky130_fd_sc_hd__clkinv_2 \l_fifo.genblk1[42].entry.input_buf[2].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[42].entry.input_buf[2].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[42].entry.input_buf[2].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[42].entry.input_buf[3].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[42].entry.input_buf[3].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[42].entry.input_buf[3].genblk1[0].mid ));
 sky130_fd_sc_hd__clkinv_2 \l_fifo.genblk1[42].entry.input_buf[3].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[42].entry.input_buf[3].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[42].entry.input_buf[3].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[42].entry.input_buf[4].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[42].entry.input_buf[4].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[42].entry.input_buf[4].genblk1[0].mid ));
 sky130_fd_sc_hd__clkinv_2 \l_fifo.genblk1[42].entry.input_buf[4].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[42].entry.input_buf[4].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[42].entry.input_buf[4].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[42].entry.input_buf[5].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[42].entry.input_buf[5].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[42].entry.input_buf[5].genblk1[0].mid ));
 sky130_fd_sc_hd__clkinv_2 \l_fifo.genblk1[42].entry.input_buf[5].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[42].entry.input_buf[5].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[42].entry.input_buf[5].X ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[42].entry.latch[0]  (.D(\l_fifo.genblk1[42].entry.input_buf[0].X ),
    .GATE(\l_fifo.genblk1[42].entry.empty ),
    .RESET_B(net14),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[41].entry.input_buf[0].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[42].entry.latch[1]  (.D(\l_fifo.genblk1[42].entry.input_buf[1].X ),
    .GATE(\l_fifo.genblk1[42].entry.empty ),
    .RESET_B(net23),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[41].entry.input_buf[1].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[42].entry.latch[2]  (.D(\l_fifo.genblk1[42].entry.input_buf[2].X ),
    .GATE(\l_fifo.genblk1[42].entry.empty ),
    .RESET_B(net33),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[41].entry.input_buf[2].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[42].entry.latch[3]  (.D(\l_fifo.genblk1[42].entry.input_buf[3].X ),
    .GATE(\l_fifo.genblk1[42].entry.empty ),
    .RESET_B(net22),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[41].entry.input_buf[3].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[42].entry.latch[4]  (.D(\l_fifo.genblk1[42].entry.input_buf[4].X ),
    .GATE(\l_fifo.genblk1[42].entry.empty ),
    .RESET_B(net34),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[41].entry.input_buf[4].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[42].entry.latch[5]  (.D(\l_fifo.genblk1[42].entry.input_buf[5].X ),
    .GATE(\l_fifo.genblk1[42].entry.empty ),
    .RESET_B(net34),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[41].entry.input_buf[5].A ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[43].entry.input_buf[0].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[43].entry.input_buf[0].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[43].entry.input_buf[0].genblk1[0].mid ));
 sky130_fd_sc_hd__inv_2 \l_fifo.genblk1[43].entry.input_buf[0].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[43].entry.input_buf[0].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[43].entry.input_buf[0].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[43].entry.input_buf[1].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[43].entry.input_buf[1].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[43].entry.input_buf[1].genblk1[0].mid ));
 sky130_fd_sc_hd__inv_2 \l_fifo.genblk1[43].entry.input_buf[1].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[43].entry.input_buf[1].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[43].entry.input_buf[1].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[43].entry.input_buf[2].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[43].entry.input_buf[2].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[43].entry.input_buf[2].genblk1[0].mid ));
 sky130_fd_sc_hd__inv_2 \l_fifo.genblk1[43].entry.input_buf[2].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[43].entry.input_buf[2].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[43].entry.input_buf[2].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[43].entry.input_buf[3].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[43].entry.input_buf[3].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[43].entry.input_buf[3].genblk1[0].mid ));
 sky130_fd_sc_hd__inv_2 \l_fifo.genblk1[43].entry.input_buf[3].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[43].entry.input_buf[3].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[43].entry.input_buf[3].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[43].entry.input_buf[4].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[43].entry.input_buf[4].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[43].entry.input_buf[4].genblk1[0].mid ));
 sky130_fd_sc_hd__inv_2 \l_fifo.genblk1[43].entry.input_buf[4].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[43].entry.input_buf[4].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[43].entry.input_buf[4].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[43].entry.input_buf[5].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[43].entry.input_buf[5].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[43].entry.input_buf[5].genblk1[0].mid ));
 sky130_fd_sc_hd__clkinv_2 \l_fifo.genblk1[43].entry.input_buf[5].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[43].entry.input_buf[5].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[43].entry.input_buf[5].X ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[43].entry.latch[0]  (.D(\l_fifo.genblk1[43].entry.input_buf[0].X ),
    .GATE(\l_fifo.genblk1[43].entry.empty ),
    .RESET_B(net24),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[42].entry.input_buf[0].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[43].entry.latch[1]  (.D(\l_fifo.genblk1[43].entry.input_buf[1].X ),
    .GATE(\l_fifo.genblk1[43].entry.empty ),
    .RESET_B(net23),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[42].entry.input_buf[1].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[43].entry.latch[2]  (.D(\l_fifo.genblk1[43].entry.input_buf[2].X ),
    .GATE(\l_fifo.genblk1[43].entry.empty ),
    .RESET_B(net24),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[42].entry.input_buf[2].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[43].entry.latch[3]  (.D(\l_fifo.genblk1[43].entry.input_buf[3].X ),
    .GATE(\l_fifo.genblk1[43].entry.empty ),
    .RESET_B(net24),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[42].entry.input_buf[3].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[43].entry.latch[4]  (.D(\l_fifo.genblk1[43].entry.input_buf[4].X ),
    .GATE(\l_fifo.genblk1[43].entry.empty ),
    .RESET_B(net42),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[42].entry.input_buf[4].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[43].entry.latch[5]  (.D(\l_fifo.genblk1[43].entry.input_buf[5].X ),
    .GATE(\l_fifo.genblk1[43].entry.empty ),
    .RESET_B(net23),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[42].entry.input_buf[5].A ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[44].entry.input_buf[0].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[44].entry.input_buf[0].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[44].entry.input_buf[0].genblk1[0].mid ));
 sky130_fd_sc_hd__clkinv_2 \l_fifo.genblk1[44].entry.input_buf[0].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[44].entry.input_buf[0].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[44].entry.input_buf[0].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[44].entry.input_buf[1].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[44].entry.input_buf[1].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[44].entry.input_buf[1].genblk1[0].mid ));
 sky130_fd_sc_hd__inv_2 \l_fifo.genblk1[44].entry.input_buf[1].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[44].entry.input_buf[1].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[44].entry.input_buf[1].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[44].entry.input_buf[2].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[44].entry.input_buf[2].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[44].entry.input_buf[2].genblk1[0].mid ));
 sky130_fd_sc_hd__inv_2 \l_fifo.genblk1[44].entry.input_buf[2].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[44].entry.input_buf[2].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[44].entry.input_buf[2].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[44].entry.input_buf[3].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[44].entry.input_buf[3].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[44].entry.input_buf[3].genblk1[0].mid ));
 sky130_fd_sc_hd__inv_2 \l_fifo.genblk1[44].entry.input_buf[3].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[44].entry.input_buf[3].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[44].entry.input_buf[3].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[44].entry.input_buf[4].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[44].entry.input_buf[4].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[44].entry.input_buf[4].genblk1[0].mid ));
 sky130_fd_sc_hd__inv_2 \l_fifo.genblk1[44].entry.input_buf[4].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[44].entry.input_buf[4].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[44].entry.input_buf[4].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[44].entry.input_buf[5].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[44].entry.input_buf[5].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[44].entry.input_buf[5].genblk1[0].mid ));
 sky130_fd_sc_hd__inv_2 \l_fifo.genblk1[44].entry.input_buf[5].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[44].entry.input_buf[5].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[44].entry.input_buf[5].X ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[44].entry.latch[0]  (.D(\l_fifo.genblk1[44].entry.input_buf[0].X ),
    .GATE(\l_fifo.genblk1[44].entry.empty ),
    .RESET_B(net24),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[43].entry.input_buf[0].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[44].entry.latch[1]  (.D(\l_fifo.genblk1[44].entry.input_buf[1].X ),
    .GATE(\l_fifo.genblk1[44].entry.empty ),
    .RESET_B(net24),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[43].entry.input_buf[1].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[44].entry.latch[2]  (.D(\l_fifo.genblk1[44].entry.input_buf[2].X ),
    .GATE(\l_fifo.genblk1[44].entry.empty ),
    .RESET_B(net24),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[43].entry.input_buf[2].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[44].entry.latch[3]  (.D(\l_fifo.genblk1[44].entry.input_buf[3].X ),
    .GATE(\l_fifo.genblk1[44].entry.empty ),
    .RESET_B(net22),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[43].entry.input_buf[3].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[44].entry.latch[4]  (.D(\l_fifo.genblk1[44].entry.input_buf[4].X ),
    .GATE(\l_fifo.genblk1[44].entry.empty ),
    .RESET_B(net23),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[43].entry.input_buf[4].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[44].entry.latch[5]  (.D(\l_fifo.genblk1[44].entry.input_buf[5].X ),
    .GATE(\l_fifo.genblk1[44].entry.empty ),
    .RESET_B(net24),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[43].entry.input_buf[5].A ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[45].entry.input_buf[0].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[45].entry.input_buf[0].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[45].entry.input_buf[0].genblk1[0].mid ));
 sky130_fd_sc_hd__inv_2 \l_fifo.genblk1[45].entry.input_buf[0].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[45].entry.input_buf[0].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[45].entry.input_buf[0].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[45].entry.input_buf[1].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[45].entry.input_buf[1].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[45].entry.input_buf[1].genblk1[0].mid ));
 sky130_fd_sc_hd__clkinv_2 \l_fifo.genblk1[45].entry.input_buf[1].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[45].entry.input_buf[1].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[45].entry.input_buf[1].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[45].entry.input_buf[2].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[45].entry.input_buf[2].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[45].entry.input_buf[2].genblk1[0].mid ));
 sky130_fd_sc_hd__inv_2 \l_fifo.genblk1[45].entry.input_buf[2].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[45].entry.input_buf[2].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[45].entry.input_buf[2].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[45].entry.input_buf[3].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[45].entry.input_buf[3].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[45].entry.input_buf[3].genblk1[0].mid ));
 sky130_fd_sc_hd__clkinv_2 \l_fifo.genblk1[45].entry.input_buf[3].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[45].entry.input_buf[3].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[45].entry.input_buf[3].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[45].entry.input_buf[4].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[45].entry.input_buf[4].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[45].entry.input_buf[4].genblk1[0].mid ));
 sky130_fd_sc_hd__inv_2 \l_fifo.genblk1[45].entry.input_buf[4].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[45].entry.input_buf[4].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[45].entry.input_buf[4].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[45].entry.input_buf[5].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[45].entry.input_buf[5].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[45].entry.input_buf[5].genblk1[0].mid ));
 sky130_fd_sc_hd__clkinv_2 \l_fifo.genblk1[45].entry.input_buf[5].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[45].entry.input_buf[5].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[45].entry.input_buf[5].X ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[45].entry.latch[0]  (.D(\l_fifo.genblk1[45].entry.input_buf[0].X ),
    .GATE(\l_fifo.genblk1[45].entry.empty ),
    .RESET_B(net28),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[44].entry.input_buf[0].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[45].entry.latch[1]  (.D(\l_fifo.genblk1[45].entry.input_buf[1].X ),
    .GATE(\l_fifo.genblk1[45].entry.empty ),
    .RESET_B(net23),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[44].entry.input_buf[1].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[45].entry.latch[2]  (.D(\l_fifo.genblk1[45].entry.input_buf[2].X ),
    .GATE(\l_fifo.genblk1[45].entry.empty ),
    .RESET_B(net28),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[44].entry.input_buf[2].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[45].entry.latch[3]  (.D(\l_fifo.genblk1[45].entry.input_buf[3].X ),
    .GATE(\l_fifo.genblk1[45].entry.empty ),
    .RESET_B(net25),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[44].entry.input_buf[3].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[45].entry.latch[4]  (.D(\l_fifo.genblk1[45].entry.input_buf[4].X ),
    .GATE(\l_fifo.genblk1[45].entry.empty ),
    .RESET_B(net28),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[44].entry.input_buf[4].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[45].entry.latch[5]  (.D(\l_fifo.genblk1[45].entry.input_buf[5].X ),
    .GATE(\l_fifo.genblk1[45].entry.empty ),
    .RESET_B(net28),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[44].entry.input_buf[5].A ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[46].entry.input_buf[0].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[46].entry.input_buf[0].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[46].entry.input_buf[0].genblk1[0].mid ));
 sky130_fd_sc_hd__inv_2 \l_fifo.genblk1[46].entry.input_buf[0].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[46].entry.input_buf[0].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[46].entry.input_buf[0].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[46].entry.input_buf[1].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[46].entry.input_buf[1].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[46].entry.input_buf[1].genblk1[0].mid ));
 sky130_fd_sc_hd__inv_2 \l_fifo.genblk1[46].entry.input_buf[1].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[46].entry.input_buf[1].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[46].entry.input_buf[1].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[46].entry.input_buf[2].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[46].entry.input_buf[2].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[46].entry.input_buf[2].genblk1[0].mid ));
 sky130_fd_sc_hd__inv_2 \l_fifo.genblk1[46].entry.input_buf[2].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[46].entry.input_buf[2].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[46].entry.input_buf[2].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[46].entry.input_buf[3].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[46].entry.input_buf[3].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[46].entry.input_buf[3].genblk1[0].mid ));
 sky130_fd_sc_hd__clkinv_2 \l_fifo.genblk1[46].entry.input_buf[3].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[46].entry.input_buf[3].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[46].entry.input_buf[3].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[46].entry.input_buf[4].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[46].entry.input_buf[4].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[46].entry.input_buf[4].genblk1[0].mid ));
 sky130_fd_sc_hd__clkinv_2 \l_fifo.genblk1[46].entry.input_buf[4].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[46].entry.input_buf[4].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[46].entry.input_buf[4].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[46].entry.input_buf[5].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[46].entry.input_buf[5].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[46].entry.input_buf[5].genblk1[0].mid ));
 sky130_fd_sc_hd__inv_2 \l_fifo.genblk1[46].entry.input_buf[5].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[46].entry.input_buf[5].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[46].entry.input_buf[5].X ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[46].entry.latch[0]  (.D(\l_fifo.genblk1[46].entry.input_buf[0].X ),
    .GATE(\l_fifo.genblk1[46].entry.empty ),
    .RESET_B(net29),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[45].entry.input_buf[0].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[46].entry.latch[1]  (.D(\l_fifo.genblk1[46].entry.input_buf[1].X ),
    .GATE(\l_fifo.genblk1[46].entry.empty ),
    .RESET_B(net23),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[45].entry.input_buf[1].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[46].entry.latch[2]  (.D(\l_fifo.genblk1[46].entry.input_buf[2].X ),
    .GATE(\l_fifo.genblk1[46].entry.empty ),
    .RESET_B(net28),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[45].entry.input_buf[2].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[46].entry.latch[3]  (.D(\l_fifo.genblk1[46].entry.input_buf[3].X ),
    .GATE(\l_fifo.genblk1[46].entry.empty ),
    .RESET_B(net27),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[45].entry.input_buf[3].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[46].entry.latch[4]  (.D(\l_fifo.genblk1[46].entry.input_buf[4].X ),
    .GATE(\l_fifo.genblk1[46].entry.empty ),
    .RESET_B(net26),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[45].entry.input_buf[4].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[46].entry.latch[5]  (.D(\l_fifo.genblk1[46].entry.input_buf[5].X ),
    .GATE(\l_fifo.genblk1[46].entry.empty ),
    .RESET_B(net28),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[45].entry.input_buf[5].A ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[47].entry.input_buf[0].genblk1[0].genblk1.inv_first  (.A(\data_in_buffer[0].X ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[47].entry.input_buf[0].genblk1[0].mid ));
 sky130_fd_sc_hd__inv_2 \l_fifo.genblk1[47].entry.input_buf[0].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[47].entry.input_buf[0].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[47].entry.input_buf[0].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[47].entry.input_buf[1].genblk1[0].genblk1.inv_first  (.A(\data_in_buffer[1].X ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[47].entry.input_buf[1].genblk1[0].mid ));
 sky130_fd_sc_hd__inv_2 \l_fifo.genblk1[47].entry.input_buf[1].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[47].entry.input_buf[1].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[47].entry.input_buf[1].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[47].entry.input_buf[2].genblk1[0].genblk1.inv_first  (.A(\data_in_buffer[2].X ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[47].entry.input_buf[2].genblk1[0].mid ));
 sky130_fd_sc_hd__inv_2 \l_fifo.genblk1[47].entry.input_buf[2].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[47].entry.input_buf[2].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[47].entry.input_buf[2].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[47].entry.input_buf[3].genblk1[0].genblk1.inv_first  (.A(\data_in_buffer[3].X ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[47].entry.input_buf[3].genblk1[0].mid ));
 sky130_fd_sc_hd__inv_2 \l_fifo.genblk1[47].entry.input_buf[3].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[47].entry.input_buf[3].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[47].entry.input_buf[3].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[47].entry.input_buf[4].genblk1[0].genblk1.inv_first  (.A(\data_in_buffer[4].X ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[47].entry.input_buf[4].genblk1[0].mid ));
 sky130_fd_sc_hd__clkinv_2 \l_fifo.genblk1[47].entry.input_buf[4].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[47].entry.input_buf[4].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[47].entry.input_buf[4].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[47].entry.input_buf[5].genblk1[0].genblk1.inv_first  (.A(\data_in_buffer[5].X ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[47].entry.input_buf[5].genblk1[0].mid ));
 sky130_fd_sc_hd__inv_2 \l_fifo.genblk1[47].entry.input_buf[5].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[47].entry.input_buf[5].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[47].entry.input_buf[5].X ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[47].entry.latch[0]  (.D(\l_fifo.genblk1[47].entry.input_buf[0].X ),
    .GATE(\l_fifo.genblk1[47].entry.empty ),
    .RESET_B(net27),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[46].entry.input_buf[0].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[47].entry.latch[1]  (.D(\l_fifo.genblk1[47].entry.input_buf[1].X ),
    .GATE(\l_fifo.genblk1[47].entry.empty ),
    .RESET_B(net28),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[46].entry.input_buf[1].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[47].entry.latch[2]  (.D(\l_fifo.genblk1[47].entry.input_buf[2].X ),
    .GATE(\l_fifo.genblk1[47].entry.empty ),
    .RESET_B(net30),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[46].entry.input_buf[2].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[47].entry.latch[3]  (.D(\l_fifo.genblk1[47].entry.input_buf[3].X ),
    .GATE(\l_fifo.genblk1[47].entry.empty ),
    .RESET_B(net27),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[46].entry.input_buf[3].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[47].entry.latch[4]  (.D(\l_fifo.genblk1[47].entry.input_buf[4].X ),
    .GATE(\l_fifo.genblk1[47].entry.empty ),
    .RESET_B(net26),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[46].entry.input_buf[4].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[47].entry.latch[5]  (.D(\l_fifo.genblk1[47].entry.input_buf[5].X ),
    .GATE(\l_fifo.genblk1[47].entry.empty ),
    .RESET_B(net27),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[46].entry.input_buf[5].A ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[4].entry.input_buf[0].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[4].entry.input_buf[0].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[4].entry.input_buf[0].genblk1[0].mid ));
 sky130_fd_sc_hd__clkinv_2 \l_fifo.genblk1[4].entry.input_buf[0].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[4].entry.input_buf[0].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[4].entry.input_buf[0].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[4].entry.input_buf[1].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[4].entry.input_buf[1].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[4].entry.input_buf[1].genblk1[0].mid ));
 sky130_fd_sc_hd__clkinv_2 \l_fifo.genblk1[4].entry.input_buf[1].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[4].entry.input_buf[1].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[4].entry.input_buf[1].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[4].entry.input_buf[2].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[4].entry.input_buf[2].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[4].entry.input_buf[2].genblk1[0].mid ));
 sky130_fd_sc_hd__clkinv_2 \l_fifo.genblk1[4].entry.input_buf[2].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[4].entry.input_buf[2].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[4].entry.input_buf[2].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[4].entry.input_buf[3].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[4].entry.input_buf[3].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[4].entry.input_buf[3].genblk1[0].mid ));
 sky130_fd_sc_hd__inv_2 \l_fifo.genblk1[4].entry.input_buf[3].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[4].entry.input_buf[3].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[4].entry.input_buf[3].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[4].entry.input_buf[4].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[4].entry.input_buf[4].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[4].entry.input_buf[4].genblk1[0].mid ));
 sky130_fd_sc_hd__inv_2 \l_fifo.genblk1[4].entry.input_buf[4].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[4].entry.input_buf[4].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[4].entry.input_buf[4].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[4].entry.input_buf[5].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[4].entry.input_buf[5].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[4].entry.input_buf[5].genblk1[0].mid ));
 sky130_fd_sc_hd__inv_2 \l_fifo.genblk1[4].entry.input_buf[5].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[4].entry.input_buf[5].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[4].entry.input_buf[5].X ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[4].entry.latch[0]  (.D(\l_fifo.genblk1[4].entry.input_buf[0].X ),
    .GATE(\l_fifo.genblk1[4].entry.empty ),
    .RESET_B(net30),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[3].entry.input_buf[0].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[4].entry.latch[1]  (.D(\l_fifo.genblk1[4].entry.input_buf[1].X ),
    .GATE(\l_fifo.genblk1[4].entry.empty ),
    .RESET_B(net30),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[3].entry.input_buf[1].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[4].entry.latch[2]  (.D(\l_fifo.genblk1[4].entry.input_buf[2].X ),
    .GATE(\l_fifo.genblk1[4].entry.empty ),
    .RESET_B(net32),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[3].entry.input_buf[2].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[4].entry.latch[3]  (.D(\l_fifo.genblk1[4].entry.input_buf[3].X ),
    .GATE(\l_fifo.genblk1[4].entry.empty ),
    .RESET_B(net32),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[3].entry.input_buf[3].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[4].entry.latch[4]  (.D(\l_fifo.genblk1[4].entry.input_buf[4].X ),
    .GATE(\l_fifo.genblk1[4].entry.empty ),
    .RESET_B(net30),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[3].entry.input_buf[4].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[4].entry.latch[5]  (.D(\l_fifo.genblk1[4].entry.input_buf[5].X ),
    .GATE(\l_fifo.genblk1[4].entry.empty ),
    .RESET_B(net31),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[3].entry.input_buf[5].A ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[5].entry.input_buf[0].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[5].entry.input_buf[0].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[5].entry.input_buf[0].genblk1[0].mid ));
 sky130_fd_sc_hd__inv_2 \l_fifo.genblk1[5].entry.input_buf[0].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[5].entry.input_buf[0].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[5].entry.input_buf[0].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[5].entry.input_buf[1].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[5].entry.input_buf[1].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[5].entry.input_buf[1].genblk1[0].mid ));
 sky130_fd_sc_hd__inv_2 \l_fifo.genblk1[5].entry.input_buf[1].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[5].entry.input_buf[1].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[5].entry.input_buf[1].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[5].entry.input_buf[2].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[5].entry.input_buf[2].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[5].entry.input_buf[2].genblk1[0].mid ));
 sky130_fd_sc_hd__inv_2 \l_fifo.genblk1[5].entry.input_buf[2].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[5].entry.input_buf[2].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[5].entry.input_buf[2].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[5].entry.input_buf[3].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[5].entry.input_buf[3].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[5].entry.input_buf[3].genblk1[0].mid ));
 sky130_fd_sc_hd__inv_2 \l_fifo.genblk1[5].entry.input_buf[3].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[5].entry.input_buf[3].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[5].entry.input_buf[3].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[5].entry.input_buf[4].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[5].entry.input_buf[4].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[5].entry.input_buf[4].genblk1[0].mid ));
 sky130_fd_sc_hd__inv_2 \l_fifo.genblk1[5].entry.input_buf[4].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[5].entry.input_buf[4].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[5].entry.input_buf[4].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[5].entry.input_buf[5].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[5].entry.input_buf[5].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[5].entry.input_buf[5].genblk1[0].mid ));
 sky130_fd_sc_hd__inv_2 \l_fifo.genblk1[5].entry.input_buf[5].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[5].entry.input_buf[5].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[5].entry.input_buf[5].X ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[5].entry.latch[0]  (.D(\l_fifo.genblk1[5].entry.input_buf[0].X ),
    .GATE(\l_fifo.genblk1[5].entry.empty ),
    .RESET_B(net30),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[4].entry.input_buf[0].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[5].entry.latch[1]  (.D(\l_fifo.genblk1[5].entry.input_buf[1].X ),
    .GATE(\l_fifo.genblk1[5].entry.empty ),
    .RESET_B(net30),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[4].entry.input_buf[1].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[5].entry.latch[2]  (.D(\l_fifo.genblk1[5].entry.input_buf[2].X ),
    .GATE(\l_fifo.genblk1[5].entry.empty ),
    .RESET_B(net30),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[4].entry.input_buf[2].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[5].entry.latch[3]  (.D(\l_fifo.genblk1[5].entry.input_buf[3].X ),
    .GATE(\l_fifo.genblk1[5].entry.empty ),
    .RESET_B(net31),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[4].entry.input_buf[3].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[5].entry.latch[4]  (.D(\l_fifo.genblk1[5].entry.input_buf[4].X ),
    .GATE(\l_fifo.genblk1[5].entry.empty ),
    .RESET_B(net30),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[4].entry.input_buf[4].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[5].entry.latch[5]  (.D(\l_fifo.genblk1[5].entry.input_buf[5].X ),
    .GATE(\l_fifo.genblk1[5].entry.empty ),
    .RESET_B(net31),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[4].entry.input_buf[5].A ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[6].entry.input_buf[0].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[6].entry.input_buf[0].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[6].entry.input_buf[0].genblk1[0].mid ));
 sky130_fd_sc_hd__inv_2 \l_fifo.genblk1[6].entry.input_buf[0].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[6].entry.input_buf[0].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[6].entry.input_buf[0].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[6].entry.input_buf[1].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[6].entry.input_buf[1].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[6].entry.input_buf[1].genblk1[0].mid ));
 sky130_fd_sc_hd__inv_2 \l_fifo.genblk1[6].entry.input_buf[1].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[6].entry.input_buf[1].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[6].entry.input_buf[1].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[6].entry.input_buf[2].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[6].entry.input_buf[2].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[6].entry.input_buf[2].genblk1[0].mid ));
 sky130_fd_sc_hd__inv_2 \l_fifo.genblk1[6].entry.input_buf[2].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[6].entry.input_buf[2].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[6].entry.input_buf[2].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[6].entry.input_buf[3].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[6].entry.input_buf[3].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[6].entry.input_buf[3].genblk1[0].mid ));
 sky130_fd_sc_hd__inv_2 \l_fifo.genblk1[6].entry.input_buf[3].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[6].entry.input_buf[3].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[6].entry.input_buf[3].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[6].entry.input_buf[4].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[6].entry.input_buf[4].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[6].entry.input_buf[4].genblk1[0].mid ));
 sky130_fd_sc_hd__inv_2 \l_fifo.genblk1[6].entry.input_buf[4].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[6].entry.input_buf[4].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[6].entry.input_buf[4].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[6].entry.input_buf[5].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[6].entry.input_buf[5].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[6].entry.input_buf[5].genblk1[0].mid ));
 sky130_fd_sc_hd__inv_2 \l_fifo.genblk1[6].entry.input_buf[5].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[6].entry.input_buf[5].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[6].entry.input_buf[5].X ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[6].entry.latch[0]  (.D(\l_fifo.genblk1[6].entry.input_buf[0].X ),
    .GATE(\l_fifo.genblk1[6].entry.empty ),
    .RESET_B(net24),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[5].entry.input_buf[0].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[6].entry.latch[1]  (.D(\l_fifo.genblk1[6].entry.input_buf[1].X ),
    .GATE(\l_fifo.genblk1[6].entry.empty ),
    .RESET_B(net29),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[5].entry.input_buf[1].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[6].entry.latch[2]  (.D(\l_fifo.genblk1[6].entry.input_buf[2].X ),
    .GATE(\l_fifo.genblk1[6].entry.empty ),
    .RESET_B(net29),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[5].entry.input_buf[2].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[6].entry.latch[3]  (.D(\l_fifo.genblk1[6].entry.input_buf[3].X ),
    .GATE(\l_fifo.genblk1[6].entry.empty ),
    .RESET_B(net29),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[5].entry.input_buf[3].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[6].entry.latch[4]  (.D(\l_fifo.genblk1[6].entry.input_buf[4].X ),
    .GATE(\l_fifo.genblk1[6].entry.empty ),
    .RESET_B(net29),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[5].entry.input_buf[4].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[6].entry.latch[5]  (.D(\l_fifo.genblk1[6].entry.input_buf[5].X ),
    .GATE(\l_fifo.genblk1[6].entry.empty ),
    .RESET_B(net29),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[5].entry.input_buf[5].A ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[7].entry.input_buf[0].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[7].entry.input_buf[0].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[7].entry.input_buf[0].genblk1[0].mid ));
 sky130_fd_sc_hd__inv_2 \l_fifo.genblk1[7].entry.input_buf[0].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[7].entry.input_buf[0].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[7].entry.input_buf[0].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[7].entry.input_buf[1].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[7].entry.input_buf[1].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[7].entry.input_buf[1].genblk1[0].mid ));
 sky130_fd_sc_hd__inv_2 \l_fifo.genblk1[7].entry.input_buf[1].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[7].entry.input_buf[1].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[7].entry.input_buf[1].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[7].entry.input_buf[2].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[7].entry.input_buf[2].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[7].entry.input_buf[2].genblk1[0].mid ));
 sky130_fd_sc_hd__inv_2 \l_fifo.genblk1[7].entry.input_buf[2].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[7].entry.input_buf[2].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[7].entry.input_buf[2].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[7].entry.input_buf[3].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[7].entry.input_buf[3].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[7].entry.input_buf[3].genblk1[0].mid ));
 sky130_fd_sc_hd__clkinv_2 \l_fifo.genblk1[7].entry.input_buf[3].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[7].entry.input_buf[3].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[7].entry.input_buf[3].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[7].entry.input_buf[4].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[7].entry.input_buf[4].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[7].entry.input_buf[4].genblk1[0].mid ));
 sky130_fd_sc_hd__clkinv_2 \l_fifo.genblk1[7].entry.input_buf[4].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[7].entry.input_buf[4].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[7].entry.input_buf[4].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[7].entry.input_buf[5].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[7].entry.input_buf[5].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[7].entry.input_buf[5].genblk1[0].mid ));
 sky130_fd_sc_hd__clkinv_2 \l_fifo.genblk1[7].entry.input_buf[5].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[7].entry.input_buf[5].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[7].entry.input_buf[5].X ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[7].entry.latch[0]  (.D(\l_fifo.genblk1[7].entry.input_buf[0].X ),
    .GATE(\l_fifo.genblk1[7].entry.empty ),
    .RESET_B(net34),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[6].entry.input_buf[0].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[7].entry.latch[1]  (.D(\l_fifo.genblk1[7].entry.input_buf[1].X ),
    .GATE(\l_fifo.genblk1[7].entry.empty ),
    .RESET_B(net34),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[6].entry.input_buf[1].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[7].entry.latch[2]  (.D(\l_fifo.genblk1[7].entry.input_buf[2].X ),
    .GATE(\l_fifo.genblk1[7].entry.empty ),
    .RESET_B(net29),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[6].entry.input_buf[2].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[7].entry.latch[3]  (.D(\l_fifo.genblk1[7].entry.input_buf[3].X ),
    .GATE(\l_fifo.genblk1[7].entry.empty ),
    .RESET_B(net25),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[6].entry.input_buf[3].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[7].entry.latch[4]  (.D(\l_fifo.genblk1[7].entry.input_buf[4].X ),
    .GATE(\l_fifo.genblk1[7].entry.empty ),
    .RESET_B(net34),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[6].entry.input_buf[4].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[7].entry.latch[5]  (.D(\l_fifo.genblk1[7].entry.input_buf[5].X ),
    .GATE(\l_fifo.genblk1[7].entry.empty ),
    .RESET_B(net42),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[6].entry.input_buf[5].A ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[8].entry.input_buf[0].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[8].entry.input_buf[0].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[8].entry.input_buf[0].genblk1[0].mid ));
 sky130_fd_sc_hd__clkinv_2 \l_fifo.genblk1[8].entry.input_buf[0].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[8].entry.input_buf[0].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[8].entry.input_buf[0].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[8].entry.input_buf[1].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[8].entry.input_buf[1].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[8].entry.input_buf[1].genblk1[0].mid ));
 sky130_fd_sc_hd__inv_2 \l_fifo.genblk1[8].entry.input_buf[1].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[8].entry.input_buf[1].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[8].entry.input_buf[1].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[8].entry.input_buf[2].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[8].entry.input_buf[2].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[8].entry.input_buf[2].genblk1[0].mid ));
 sky130_fd_sc_hd__inv_2 \l_fifo.genblk1[8].entry.input_buf[2].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[8].entry.input_buf[2].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[8].entry.input_buf[2].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[8].entry.input_buf[3].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[8].entry.input_buf[3].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[8].entry.input_buf[3].genblk1[0].mid ));
 sky130_fd_sc_hd__inv_2 \l_fifo.genblk1[8].entry.input_buf[3].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[8].entry.input_buf[3].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[8].entry.input_buf[3].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[8].entry.input_buf[4].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[8].entry.input_buf[4].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[8].entry.input_buf[4].genblk1[0].mid ));
 sky130_fd_sc_hd__inv_2 \l_fifo.genblk1[8].entry.input_buf[4].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[8].entry.input_buf[4].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[8].entry.input_buf[4].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[8].entry.input_buf[5].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[8].entry.input_buf[5].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[8].entry.input_buf[5].genblk1[0].mid ));
 sky130_fd_sc_hd__inv_2 \l_fifo.genblk1[8].entry.input_buf[5].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[8].entry.input_buf[5].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[8].entry.input_buf[5].X ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[8].entry.latch[0]  (.D(\l_fifo.genblk1[8].entry.input_buf[0].X ),
    .GATE(\l_fifo.genblk1[8].entry.empty ),
    .RESET_B(net34),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[7].entry.input_buf[0].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[8].entry.latch[1]  (.D(\l_fifo.genblk1[8].entry.input_buf[1].X ),
    .GATE(\l_fifo.genblk1[8].entry.empty ),
    .RESET_B(net34),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[7].entry.input_buf[1].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[8].entry.latch[2]  (.D(\l_fifo.genblk1[8].entry.input_buf[2].X ),
    .GATE(\l_fifo.genblk1[8].entry.empty ),
    .RESET_B(net43),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[7].entry.input_buf[2].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[8].entry.latch[3]  (.D(\l_fifo.genblk1[8].entry.input_buf[3].X ),
    .GATE(\l_fifo.genblk1[8].entry.empty ),
    .RESET_B(net34),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[7].entry.input_buf[3].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[8].entry.latch[4]  (.D(\l_fifo.genblk1[8].entry.input_buf[4].X ),
    .GATE(\l_fifo.genblk1[8].entry.empty ),
    .RESET_B(net34),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[7].entry.input_buf[4].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[8].entry.latch[5]  (.D(\l_fifo.genblk1[8].entry.input_buf[5].X ),
    .GATE(\l_fifo.genblk1[8].entry.empty ),
    .RESET_B(net42),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[7].entry.input_buf[5].A ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[9].entry.input_buf[0].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[9].entry.input_buf[0].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[9].entry.input_buf[0].genblk1[0].mid ));
 sky130_fd_sc_hd__inv_2 \l_fifo.genblk1[9].entry.input_buf[0].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[9].entry.input_buf[0].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[9].entry.input_buf[0].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[9].entry.input_buf[1].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[9].entry.input_buf[1].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[9].entry.input_buf[1].genblk1[0].mid ));
 sky130_fd_sc_hd__clkinv_2 \l_fifo.genblk1[9].entry.input_buf[1].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[9].entry.input_buf[1].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[9].entry.input_buf[1].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[9].entry.input_buf[2].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[9].entry.input_buf[2].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[9].entry.input_buf[2].genblk1[0].mid ));
 sky130_fd_sc_hd__inv_2 \l_fifo.genblk1[9].entry.input_buf[2].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[9].entry.input_buf[2].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[9].entry.input_buf[2].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[9].entry.input_buf[3].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[9].entry.input_buf[3].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[9].entry.input_buf[3].genblk1[0].mid ));
 sky130_fd_sc_hd__inv_2 \l_fifo.genblk1[9].entry.input_buf[3].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[9].entry.input_buf[3].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[9].entry.input_buf[3].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[9].entry.input_buf[4].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[9].entry.input_buf[4].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[9].entry.input_buf[4].genblk1[0].mid ));
 sky130_fd_sc_hd__inv_2 \l_fifo.genblk1[9].entry.input_buf[4].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[9].entry.input_buf[4].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[9].entry.input_buf[4].X ));
 sky130_fd_sc_hd__inv_1 \l_fifo.genblk1[9].entry.input_buf[5].genblk1[0].genblk1.inv_first  (.A(\l_fifo.genblk1[9].entry.input_buf[5].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[9].entry.input_buf[5].genblk1[0].mid ));
 sky130_fd_sc_hd__inv_2 \l_fifo.genblk1[9].entry.input_buf[5].genblk1[0].genblk2.inv_last  (.A(\l_fifo.genblk1[9].entry.input_buf[5].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\l_fifo.genblk1[9].entry.input_buf[5].X ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[9].entry.latch[0]  (.D(\l_fifo.genblk1[9].entry.input_buf[0].X ),
    .GATE(\l_fifo.genblk1[10].entry.next_is_empty ),
    .RESET_B(net42),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[8].entry.input_buf[0].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[9].entry.latch[1]  (.D(\l_fifo.genblk1[9].entry.input_buf[1].X ),
    .GATE(\l_fifo.genblk1[10].entry.next_is_empty ),
    .RESET_B(net42),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[8].entry.input_buf[1].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[9].entry.latch[2]  (.D(\l_fifo.genblk1[9].entry.input_buf[2].X ),
    .GATE(\l_fifo.genblk1[10].entry.next_is_empty ),
    .RESET_B(net43),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[8].entry.input_buf[2].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[9].entry.latch[3]  (.D(\l_fifo.genblk1[9].entry.input_buf[3].X ),
    .GATE(\l_fifo.genblk1[10].entry.next_is_empty ),
    .RESET_B(net43),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[8].entry.input_buf[3].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[9].entry.latch[4]  (.D(\l_fifo.genblk1[9].entry.input_buf[4].X ),
    .GATE(\l_fifo.genblk1[10].entry.next_is_empty ),
    .RESET_B(net35),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[8].entry.input_buf[4].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[9].entry.latch[5]  (.D(\l_fifo.genblk1[9].entry.input_buf[5].X ),
    .GATE(\l_fifo.genblk1[10].entry.next_is_empty ),
    .RESET_B(net25),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[8].entry.input_buf[5].A ));
endmodule
