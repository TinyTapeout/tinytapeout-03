// This is the unpowered netlist.
module scan_controller (clk,
    la_scan_clk_in,
    la_scan_data_in,
    la_scan_data_out,
    la_scan_latch_en,
    la_scan_select,
    ready,
    reset,
    scan_clk_in,
    scan_clk_out,
    scan_data_in,
    scan_data_out,
    scan_latch_en,
    scan_select,
    set_clk_div,
    slow_clk,
    active_select,
    driver_sel,
    inputs,
    oeb,
    outputs);
 input clk;
 input la_scan_clk_in;
 input la_scan_data_in;
 output la_scan_data_out;
 input la_scan_latch_en;
 input la_scan_select;
 output ready;
 input reset;
 input scan_clk_in;
 output scan_clk_out;
 input scan_data_in;
 output scan_data_out;
 output scan_latch_en;
 output scan_select;
 input set_clk_div;
 output slow_clk;
 input [8:0] active_select;
 input [1:0] driver_sel;
 input [7:0] inputs;
 output [37:0] oeb;
 output [7:0] outputs;

 wire net43;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net44;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net45;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _039_;
 wire _041_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire _203_;
 wire _204_;
 wire _205_;
 wire _206_;
 wire _207_;
 wire _208_;
 wire _209_;
 wire _210_;
 wire _211_;
 wire _212_;
 wire _213_;
 wire _214_;
 wire _215_;
 wire _216_;
 wire _217_;
 wire _218_;
 wire _219_;
 wire _220_;
 wire _221_;
 wire _222_;
 wire _223_;
 wire _224_;
 wire _225_;
 wire _226_;
 wire _227_;
 wire _228_;
 wire _229_;
 wire _230_;
 wire _231_;
 wire _232_;
 wire _233_;
 wire _234_;
 wire _235_;
 wire _236_;
 wire _237_;
 wire _238_;
 wire _239_;
 wire _240_;
 wire _241_;
 wire _242_;
 wire _243_;
 wire _244_;
 wire _245_;
 wire _246_;
 wire _247_;
 wire _248_;
 wire _249_;
 wire _250_;
 wire _251_;
 wire _252_;
 wire _253_;
 wire _254_;
 wire _255_;
 wire _256_;
 wire _257_;
 wire _258_;
 wire _259_;
 wire _260_;
 wire _261_;
 wire _262_;
 wire _263_;
 wire _264_;
 wire _265_;
 wire _266_;
 wire _267_;
 wire _268_;
 wire _269_;
 wire _270_;
 wire _271_;
 wire _272_;
 wire _273_;
 wire _274_;
 wire _275_;
 wire _276_;
 wire _277_;
 wire _278_;
 wire _279_;
 wire _280_;
 wire _281_;
 wire _282_;
 wire _283_;
 wire _284_;
 wire _285_;
 wire _286_;
 wire _287_;
 wire _288_;
 wire _289_;
 wire _290_;
 wire _291_;
 wire _292_;
 wire _293_;
 wire _294_;
 wire _295_;
 wire _296_;
 wire _297_;
 wire _298_;
 wire _299_;
 wire _300_;
 wire _301_;
 wire _302_;
 wire _303_;
 wire _304_;
 wire _305_;
 wire _306_;
 wire _307_;
 wire _308_;
 wire _309_;
 wire _310_;
 wire _311_;
 wire _312_;
 wire _313_;
 wire _314_;
 wire _315_;
 wire _316_;
 wire _317_;
 wire _318_;
 wire _319_;
 wire _320_;
 wire _321_;
 wire _322_;
 wire _323_;
 wire _324_;
 wire _325_;
 wire _326_;
 wire _327_;
 wire _328_;
 wire _329_;
 wire _330_;
 wire _331_;
 wire _332_;
 wire _333_;
 wire _334_;
 wire _335_;
 wire _336_;
 wire _337_;
 wire _338_;
 wire _339_;
 wire active;
 wire \aio_input_reg[0] ;
 wire \aio_input_reg[1] ;
 wire \aio_input_reg[2] ;
 wire \aio_input_reg[3] ;
 wire \aio_input_reg[4] ;
 wire \aio_input_reg[5] ;
 wire \aio_input_reg[6] ;
 wire \aio_input_reg[7] ;
 wire aio_input_sh;
 wire \aio_input_shift[0] ;
 wire \aio_input_shift[1] ;
 wire \aio_input_shift[2] ;
 wire \aio_input_shift[3] ;
 wire \aio_input_shift[4] ;
 wire \aio_input_shift[5] ;
 wire \aio_input_shift[6] ;
 wire \aio_input_shift[7] ;
 wire \aio_input_sync[0] ;
 wire \aio_input_sync[1] ;
 wire \aio_input_sync[2] ;
 wire \aio_input_sync[3] ;
 wire \aio_input_sync[4] ;
 wire \aio_input_sync[5] ;
 wire \aio_input_sync[6] ;
 wire \aio_input_sync[7] ;
 wire aio_output_cap;
 wire \aio_output_reg[0] ;
 wire \aio_output_reg[1] ;
 wire \aio_output_reg[2] ;
 wire \aio_output_reg[3] ;
 wire \aio_output_reg[4] ;
 wire \aio_output_reg[5] ;
 wire \aio_output_reg[6] ;
 wire \aio_output_reg[7] ;
 wire \aio_output_shift[0] ;
 wire \aio_output_shift[1] ;
 wire \aio_output_shift[2] ;
 wire \aio_output_shift[3] ;
 wire \aio_output_shift[4] ;
 wire \aio_output_shift[5] ;
 wire \aio_output_shift[6] ;
 wire \aio_output_shift[7] ;
 wire \bit_cnt[0] ;
 wire \bit_cnt[1] ;
 wire \bit_cnt[2] ;
 wire \clk_divider_I.active ;
 wire \clk_divider_I.ce ;
 wire \clk_divider_I.compare[0] ;
 wire \clk_divider_I.compare[1] ;
 wire \clk_divider_I.compare[2] ;
 wire \clk_divider_I.compare[3] ;
 wire \clk_divider_I.compare[4] ;
 wire \clk_divider_I.compare[5] ;
 wire \clk_divider_I.compare[6] ;
 wire \clk_divider_I.compare[7] ;
 wire \clk_divider_I.counter[0] ;
 wire \clk_divider_I.counter[1] ;
 wire \clk_divider_I.counter[2] ;
 wire \clk_divider_I.counter[3] ;
 wire \clk_divider_I.counter[4] ;
 wire \clk_divider_I.counter[5] ;
 wire \clk_divider_I.counter[6] ;
 wire \clk_divider_I.counter[7] ;
 wire \clk_divider_I.reset ;
 wire \clk_divider_I.set_now ;
 wire \clk_divider_I.set_sync[0] ;
 wire \clk_divider_I.set_sync[1] ;
 wire clknet_0_clk;
 wire clknet_0_scan_clk_in;
 wire clknet_1_0__leaf_scan_clk_in;
 wire clknet_1_1__leaf_scan_clk_in;
 wire clknet_3_0__leaf_clk;
 wire clknet_3_1__leaf_clk;
 wire clknet_3_2__leaf_clk;
 wire clknet_3_3__leaf_clk;
 wire clknet_3_4__leaf_clk;
 wire clknet_3_5__leaf_clk;
 wire clknet_3_6__leaf_clk;
 wire clknet_3_7__leaf_clk;
 wire int_scan_clk_out;
 wire int_scan_data_out;
 wire int_scan_latch_en;
 wire int_scan_select;
 wire net1;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net2;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net3;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net4;
 wire net40;
 wire net41;
 wire net42;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net9;
 wire net90;
 wire net91;
 wire \proj_cnt[0] ;
 wire \proj_cnt[1] ;
 wire \proj_cnt[2] ;
 wire \proj_cnt[3] ;
 wire \proj_cnt[4] ;
 wire \proj_cnt[5] ;
 wire \proj_cnt[6] ;
 wire \proj_cnt[7] ;
 wire \proj_cnt[8] ;
 wire \rst_shift[0] ;
 wire \rst_shift[1] ;
 wire \state[0] ;
 wire \state[12] ;
 wire \state[13] ;
 wire \state[1] ;
 wire \state[2] ;
 wire \state[3] ;
 wire \state[4] ;
 wire \state[5] ;
 wire \state[6] ;
 wire \state[8] ;
 wire \state[9] ;
 wire \ws_cfg[0] ;
 wire \ws_cfg[1] ;
 wire \ws_cfg[2] ;
 wire \ws_cfg[3] ;
 wire \ws_cfg[4] ;
 wire \ws_cfg[5] ;
 wire \ws_cfg[6] ;
 wire \ws_cfg[7] ;
 wire \ws_cnt[0] ;
 wire \ws_cnt[1] ;
 wire \ws_cnt[2] ;
 wire \ws_cnt[3] ;
 wire \ws_cnt[4] ;
 wire \ws_cnt[5] ;
 wire \ws_cnt[6] ;
 wire \ws_cnt[7] ;
 wire ws_set_now;
 wire \ws_set_sync[0] ;
 wire \ws_set_sync[1] ;
 wire \ws_set_sync[2] ;

 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(net19));
 sky130_fd_sc_hd__fill_2 FILLER_0_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_202 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_210 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_258 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_398 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_471 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_115 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_173 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_264 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_275 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_292 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_360 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_457 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_59 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_108 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_144 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_164 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_20 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_202 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_286 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_316 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_348 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_411 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_96 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_13 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_186 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_207 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_224 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_26 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_298 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_42 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_457 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_471 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_50 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_96 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_243 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_256 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_344 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_43 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_62 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_154 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_235 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_39 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_56 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_135 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_180 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_192 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_230 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_242 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_256 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_319 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_406 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_95 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_128 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_132 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_176 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_214 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_267 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_288 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_392 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_60 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_124 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_136 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_348 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_403 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_68 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_100 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_392 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_404 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_451 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_144 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_178 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_303 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_403 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_420 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_471 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_64 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_144 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_20 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_32 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_44 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_124 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_192 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_227 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_236 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_428 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_67 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_143 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_151 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_176 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_247 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_308 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_32 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_354 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_425 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_472 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_64 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_154 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_23 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_230 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_300 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_427 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_456 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_471 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_32 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_44 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_471 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_202 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_214 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_471 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_17 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_210 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_266 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_272 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_314 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_322 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_398 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_406 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_42 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_62 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_70 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_76 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_152 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_156 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_215 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_457 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_471 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_207 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_100 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_112 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_152 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_290 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_471 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_96 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_156 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_20 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_248 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_286 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_32 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_351 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_42 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_8 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_99 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_159 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_208 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_471 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_353 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_376 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_48 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_67 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_158 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_202 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_26 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_272 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_176 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_199 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_243 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_295 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_364 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_40 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_410 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_422 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_67 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_93 ();
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_56 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_57 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_58 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_59 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_60 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_61 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_62 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_63 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_64 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_65 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_66 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_67 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_68 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_69 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_70 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_71 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_72 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_73 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_74 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_75 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_76 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_77 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_78 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_79 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_80 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_81 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_82 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_83 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_84 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_85 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_86 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_87 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_88 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_89 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_90 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_91 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_92 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_93 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_94 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_95 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_96 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_97 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_98 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_99 ();
 sky130_fd_sc_hd__xor2_1 _341_ (.A(\clk_divider_I.counter[6] ),
    .B(\clk_divider_I.compare[6] ),
    .X(_126_));
 sky130_fd_sc_hd__xor2_1 _342_ (.A(\clk_divider_I.counter[7] ),
    .B(\clk_divider_I.compare[7] ),
    .X(_127_));
 sky130_fd_sc_hd__xor2_1 _343_ (.A(\clk_divider_I.counter[1] ),
    .B(\clk_divider_I.compare[1] ),
    .X(_128_));
 sky130_fd_sc_hd__xor2_1 _344_ (.A(\clk_divider_I.counter[0] ),
    .B(\clk_divider_I.compare[0] ),
    .X(_129_));
 sky130_fd_sc_hd__or4_1 _345_ (.A(_126_),
    .B(_127_),
    .C(_128_),
    .D(_129_),
    .X(_130_));
 sky130_fd_sc_hd__xor2_1 _346_ (.A(\clk_divider_I.counter[5] ),
    .B(\clk_divider_I.compare[5] ),
    .X(_131_));
 sky130_fd_sc_hd__xor2_1 _347_ (.A(\clk_divider_I.counter[2] ),
    .B(\clk_divider_I.compare[2] ),
    .X(_132_));
 sky130_fd_sc_hd__xor2_1 _348_ (.A(\clk_divider_I.counter[4] ),
    .B(\clk_divider_I.compare[4] ),
    .X(_133_));
 sky130_fd_sc_hd__xor2_1 _349_ (.A(\clk_divider_I.counter[3] ),
    .B(\clk_divider_I.compare[3] ),
    .X(_134_));
 sky130_fd_sc_hd__or4_1 _350_ (.A(_131_),
    .B(_132_),
    .C(_133_),
    .D(_134_),
    .X(_135_));
 sky130_fd_sc_hd__nor2_1 _351_ (.A(_130_),
    .B(_135_),
    .Y(_136_));
 sky130_fd_sc_hd__nand2_2 _352_ (.A(\clk_divider_I.ce ),
    .B(_136_),
    .Y(_137_));
 sky130_fd_sc_hd__xnor2_1 _353_ (.A(net41),
    .B(_137_),
    .Y(_125_));
 sky130_fd_sc_hd__and4_1 _354_ (.A(\clk_divider_I.ce ),
    .B(\clk_divider_I.counter[2] ),
    .C(\clk_divider_I.counter[1] ),
    .D(\clk_divider_I.counter[0] ),
    .X(_138_));
 sky130_fd_sc_hd__and3_1 _355_ (.A(\clk_divider_I.counter[4] ),
    .B(\clk_divider_I.counter[3] ),
    .C(_138_),
    .X(_139_));
 sky130_fd_sc_hd__and3_1 _356_ (.A(\clk_divider_I.counter[6] ),
    .B(\clk_divider_I.counter[5] ),
    .C(_139_),
    .X(_140_));
 sky130_fd_sc_hd__or2_1 _357_ (.A(\clk_divider_I.counter[7] ),
    .B(_140_),
    .X(_141_));
 sky130_fd_sc_hd__nand2_1 _358_ (.A(\clk_divider_I.counter[7] ),
    .B(_140_),
    .Y(_142_));
 sky130_fd_sc_hd__and3_1 _359_ (.A(_137_),
    .B(_141_),
    .C(_142_),
    .X(_143_));
 sky130_fd_sc_hd__clkbuf_1 _360_ (.A(_143_),
    .X(_124_));
 sky130_fd_sc_hd__clkbuf_4 _361_ (.A(\clk_divider_I.ce ),
    .X(_144_));
 sky130_fd_sc_hd__nand2_1 _362_ (.A(\clk_divider_I.counter[5] ),
    .B(_139_),
    .Y(_145_));
 sky130_fd_sc_hd__inv_2 _363_ (.A(\clk_divider_I.counter[6] ),
    .Y(_146_));
 sky130_fd_sc_hd__a221oi_1 _364_ (.A1(_144_),
    .A2(_136_),
    .B1(_145_),
    .B2(_146_),
    .C1(_140_),
    .Y(_123_));
 sky130_fd_sc_hd__or2_1 _365_ (.A(\clk_divider_I.counter[5] ),
    .B(_139_),
    .X(_147_));
 sky130_fd_sc_hd__and3_1 _366_ (.A(_137_),
    .B(_145_),
    .C(_147_),
    .X(_148_));
 sky130_fd_sc_hd__clkbuf_1 _367_ (.A(_148_),
    .X(_122_));
 sky130_fd_sc_hd__clkinv_2 _368_ (.A(_139_),
    .Y(_149_));
 sky130_fd_sc_hd__a21o_1 _369_ (.A1(\clk_divider_I.counter[3] ),
    .A2(_138_),
    .B1(\clk_divider_I.counter[4] ),
    .X(_150_));
 sky130_fd_sc_hd__and3_1 _370_ (.A(_137_),
    .B(_149_),
    .C(_150_),
    .X(_151_));
 sky130_fd_sc_hd__clkbuf_1 _371_ (.A(_151_),
    .X(_121_));
 sky130_fd_sc_hd__nand2_1 _372_ (.A(\clk_divider_I.counter[3] ),
    .B(_138_),
    .Y(_152_));
 sky130_fd_sc_hd__or2_1 _373_ (.A(\clk_divider_I.counter[3] ),
    .B(_138_),
    .X(_153_));
 sky130_fd_sc_hd__and3_1 _374_ (.A(_137_),
    .B(_152_),
    .C(_153_),
    .X(_154_));
 sky130_fd_sc_hd__clkbuf_1 _375_ (.A(_154_),
    .X(_120_));
 sky130_fd_sc_hd__clkinv_2 _376_ (.A(_138_),
    .Y(_155_));
 sky130_fd_sc_hd__a31o_1 _377_ (.A1(\clk_divider_I.ce ),
    .A2(\clk_divider_I.counter[1] ),
    .A3(\clk_divider_I.counter[0] ),
    .B1(\clk_divider_I.counter[2] ),
    .X(_156_));
 sky130_fd_sc_hd__and3_1 _378_ (.A(_137_),
    .B(_155_),
    .C(_156_),
    .X(_157_));
 sky130_fd_sc_hd__clkbuf_1 _379_ (.A(_157_),
    .X(_119_));
 sky130_fd_sc_hd__nand3_1 _380_ (.A(\clk_divider_I.ce ),
    .B(\clk_divider_I.counter[1] ),
    .C(\clk_divider_I.counter[0] ),
    .Y(_158_));
 sky130_fd_sc_hd__a21o_1 _381_ (.A1(\clk_divider_I.ce ),
    .A2(\clk_divider_I.counter[0] ),
    .B1(\clk_divider_I.counter[1] ),
    .X(_159_));
 sky130_fd_sc_hd__and3_1 _382_ (.A(_137_),
    .B(_158_),
    .C(_159_),
    .X(_160_));
 sky130_fd_sc_hd__clkbuf_1 _383_ (.A(_160_),
    .X(_118_));
 sky130_fd_sc_hd__nand2_1 _384_ (.A(\clk_divider_I.ce ),
    .B(\clk_divider_I.counter[0] ),
    .Y(_161_));
 sky130_fd_sc_hd__or2_1 _385_ (.A(\clk_divider_I.ce ),
    .B(\clk_divider_I.counter[0] ),
    .X(_162_));
 sky130_fd_sc_hd__and3_1 _386_ (.A(_137_),
    .B(_161_),
    .C(_162_),
    .X(_163_));
 sky130_fd_sc_hd__clkbuf_1 _387_ (.A(_163_),
    .X(_117_));
 sky130_fd_sc_hd__inv_2 _388_ (.A(net24),
    .Y(_041_));
 sky130_fd_sc_hd__inv_2 _389_ (.A(net24),
    .Y(_039_));
 sky130_fd_sc_hd__inv_2 _390_ (.A(net24),
    .Y(_037_));
 sky130_fd_sc_hd__mux2_1 _391_ (.A0(\ws_cfg[7] ),
    .A1(net19),
    .S(ws_set_now),
    .X(_164_));
 sky130_fd_sc_hd__clkbuf_1 _392_ (.A(_164_),
    .X(_072_));
 sky130_fd_sc_hd__mux2_1 _393_ (.A0(\ws_cfg[6] ),
    .A1(net18),
    .S(ws_set_now),
    .X(_165_));
 sky130_fd_sc_hd__clkbuf_1 _394_ (.A(_165_),
    .X(_071_));
 sky130_fd_sc_hd__mux2_1 _395_ (.A0(\ws_cfg[5] ),
    .A1(net17),
    .S(ws_set_now),
    .X(_166_));
 sky130_fd_sc_hd__clkbuf_1 _396_ (.A(_166_),
    .X(_070_));
 sky130_fd_sc_hd__mux2_1 _397_ (.A0(\ws_cfg[4] ),
    .A1(net16),
    .S(ws_set_now),
    .X(_167_));
 sky130_fd_sc_hd__clkbuf_1 _398_ (.A(_167_),
    .X(_069_));
 sky130_fd_sc_hd__mux2_1 _399_ (.A0(\ws_cfg[3] ),
    .A1(net15),
    .S(ws_set_now),
    .X(_168_));
 sky130_fd_sc_hd__clkbuf_1 _400_ (.A(_168_),
    .X(_068_));
 sky130_fd_sc_hd__mux2_1 _401_ (.A0(\ws_cfg[2] ),
    .A1(net14),
    .S(ws_set_now),
    .X(_169_));
 sky130_fd_sc_hd__clkbuf_1 _402_ (.A(_169_),
    .X(_067_));
 sky130_fd_sc_hd__mux2_1 _403_ (.A0(\ws_cfg[1] ),
    .A1(net13),
    .S(ws_set_now),
    .X(_170_));
 sky130_fd_sc_hd__clkbuf_1 _404_ (.A(_170_),
    .X(_066_));
 sky130_fd_sc_hd__mux2_1 _405_ (.A0(\ws_cfg[0] ),
    .A1(net12),
    .S(ws_set_now),
    .X(_171_));
 sky130_fd_sc_hd__clkbuf_1 _406_ (.A(_171_),
    .X(_065_));
 sky130_fd_sc_hd__inv_2 _407_ (.A(\ws_cnt[0] ),
    .Y(_172_));
 sky130_fd_sc_hd__inv_2 _408_ (.A(\ws_cnt[7] ),
    .Y(_173_));
 sky130_fd_sc_hd__xnor2_1 _409_ (.A(\ws_cfg[5] ),
    .B(\ws_cnt[5] ),
    .Y(_174_));
 sky130_fd_sc_hd__o221a_1 _410_ (.A1(\ws_cfg[0] ),
    .A2(_172_),
    .B1(_173_),
    .B2(\ws_cfg[7] ),
    .C1(_174_),
    .X(_175_));
 sky130_fd_sc_hd__inv_2 _411_ (.A(\ws_cfg[6] ),
    .Y(_176_));
 sky130_fd_sc_hd__a22o_1 _412_ (.A1(\ws_cfg[0] ),
    .A2(_172_),
    .B1(\ws_cnt[6] ),
    .B2(_176_),
    .X(_177_));
 sky130_fd_sc_hd__o2bb2a_1 _413_ (.A1_N(\ws_cfg[7] ),
    .A2_N(_173_),
    .B1(_176_),
    .B2(\ws_cnt[6] ),
    .X(_178_));
 sky130_fd_sc_hd__nand2_1 _414_ (.A(\ws_cfg[4] ),
    .B(\ws_cnt[4] ),
    .Y(_179_));
 sky130_fd_sc_hd__or2_1 _415_ (.A(\ws_cfg[4] ),
    .B(\ws_cnt[4] ),
    .X(_180_));
 sky130_fd_sc_hd__xor2_1 _416_ (.A(\ws_cfg[1] ),
    .B(\ws_cnt[1] ),
    .X(_181_));
 sky130_fd_sc_hd__a21oi_1 _417_ (.A1(_179_),
    .A2(_180_),
    .B1(_181_),
    .Y(_182_));
 sky130_fd_sc_hd__nand2_1 _418_ (.A(\ws_cfg[2] ),
    .B(\ws_cnt[2] ),
    .Y(_183_));
 sky130_fd_sc_hd__or2_1 _419_ (.A(\ws_cfg[2] ),
    .B(\ws_cnt[2] ),
    .X(_184_));
 sky130_fd_sc_hd__xor2_1 _420_ (.A(\ws_cfg[3] ),
    .B(\ws_cnt[3] ),
    .X(_185_));
 sky130_fd_sc_hd__a21oi_1 _421_ (.A1(_183_),
    .A2(_184_),
    .B1(_185_),
    .Y(_186_));
 sky130_fd_sc_hd__and4b_1 _422_ (.A_N(_177_),
    .B(_178_),
    .C(_182_),
    .D(_186_),
    .X(_187_));
 sky130_fd_sc_hd__and2_1 _423_ (.A(_175_),
    .B(_187_),
    .X(_188_));
 sky130_fd_sc_hd__mux2_1 _424_ (.A0(\state[8] ),
    .A1(\state[1] ),
    .S(_188_),
    .X(_189_));
 sky130_fd_sc_hd__clkbuf_1 _425_ (.A(_189_),
    .X(_056_));
 sky130_fd_sc_hd__nand2_1 _426_ (.A(_175_),
    .B(_187_),
    .Y(_190_));
 sky130_fd_sc_hd__a21o_1 _427_ (.A1(\state[1] ),
    .A2(_190_),
    .B1(\state[13] ),
    .X(_008_));
 sky130_fd_sc_hd__and2_1 _428_ (.A(\proj_cnt[5] ),
    .B(\proj_cnt[4] ),
    .X(_191_));
 sky130_fd_sc_hd__inv_2 _429_ (.A(\proj_cnt[8] ),
    .Y(_192_));
 sky130_fd_sc_hd__and4_1 _430_ (.A(_192_),
    .B(\proj_cnt[7] ),
    .C(\proj_cnt[6] ),
    .D(\proj_cnt[3] ),
    .X(_193_));
 sky130_fd_sc_hd__nand2_1 _431_ (.A(_191_),
    .B(_193_),
    .Y(_194_));
 sky130_fd_sc_hd__nand3_1 _432_ (.A(\bit_cnt[2] ),
    .B(\bit_cnt[1] ),
    .C(\bit_cnt[0] ),
    .Y(_195_));
 sky130_fd_sc_hd__or4b_1 _433_ (.A(\proj_cnt[2] ),
    .B(\proj_cnt[0] ),
    .C(_195_),
    .D_N(\proj_cnt[1] ),
    .X(_196_));
 sky130_fd_sc_hd__or2_1 _434_ (.A(_194_),
    .B(_196_),
    .X(_197_));
 sky130_fd_sc_hd__a22o_1 _435_ (.A1(\state[8] ),
    .A2(_188_),
    .B1(_197_),
    .B2(\state[12] ),
    .X(_012_));
 sky130_fd_sc_hd__a21o_1 _436_ (.A1(\state[6] ),
    .A2(_190_),
    .B1(\state[9] ),
    .X(_013_));
 sky130_fd_sc_hd__clkbuf_4 _437_ (.A(aio_input_sh),
    .X(_198_));
 sky130_fd_sc_hd__inv_2 _438_ (.A(net1),
    .Y(_199_));
 sky130_fd_sc_hd__inv_2 _439_ (.A(net3),
    .Y(_200_));
 sky130_fd_sc_hd__inv_2 _440_ (.A(net4),
    .Y(_201_));
 sky130_fd_sc_hd__nor2_1 _441_ (.A(\proj_cnt[3] ),
    .B(_201_),
    .Y(_202_));
 sky130_fd_sc_hd__a221o_1 _442_ (.A1(\proj_cnt[0] ),
    .A2(_199_),
    .B1(_200_),
    .B2(\proj_cnt[2] ),
    .C1(_202_),
    .X(_203_));
 sky130_fd_sc_hd__inv_2 _443_ (.A(\proj_cnt[6] ),
    .Y(_204_));
 sky130_fd_sc_hd__o22a_1 _444_ (.A1(\proj_cnt[2] ),
    .A2(_200_),
    .B1(net7),
    .B2(_204_),
    .X(_205_));
 sky130_fd_sc_hd__or2_1 _445_ (.A(\proj_cnt[7] ),
    .B(net8),
    .X(_206_));
 sky130_fd_sc_hd__nand2_1 _446_ (.A(\proj_cnt[7] ),
    .B(net8),
    .Y(_207_));
 sky130_fd_sc_hd__or2_1 _447_ (.A(\proj_cnt[1] ),
    .B(net2),
    .X(_208_));
 sky130_fd_sc_hd__nand2_1 _448_ (.A(\proj_cnt[1] ),
    .B(net2),
    .Y(_209_));
 sky130_fd_sc_hd__a22o_1 _449_ (.A1(_206_),
    .A2(_207_),
    .B1(_208_),
    .B2(_209_),
    .X(_210_));
 sky130_fd_sc_hd__a221o_1 _450_ (.A1(\proj_cnt[3] ),
    .A2(_201_),
    .B1(net7),
    .B2(_204_),
    .C1(_195_),
    .X(_211_));
 sky130_fd_sc_hd__inv_2 _451_ (.A(net6),
    .Y(_212_));
 sky130_fd_sc_hd__xor2_1 _452_ (.A(\proj_cnt[4] ),
    .B(net5),
    .X(_213_));
 sky130_fd_sc_hd__a221o_1 _453_ (.A1(\proj_cnt[5] ),
    .A2(_212_),
    .B1(net9),
    .B2(_192_),
    .C1(_213_),
    .X(_214_));
 sky130_fd_sc_hd__or2b_1 _454_ (.A(net9),
    .B_N(\proj_cnt[8] ),
    .X(_215_));
 sky130_fd_sc_hd__o221a_1 _455_ (.A1(\proj_cnt[0] ),
    .A2(_199_),
    .B1(_212_),
    .B2(\proj_cnt[5] ),
    .C1(_215_),
    .X(_216_));
 sky130_fd_sc_hd__nor4b_1 _456_ (.A(_210_),
    .B(_211_),
    .C(_214_),
    .D_N(_216_),
    .Y(_217_));
 sky130_fd_sc_hd__nand3b_1 _457_ (.A_N(_203_),
    .B(_205_),
    .C(_217_),
    .Y(_218_));
 sky130_fd_sc_hd__a21o_1 _458_ (.A1(_198_),
    .A2(_218_),
    .B1(_144_),
    .X(_011_));
 sky130_fd_sc_hd__clkinv_2 _459_ (.A(_198_),
    .Y(_219_));
 sky130_fd_sc_hd__a2bb2o_1 _460_ (.A1_N(_219_),
    .A2_N(_218_),
    .B1(_190_),
    .B2(\state[2] ),
    .X(_009_));
 sky130_fd_sc_hd__clkinv_2 _461_ (.A(\state[12] ),
    .Y(_220_));
 sky130_fd_sc_hd__a2bb2o_1 _462_ (.A1_N(_220_),
    .A2_N(_197_),
    .B1(_190_),
    .B2(\state[3] ),
    .X(_010_));
 sky130_fd_sc_hd__buf_2 _463_ (.A(\state[0] ),
    .X(_221_));
 sky130_fd_sc_hd__inv_2 _464_ (.A(active),
    .Y(_222_));
 sky130_fd_sc_hd__a21o_1 _465_ (.A1(_221_),
    .A2(_222_),
    .B1(aio_output_cap),
    .X(_007_));
 sky130_fd_sc_hd__clkbuf_2 _466_ (.A(net11),
    .X(_223_));
 sky130_fd_sc_hd__and2_1 _467_ (.A(_223_),
    .B(net10),
    .X(_224_));
 sky130_fd_sc_hd__clkbuf_1 _468_ (.A(_224_),
    .X(_003_));
 sky130_fd_sc_hd__clkbuf_4 _469_ (.A(net11),
    .X(_225_));
 sky130_fd_sc_hd__mux2_2 _470_ (.A0(clknet_1_1__leaf_scan_clk_in),
    .A1(\aio_output_reg[0] ),
    .S(_225_),
    .X(_226_));
 sky130_fd_sc_hd__buf_1 _471_ (.A(_226_),
    .X(net28));
 sky130_fd_sc_hd__mux2_1 _472_ (.A0(net25),
    .A1(\aio_output_reg[1] ),
    .S(_225_),
    .X(_227_));
 sky130_fd_sc_hd__clkbuf_1 _473_ (.A(_227_),
    .X(net29));
 sky130_fd_sc_hd__and2_1 _474_ (.A(_223_),
    .B(\aio_output_reg[2] ),
    .X(_228_));
 sky130_fd_sc_hd__clkbuf_1 _475_ (.A(_228_),
    .X(net30));
 sky130_fd_sc_hd__and2_1 _476_ (.A(_223_),
    .B(\aio_output_reg[3] ),
    .X(_229_));
 sky130_fd_sc_hd__clkbuf_1 _477_ (.A(_229_),
    .X(net31));
 sky130_fd_sc_hd__and2_1 _478_ (.A(_223_),
    .B(\aio_output_reg[4] ),
    .X(_230_));
 sky130_fd_sc_hd__clkbuf_1 _479_ (.A(_230_),
    .X(net32));
 sky130_fd_sc_hd__and2_1 _480_ (.A(_223_),
    .B(\aio_output_reg[5] ),
    .X(_231_));
 sky130_fd_sc_hd__clkbuf_1 _481_ (.A(_231_),
    .X(net33));
 sky130_fd_sc_hd__and2_1 _482_ (.A(_223_),
    .B(\aio_output_reg[6] ),
    .X(_232_));
 sky130_fd_sc_hd__clkbuf_1 _483_ (.A(_232_),
    .X(net34));
 sky130_fd_sc_hd__and2_1 _484_ (.A(_223_),
    .B(\aio_output_reg[7] ),
    .X(_233_));
 sky130_fd_sc_hd__clkbuf_1 _485_ (.A(_233_),
    .X(net35));
 sky130_fd_sc_hd__mux2_1 _486_ (.A0(net12),
    .A1(net20),
    .S(net10),
    .X(_234_));
 sky130_fd_sc_hd__mux2_1 _487_ (.A0(_234_),
    .A1(int_scan_clk_out),
    .S(_225_),
    .X(_235_));
 sky130_fd_sc_hd__clkbuf_1 _488_ (.A(_235_),
    .X(net37));
 sky130_fd_sc_hd__mux2_1 _489_ (.A0(net13),
    .A1(net21),
    .S(net10),
    .X(_236_));
 sky130_fd_sc_hd__mux2_1 _490_ (.A0(_236_),
    .A1(int_scan_data_out),
    .S(_225_),
    .X(_237_));
 sky130_fd_sc_hd__clkbuf_1 _491_ (.A(_237_),
    .X(net38));
 sky130_fd_sc_hd__mux2_1 _492_ (.A0(net14),
    .A1(net23),
    .S(net10),
    .X(_238_));
 sky130_fd_sc_hd__mux2_1 _493_ (.A0(_238_),
    .A1(int_scan_select),
    .S(_225_),
    .X(_239_));
 sky130_fd_sc_hd__clkbuf_1 _494_ (.A(_239_),
    .X(net40));
 sky130_fd_sc_hd__mux2_1 _495_ (.A0(net15),
    .A1(net22),
    .S(net10),
    .X(_240_));
 sky130_fd_sc_hd__mux2_1 _496_ (.A0(_240_),
    .A1(int_scan_latch_en),
    .S(net11),
    .X(_241_));
 sky130_fd_sc_hd__clkbuf_1 _497_ (.A(_241_),
    .X(net39));
 sky130_fd_sc_hd__and3_1 _498_ (.A(\state[3] ),
    .B(_175_),
    .C(_187_),
    .X(_242_));
 sky130_fd_sc_hd__clkbuf_1 _499_ (.A(_242_),
    .X(_005_));
 sky130_fd_sc_hd__and3_1 _500_ (.A(\state[2] ),
    .B(_175_),
    .C(_187_),
    .X(_243_));
 sky130_fd_sc_hd__clkbuf_1 _501_ (.A(_243_),
    .X(_004_));
 sky130_fd_sc_hd__and2_1 _502_ (.A(\state[0] ),
    .B(active),
    .X(_244_));
 sky130_fd_sc_hd__clkbuf_1 _503_ (.A(_244_),
    .X(net36));
 sky130_fd_sc_hd__and3_1 _504_ (.A(\state[6] ),
    .B(_175_),
    .C(_187_),
    .X(_245_));
 sky130_fd_sc_hd__clkbuf_1 _505_ (.A(_245_),
    .X(_006_));
 sky130_fd_sc_hd__or3_1 _506_ (.A(\state[13] ),
    .B(\state[12] ),
    .C(_198_),
    .X(_246_));
 sky130_fd_sc_hd__clkbuf_1 _507_ (.A(_246_),
    .X(_000_));
 sky130_fd_sc_hd__or3_1 _508_ (.A(\state[1] ),
    .B(\state[13] ),
    .C(\state[6] ),
    .X(_247_));
 sky130_fd_sc_hd__clkbuf_1 _509_ (.A(_247_),
    .X(_001_));
 sky130_fd_sc_hd__and2b_1 _510_ (.A_N(\ws_set_sync[2] ),
    .B(\ws_set_sync[1] ),
    .X(_248_));
 sky130_fd_sc_hd__clkbuf_1 _511_ (.A(_248_),
    .X(_002_));
 sky130_fd_sc_hd__and2b_1 _512_ (.A_N(\clk_divider_I.active ),
    .B(\clk_divider_I.set_sync[1] ),
    .X(_249_));
 sky130_fd_sc_hd__clkbuf_1 _513_ (.A(_249_),
    .X(_014_));
 sky130_fd_sc_hd__clkbuf_4 _514_ (.A(\clk_divider_I.reset ),
    .X(_250_));
 sky130_fd_sc_hd__buf_4 _515_ (.A(_250_),
    .X(_251_));
 sky130_fd_sc_hd__inv_2 _516_ (.A(_251_),
    .Y(_015_));
 sky130_fd_sc_hd__mux2_1 _517_ (.A0(\aio_input_shift[1] ),
    .A1(\aio_input_shift[0] ),
    .S(_198_),
    .X(_252_));
 sky130_fd_sc_hd__mux2_1 _518_ (.A0(_252_),
    .A1(\aio_input_reg[1] ),
    .S(_144_),
    .X(_253_));
 sky130_fd_sc_hd__clkbuf_1 _519_ (.A(_253_),
    .X(_057_));
 sky130_fd_sc_hd__mux2_1 _520_ (.A0(\aio_input_shift[2] ),
    .A1(\aio_input_shift[1] ),
    .S(_198_),
    .X(_254_));
 sky130_fd_sc_hd__mux2_1 _521_ (.A0(_254_),
    .A1(\aio_input_reg[2] ),
    .S(_144_),
    .X(_255_));
 sky130_fd_sc_hd__clkbuf_1 _522_ (.A(_255_),
    .X(_058_));
 sky130_fd_sc_hd__mux2_1 _523_ (.A0(\aio_input_shift[3] ),
    .A1(\aio_input_shift[2] ),
    .S(_198_),
    .X(_256_));
 sky130_fd_sc_hd__mux2_1 _524_ (.A0(_256_),
    .A1(\aio_input_reg[3] ),
    .S(_144_),
    .X(_257_));
 sky130_fd_sc_hd__clkbuf_1 _525_ (.A(_257_),
    .X(_059_));
 sky130_fd_sc_hd__mux2_1 _526_ (.A0(\aio_input_shift[4] ),
    .A1(\aio_input_shift[3] ),
    .S(_198_),
    .X(_258_));
 sky130_fd_sc_hd__mux2_1 _527_ (.A0(_258_),
    .A1(\aio_input_reg[4] ),
    .S(_144_),
    .X(_259_));
 sky130_fd_sc_hd__clkbuf_1 _528_ (.A(_259_),
    .X(_060_));
 sky130_fd_sc_hd__mux2_1 _529_ (.A0(\aio_input_shift[5] ),
    .A1(\aio_input_shift[4] ),
    .S(_198_),
    .X(_260_));
 sky130_fd_sc_hd__mux2_1 _530_ (.A0(_260_),
    .A1(\aio_input_reg[5] ),
    .S(_144_),
    .X(_261_));
 sky130_fd_sc_hd__clkbuf_1 _531_ (.A(_261_),
    .X(_061_));
 sky130_fd_sc_hd__mux2_1 _532_ (.A0(\aio_input_shift[6] ),
    .A1(\aio_input_shift[5] ),
    .S(aio_input_sh),
    .X(_262_));
 sky130_fd_sc_hd__mux2_1 _533_ (.A0(_262_),
    .A1(\aio_input_reg[6] ),
    .S(_144_),
    .X(_263_));
 sky130_fd_sc_hd__clkbuf_1 _534_ (.A(_263_),
    .X(_062_));
 sky130_fd_sc_hd__mux2_1 _535_ (.A0(\aio_input_shift[7] ),
    .A1(\aio_input_shift[6] ),
    .S(aio_input_sh),
    .X(_264_));
 sky130_fd_sc_hd__mux2_1 _536_ (.A0(_264_),
    .A1(\aio_input_reg[7] ),
    .S(\clk_divider_I.ce ),
    .X(_265_));
 sky130_fd_sc_hd__clkbuf_1 _537_ (.A(_265_),
    .X(_063_));
 sky130_fd_sc_hd__inv_2 _538_ (.A(_251_),
    .Y(_016_));
 sky130_fd_sc_hd__inv_2 _539_ (.A(_251_),
    .Y(_017_));
 sky130_fd_sc_hd__inv_2 _540_ (.A(_251_),
    .Y(_018_));
 sky130_fd_sc_hd__inv_2 _541_ (.A(_251_),
    .Y(_019_));
 sky130_fd_sc_hd__inv_2 _542_ (.A(_251_),
    .Y(_020_));
 sky130_fd_sc_hd__inv_2 _543_ (.A(_251_),
    .Y(_021_));
 sky130_fd_sc_hd__inv_2 _544_ (.A(_251_),
    .Y(_022_));
 sky130_fd_sc_hd__inv_2 _545_ (.A(_251_),
    .Y(_023_));
 sky130_fd_sc_hd__inv_2 _546_ (.A(_251_),
    .Y(_024_));
 sky130_fd_sc_hd__buf_4 _547_ (.A(_250_),
    .X(_266_));
 sky130_fd_sc_hd__inv_2 _548_ (.A(_266_),
    .Y(_025_));
 sky130_fd_sc_hd__inv_2 _549_ (.A(_266_),
    .Y(_026_));
 sky130_fd_sc_hd__inv_2 _550_ (.A(_266_),
    .Y(_027_));
 sky130_fd_sc_hd__inv_2 _551_ (.A(_266_),
    .Y(_028_));
 sky130_fd_sc_hd__nor2_1 _552_ (.A(_144_),
    .B(_198_),
    .Y(_267_));
 sky130_fd_sc_hd__mux2_1 _553_ (.A0(\aio_input_reg[0] ),
    .A1(net41),
    .S(\clk_divider_I.active ),
    .X(_268_));
 sky130_fd_sc_hd__a22o_1 _554_ (.A1(\aio_input_shift[0] ),
    .A2(_267_),
    .B1(_268_),
    .B2(_144_),
    .X(_064_));
 sky130_fd_sc_hd__inv_2 _555_ (.A(_266_),
    .Y(_029_));
 sky130_fd_sc_hd__inv_2 _556_ (.A(_266_),
    .Y(_030_));
 sky130_fd_sc_hd__inv_2 _557_ (.A(_266_),
    .Y(_031_));
 sky130_fd_sc_hd__inv_2 _558_ (.A(_266_),
    .Y(_032_));
 sky130_fd_sc_hd__inv_2 _559_ (.A(_266_),
    .Y(_033_));
 sky130_fd_sc_hd__inv_2 _560_ (.A(_266_),
    .Y(_034_));
 sky130_fd_sc_hd__buf_4 _561_ (.A(_250_),
    .X(_269_));
 sky130_fd_sc_hd__inv_2 _562_ (.A(_269_),
    .Y(_035_));
 sky130_fd_sc_hd__inv_2 _563_ (.A(_269_),
    .Y(_036_));
 sky130_fd_sc_hd__inv_2 _564__1 (.A(clknet_3_1__leaf_clk),
    .Y(net81));
 sky130_fd_sc_hd__inv_2 _565__2 (.A(clknet_3_1__leaf_clk),
    .Y(net82));
 sky130_fd_sc_hd__inv_2 _566__3 (.A(clknet_3_1__leaf_clk),
    .Y(net83));
 sky130_fd_sc_hd__mux2_1 _567_ (.A0(\clk_divider_I.compare[0] ),
    .A1(net12),
    .S(\clk_divider_I.set_now ),
    .X(_270_));
 sky130_fd_sc_hd__clkbuf_1 _568_ (.A(_270_),
    .X(_073_));
 sky130_fd_sc_hd__mux2_1 _569_ (.A0(\clk_divider_I.compare[1] ),
    .A1(net13),
    .S(\clk_divider_I.set_now ),
    .X(_271_));
 sky130_fd_sc_hd__clkbuf_1 _570_ (.A(_271_),
    .X(_074_));
 sky130_fd_sc_hd__mux2_1 _571_ (.A0(\clk_divider_I.compare[2] ),
    .A1(net14),
    .S(\clk_divider_I.set_now ),
    .X(_272_));
 sky130_fd_sc_hd__clkbuf_1 _572_ (.A(_272_),
    .X(_075_));
 sky130_fd_sc_hd__mux2_1 _573_ (.A0(\clk_divider_I.compare[3] ),
    .A1(net15),
    .S(\clk_divider_I.set_now ),
    .X(_273_));
 sky130_fd_sc_hd__clkbuf_1 _574_ (.A(_273_),
    .X(_076_));
 sky130_fd_sc_hd__mux2_1 _575_ (.A0(\clk_divider_I.compare[4] ),
    .A1(net16),
    .S(\clk_divider_I.set_now ),
    .X(_274_));
 sky130_fd_sc_hd__clkbuf_1 _576_ (.A(_274_),
    .X(_077_));
 sky130_fd_sc_hd__mux2_1 _577_ (.A0(\clk_divider_I.compare[5] ),
    .A1(net17),
    .S(\clk_divider_I.set_now ),
    .X(_275_));
 sky130_fd_sc_hd__clkbuf_1 _578_ (.A(_275_),
    .X(_078_));
 sky130_fd_sc_hd__mux2_1 _579_ (.A0(\clk_divider_I.compare[6] ),
    .A1(net18),
    .S(\clk_divider_I.set_now ),
    .X(_276_));
 sky130_fd_sc_hd__clkbuf_1 _580_ (.A(_276_),
    .X(_079_));
 sky130_fd_sc_hd__mux2_1 _581_ (.A0(\clk_divider_I.compare[7] ),
    .A1(net19),
    .S(\clk_divider_I.set_now ),
    .X(_277_));
 sky130_fd_sc_hd__clkbuf_1 _582_ (.A(_277_),
    .X(_080_));
 sky130_fd_sc_hd__inv_2 _583_ (.A(_269_),
    .Y(_043_));
 sky130_fd_sc_hd__o21a_1 _584_ (.A1(\state[12] ),
    .A2(aio_input_sh),
    .B1(\bit_cnt[0] ),
    .X(_278_));
 sky130_fd_sc_hd__nor2_1 _585_ (.A(\state[0] ),
    .B(_278_),
    .Y(_279_));
 sky130_fd_sc_hd__o31a_1 _586_ (.A1(\bit_cnt[0] ),
    .A2(\state[12] ),
    .A3(_198_),
    .B1(_279_),
    .X(_081_));
 sky130_fd_sc_hd__and2_1 _587_ (.A(\bit_cnt[1] ),
    .B(_278_),
    .X(_280_));
 sky130_fd_sc_hd__nor2_1 _588_ (.A(_221_),
    .B(_280_),
    .Y(_281_));
 sky130_fd_sc_hd__o21a_1 _589_ (.A1(\bit_cnt[1] ),
    .A2(_278_),
    .B1(_281_),
    .X(_082_));
 sky130_fd_sc_hd__o2111a_1 _590_ (.A1(\state[12] ),
    .A2(aio_input_sh),
    .B1(\bit_cnt[2] ),
    .C1(\bit_cnt[1] ),
    .D1(\bit_cnt[0] ),
    .X(_282_));
 sky130_fd_sc_hd__nor2_1 _591_ (.A(_221_),
    .B(_282_),
    .Y(_283_));
 sky130_fd_sc_hd__o21a_1 _592_ (.A1(\bit_cnt[2] ),
    .A2(_280_),
    .B1(_283_),
    .X(_083_));
 sky130_fd_sc_hd__and2_1 _593_ (.A(\proj_cnt[0] ),
    .B(_282_),
    .X(_284_));
 sky130_fd_sc_hd__nor2_1 _594_ (.A(_221_),
    .B(_284_),
    .Y(_285_));
 sky130_fd_sc_hd__o21a_1 _595_ (.A1(\proj_cnt[0] ),
    .A2(_282_),
    .B1(_285_),
    .X(_084_));
 sky130_fd_sc_hd__and2_1 _596_ (.A(\proj_cnt[1] ),
    .B(\proj_cnt[0] ),
    .X(_286_));
 sky130_fd_sc_hd__and2_1 _597_ (.A(_282_),
    .B(_286_),
    .X(_287_));
 sky130_fd_sc_hd__nor2_1 _598_ (.A(_221_),
    .B(_287_),
    .Y(_288_));
 sky130_fd_sc_hd__o21a_1 _599_ (.A1(\proj_cnt[1] ),
    .A2(_284_),
    .B1(_288_),
    .X(_085_));
 sky130_fd_sc_hd__and3_1 _600_ (.A(\proj_cnt[2] ),
    .B(_282_),
    .C(_286_),
    .X(_289_));
 sky130_fd_sc_hd__nor2_1 _601_ (.A(_221_),
    .B(_289_),
    .Y(_290_));
 sky130_fd_sc_hd__o21a_1 _602_ (.A1(\proj_cnt[2] ),
    .A2(_287_),
    .B1(_290_),
    .X(_086_));
 sky130_fd_sc_hd__and4_1 _603_ (.A(\proj_cnt[3] ),
    .B(\proj_cnt[2] ),
    .C(_282_),
    .D(_286_),
    .X(_291_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _604_ (.A(_291_),
    .X(_292_));
 sky130_fd_sc_hd__nor2_1 _605_ (.A(_221_),
    .B(_292_),
    .Y(_293_));
 sky130_fd_sc_hd__o21a_1 _606_ (.A1(\proj_cnt[3] ),
    .A2(_289_),
    .B1(_293_),
    .X(_087_));
 sky130_fd_sc_hd__and2_1 _607_ (.A(\proj_cnt[4] ),
    .B(_292_),
    .X(_294_));
 sky130_fd_sc_hd__nor2_1 _608_ (.A(\state[0] ),
    .B(_294_),
    .Y(_295_));
 sky130_fd_sc_hd__o21a_1 _609_ (.A1(\proj_cnt[4] ),
    .A2(_292_),
    .B1(_295_),
    .X(_088_));
 sky130_fd_sc_hd__a21oi_1 _610_ (.A1(_191_),
    .A2(_292_),
    .B1(_221_),
    .Y(_296_));
 sky130_fd_sc_hd__o21a_1 _611_ (.A1(\proj_cnt[5] ),
    .A2(_294_),
    .B1(_296_),
    .X(_089_));
 sky130_fd_sc_hd__a21oi_1 _612_ (.A1(_191_),
    .A2(_292_),
    .B1(\proj_cnt[6] ),
    .Y(_297_));
 sky130_fd_sc_hd__and3_1 _613_ (.A(\proj_cnt[6] ),
    .B(_191_),
    .C(_292_),
    .X(_298_));
 sky130_fd_sc_hd__nor3_1 _614_ (.A(_221_),
    .B(_297_),
    .C(_298_),
    .Y(_090_));
 sky130_fd_sc_hd__a21oi_1 _615_ (.A1(\proj_cnt[7] ),
    .A2(_298_),
    .B1(_221_),
    .Y(_299_));
 sky130_fd_sc_hd__o21a_1 _616_ (.A1(\proj_cnt[7] ),
    .A2(_298_),
    .B1(_299_),
    .X(_091_));
 sky130_fd_sc_hd__a21oi_1 _617_ (.A1(\proj_cnt[7] ),
    .A2(_298_),
    .B1(\proj_cnt[8] ),
    .Y(_300_));
 sky130_fd_sc_hd__a31o_1 _618_ (.A1(\proj_cnt[8] ),
    .A2(\proj_cnt[7] ),
    .A3(_298_),
    .B1(\state[0] ),
    .X(_301_));
 sky130_fd_sc_hd__nor2_1 _619_ (.A(_300_),
    .B(_301_),
    .Y(_092_));
 sky130_fd_sc_hd__and2_1 _620_ (.A(_223_),
    .B(\aio_input_sync[0] ),
    .X(_302_));
 sky130_fd_sc_hd__clkbuf_1 _621_ (.A(_302_),
    .X(_093_));
 sky130_fd_sc_hd__and2_1 _622_ (.A(_223_),
    .B(\aio_input_sync[1] ),
    .X(_303_));
 sky130_fd_sc_hd__clkbuf_1 _623_ (.A(_303_),
    .X(_094_));
 sky130_fd_sc_hd__and2_1 _624_ (.A(_223_),
    .B(\aio_input_sync[2] ),
    .X(_304_));
 sky130_fd_sc_hd__clkbuf_1 _625_ (.A(_304_),
    .X(_095_));
 sky130_fd_sc_hd__and2_1 _626_ (.A(_225_),
    .B(\aio_input_sync[3] ),
    .X(_305_));
 sky130_fd_sc_hd__clkbuf_1 _627_ (.A(_305_),
    .X(_096_));
 sky130_fd_sc_hd__and2_1 _628_ (.A(_225_),
    .B(\aio_input_sync[4] ),
    .X(_306_));
 sky130_fd_sc_hd__clkbuf_1 _629_ (.A(_306_),
    .X(_097_));
 sky130_fd_sc_hd__and2_1 _630_ (.A(_225_),
    .B(\aio_input_sync[5] ),
    .X(_307_));
 sky130_fd_sc_hd__clkbuf_1 _631_ (.A(_307_),
    .X(_098_));
 sky130_fd_sc_hd__and2_1 _632_ (.A(_225_),
    .B(\aio_input_sync[6] ),
    .X(_308_));
 sky130_fd_sc_hd__clkbuf_1 _633_ (.A(_308_),
    .X(_099_));
 sky130_fd_sc_hd__and2_1 _634_ (.A(_225_),
    .B(\aio_input_sync[7] ),
    .X(_309_));
 sky130_fd_sc_hd__clkbuf_1 _635_ (.A(_309_),
    .X(_100_));
 sky130_fd_sc_hd__mux2_1 _636_ (.A0(\aio_output_reg[0] ),
    .A1(net86),
    .S(aio_output_cap),
    .X(_310_));
 sky130_fd_sc_hd__clkbuf_1 _637_ (.A(_310_),
    .X(_101_));
 sky130_fd_sc_hd__mux2_1 _638_ (.A0(\aio_output_reg[1] ),
    .A1(net90),
    .S(aio_output_cap),
    .X(_311_));
 sky130_fd_sc_hd__clkbuf_1 _639_ (.A(_311_),
    .X(_102_));
 sky130_fd_sc_hd__mux2_1 _640_ (.A0(\aio_output_reg[2] ),
    .A1(net87),
    .S(aio_output_cap),
    .X(_312_));
 sky130_fd_sc_hd__clkbuf_1 _641_ (.A(_312_),
    .X(_103_));
 sky130_fd_sc_hd__mux2_1 _642_ (.A0(\aio_output_reg[3] ),
    .A1(net85),
    .S(aio_output_cap),
    .X(_313_));
 sky130_fd_sc_hd__clkbuf_1 _643_ (.A(_313_),
    .X(_104_));
 sky130_fd_sc_hd__mux2_1 _644_ (.A0(\aio_output_reg[4] ),
    .A1(net89),
    .S(aio_output_cap),
    .X(_314_));
 sky130_fd_sc_hd__clkbuf_1 _645_ (.A(_314_),
    .X(_105_));
 sky130_fd_sc_hd__mux2_1 _646_ (.A0(\aio_output_reg[5] ),
    .A1(net88),
    .S(aio_output_cap),
    .X(_315_));
 sky130_fd_sc_hd__clkbuf_1 _647_ (.A(_315_),
    .X(_106_));
 sky130_fd_sc_hd__mux2_1 _648_ (.A0(\aio_output_reg[6] ),
    .A1(net91),
    .S(aio_output_cap),
    .X(_316_));
 sky130_fd_sc_hd__clkbuf_1 _649_ (.A(_316_),
    .X(_107_));
 sky130_fd_sc_hd__mux2_1 _650_ (.A0(\aio_output_reg[7] ),
    .A1(net84),
    .S(aio_output_cap),
    .X(_317_));
 sky130_fd_sc_hd__clkbuf_1 _651_ (.A(_317_),
    .X(_108_));
 sky130_fd_sc_hd__inv_2 _652_ (.A(_269_),
    .Y(_044_));
 sky130_fd_sc_hd__inv_2 _653_ (.A(_269_),
    .Y(_045_));
 sky130_fd_sc_hd__inv_2 _654_ (.A(_269_),
    .Y(_046_));
 sky130_fd_sc_hd__or4_1 _655_ (.A(\state[1] ),
    .B(\state[6] ),
    .C(\state[2] ),
    .D(\state[3] ),
    .X(_318_));
 sky130_fd_sc_hd__o2bb2a_2 _656_ (.A1_N(_175_),
    .A2_N(_187_),
    .B1(_318_),
    .B2(\state[8] ),
    .X(_319_));
 sky130_fd_sc_hd__and2_1 _657_ (.A(_172_),
    .B(_319_),
    .X(_320_));
 sky130_fd_sc_hd__clkbuf_1 _658_ (.A(_320_),
    .X(_109_));
 sky130_fd_sc_hd__or2_1 _659_ (.A(\ws_cnt[0] ),
    .B(\ws_cnt[1] ),
    .X(_321_));
 sky130_fd_sc_hd__nand2_1 _660_ (.A(\ws_cnt[0] ),
    .B(\ws_cnt[1] ),
    .Y(_322_));
 sky130_fd_sc_hd__and3_1 _661_ (.A(_319_),
    .B(_321_),
    .C(_322_),
    .X(_323_));
 sky130_fd_sc_hd__clkbuf_1 _662_ (.A(_323_),
    .X(_110_));
 sky130_fd_sc_hd__nand3_1 _663_ (.A(\ws_cnt[0] ),
    .B(\ws_cnt[1] ),
    .C(\ws_cnt[2] ),
    .Y(_324_));
 sky130_fd_sc_hd__a21o_1 _664_ (.A1(\ws_cnt[0] ),
    .A2(\ws_cnt[1] ),
    .B1(\ws_cnt[2] ),
    .X(_325_));
 sky130_fd_sc_hd__and3_1 _665_ (.A(_319_),
    .B(_324_),
    .C(_325_),
    .X(_326_));
 sky130_fd_sc_hd__clkbuf_1 _666_ (.A(_326_),
    .X(_111_));
 sky130_fd_sc_hd__and4_1 _667_ (.A(\ws_cnt[0] ),
    .B(\ws_cnt[1] ),
    .C(\ws_cnt[2] ),
    .D(\ws_cnt[3] ),
    .X(_327_));
 sky130_fd_sc_hd__a31o_1 _668_ (.A1(\ws_cnt[0] ),
    .A2(\ws_cnt[1] ),
    .A3(\ws_cnt[2] ),
    .B1(\ws_cnt[3] ),
    .X(_328_));
 sky130_fd_sc_hd__and3b_1 _669_ (.A_N(_327_),
    .B(_328_),
    .C(_319_),
    .X(_329_));
 sky130_fd_sc_hd__clkbuf_1 _670_ (.A(_329_),
    .X(_112_));
 sky130_fd_sc_hd__and2_1 _671_ (.A(\ws_cnt[4] ),
    .B(_327_),
    .X(_330_));
 sky130_fd_sc_hd__or2_1 _672_ (.A(\ws_cnt[4] ),
    .B(_327_),
    .X(_331_));
 sky130_fd_sc_hd__and3b_1 _673_ (.A_N(_330_),
    .B(_331_),
    .C(_319_),
    .X(_332_));
 sky130_fd_sc_hd__clkbuf_1 _674_ (.A(_332_),
    .X(_113_));
 sky130_fd_sc_hd__and3_1 _675_ (.A(\ws_cnt[4] ),
    .B(\ws_cnt[5] ),
    .C(_327_),
    .X(_333_));
 sky130_fd_sc_hd__or2_1 _676_ (.A(\ws_cnt[5] ),
    .B(_330_),
    .X(_334_));
 sky130_fd_sc_hd__and3b_1 _677_ (.A_N(_333_),
    .B(_334_),
    .C(_319_),
    .X(_335_));
 sky130_fd_sc_hd__clkbuf_1 _678_ (.A(_335_),
    .X(_114_));
 sky130_fd_sc_hd__or2_1 _679_ (.A(\ws_cnt[6] ),
    .B(_333_),
    .X(_336_));
 sky130_fd_sc_hd__nand2_1 _680_ (.A(\ws_cnt[6] ),
    .B(_333_),
    .Y(_337_));
 sky130_fd_sc_hd__and3_1 _681_ (.A(_319_),
    .B(_336_),
    .C(_337_),
    .X(_338_));
 sky130_fd_sc_hd__clkbuf_1 _682_ (.A(_338_),
    .X(_115_));
 sky130_fd_sc_hd__nand2_1 _683_ (.A(_173_),
    .B(_337_),
    .Y(_339_));
 sky130_fd_sc_hd__o211a_1 _684_ (.A1(_173_),
    .A2(_337_),
    .B1(_339_),
    .C1(_319_),
    .X(_116_));
 sky130_fd_sc_hd__inv_2 _685_ (.A(_269_),
    .Y(_047_));
 sky130_fd_sc_hd__inv_2 _686_ (.A(_269_),
    .Y(_048_));
 sky130_fd_sc_hd__inv_2 _687_ (.A(_269_),
    .Y(_049_));
 sky130_fd_sc_hd__inv_2 _688_ (.A(_269_),
    .Y(_050_));
 sky130_fd_sc_hd__inv_2 _689_ (.A(_250_),
    .Y(_051_));
 sky130_fd_sc_hd__inv_2 _690_ (.A(_250_),
    .Y(_052_));
 sky130_fd_sc_hd__inv_2 _691_ (.A(_250_),
    .Y(_053_));
 sky130_fd_sc_hd__inv_2 _692_ (.A(_250_),
    .Y(_054_));
 sky130_fd_sc_hd__inv_2 _693_ (.A(_250_),
    .Y(_055_));
 sky130_fd_sc_hd__dfrtp_1 _694_ (.CLK(clknet_3_3__leaf_clk),
    .D(_056_),
    .RESET_B(_015_),
    .Q(\state[8] ));
 sky130_fd_sc_hd__dfxtp_1 _695_ (.CLK(clknet_3_1__leaf_clk),
    .D(_057_),
    .Q(\aio_input_shift[1] ));
 sky130_fd_sc_hd__dfxtp_1 _696_ (.CLK(clknet_3_3__leaf_clk),
    .D(_058_),
    .Q(\aio_input_shift[2] ));
 sky130_fd_sc_hd__dfxtp_1 _697_ (.CLK(clknet_3_4__leaf_clk),
    .D(_059_),
    .Q(\aio_input_shift[3] ));
 sky130_fd_sc_hd__dfxtp_1 _698_ (.CLK(clknet_3_4__leaf_clk),
    .D(_060_),
    .Q(\aio_input_shift[4] ));
 sky130_fd_sc_hd__dfxtp_1 _699_ (.CLK(clknet_3_5__leaf_clk),
    .D(_061_),
    .Q(\aio_input_shift[5] ));
 sky130_fd_sc_hd__dfxtp_1 _700_ (.CLK(clknet_3_5__leaf_clk),
    .D(_062_),
    .Q(\aio_input_shift[6] ));
 sky130_fd_sc_hd__dfxtp_1 _701_ (.CLK(clknet_3_5__leaf_clk),
    .D(_063_),
    .Q(\aio_input_shift[7] ));
 sky130_fd_sc_hd__dfstp_1 _702_ (.CLK(clknet_3_6__leaf_clk),
    .D(_007_),
    .SET_B(_016_),
    .Q(\state[0] ));
 sky130_fd_sc_hd__dfrtp_1 _703_ (.CLK(clknet_3_6__leaf_clk),
    .D(_008_),
    .RESET_B(_017_),
    .Q(\state[1] ));
 sky130_fd_sc_hd__dfrtp_1 _704_ (.CLK(clknet_3_6__leaf_clk),
    .D(_009_),
    .RESET_B(_018_),
    .Q(\state[2] ));
 sky130_fd_sc_hd__dfrtp_1 _705_ (.CLK(clknet_3_3__leaf_clk),
    .D(_010_),
    .RESET_B(_019_),
    .Q(\state[3] ));
 sky130_fd_sc_hd__dfrtp_1 _706_ (.CLK(clknet_3_4__leaf_clk),
    .D(_011_),
    .RESET_B(_020_),
    .Q(\state[4] ));
 sky130_fd_sc_hd__dfrtp_1 _707_ (.CLK(clknet_3_6__leaf_clk),
    .D(_012_),
    .RESET_B(_021_),
    .Q(\state[5] ));
 sky130_fd_sc_hd__dfrtp_1 _708_ (.CLK(clknet_3_6__leaf_clk),
    .D(_013_),
    .RESET_B(_022_),
    .Q(\state[6] ));
 sky130_fd_sc_hd__dfrtp_4 _709_ (.CLK(clknet_3_5__leaf_clk),
    .D(net36),
    .RESET_B(_023_),
    .Q(\clk_divider_I.ce ));
 sky130_fd_sc_hd__dfrtp_1 _710_ (.CLK(clknet_3_3__leaf_clk),
    .D(_004_),
    .RESET_B(_024_),
    .Q(\state[9] ));
 sky130_fd_sc_hd__dfrtp_4 _711_ (.CLK(clknet_3_3__leaf_clk),
    .D(_005_),
    .RESET_B(_025_),
    .Q(aio_output_cap));
 sky130_fd_sc_hd__dfrtp_2 _712_ (.CLK(clknet_3_4__leaf_clk),
    .D(\state[4] ),
    .RESET_B(_026_),
    .Q(aio_input_sh));
 sky130_fd_sc_hd__dfrtp_2 _713_ (.CLK(clknet_3_6__leaf_clk),
    .D(\state[5] ),
    .RESET_B(_027_),
    .Q(\state[12] ));
 sky130_fd_sc_hd__dfrtp_1 _714_ (.CLK(clknet_3_6__leaf_clk),
    .D(_006_),
    .RESET_B(_028_),
    .Q(\state[13] ));
 sky130_fd_sc_hd__dfxtp_1 _715_ (.CLK(clknet_3_4__leaf_clk),
    .D(_064_),
    .Q(\aio_input_shift[0] ));
 sky130_fd_sc_hd__dfrtp_1 _716_ (.CLK(clknet_3_2__leaf_clk),
    .D(_065_),
    .RESET_B(_029_),
    .Q(\ws_cfg[0] ));
 sky130_fd_sc_hd__dfstp_1 _717_ (.CLK(clknet_3_2__leaf_clk),
    .D(_066_),
    .SET_B(_030_),
    .Q(\ws_cfg[1] ));
 sky130_fd_sc_hd__dfrtp_1 _718_ (.CLK(clknet_3_3__leaf_clk),
    .D(_067_),
    .RESET_B(_031_),
    .Q(\ws_cfg[2] ));
 sky130_fd_sc_hd__dfstp_1 _719_ (.CLK(clknet_3_3__leaf_clk),
    .D(_068_),
    .SET_B(_032_),
    .Q(\ws_cfg[3] ));
 sky130_fd_sc_hd__dfrtp_1 _720_ (.CLK(clknet_3_2__leaf_clk),
    .D(_069_),
    .RESET_B(_033_),
    .Q(\ws_cfg[4] ));
 sky130_fd_sc_hd__dfrtp_1 _721_ (.CLK(clknet_3_2__leaf_clk),
    .D(_070_),
    .RESET_B(_034_),
    .Q(\ws_cfg[5] ));
 sky130_fd_sc_hd__dfrtp_1 _722_ (.CLK(clknet_3_1__leaf_clk),
    .D(_071_),
    .RESET_B(_035_),
    .Q(\ws_cfg[6] ));
 sky130_fd_sc_hd__dfrtp_1 _723_ (.CLK(clknet_3_3__leaf_clk),
    .D(_072_),
    .RESET_B(_036_),
    .Q(\ws_cfg[7] ));
 sky130_fd_sc_hd__dfstp_1 _724_ (.CLK(net81),
    .D(net42),
    .SET_B(_037_),
    .Q(\rst_shift[0] ));
 sky130_fd_sc_hd__conb_1 _724__42 (.LO(net42));
 sky130_fd_sc_hd__dfstp_1 _725_ (.CLK(net82),
    .D(\rst_shift[0] ),
    .SET_B(_039_),
    .Q(\rst_shift[1] ));
 sky130_fd_sc_hd__dfstp_1 _726_ (.CLK(net83),
    .D(\rst_shift[1] ),
    .SET_B(_041_),
    .Q(\clk_divider_I.reset ));
 sky130_fd_sc_hd__dfxtp_1 _727_ (.CLK(clknet_3_1__leaf_clk),
    .D(net12),
    .Q(\aio_input_sync[0] ));
 sky130_fd_sc_hd__dfxtp_1 _728_ (.CLK(clknet_3_1__leaf_clk),
    .D(net13),
    .Q(\aio_input_sync[1] ));
 sky130_fd_sc_hd__dfxtp_1 _729_ (.CLK(clknet_3_3__leaf_clk),
    .D(net14),
    .Q(\aio_input_sync[2] ));
 sky130_fd_sc_hd__dfxtp_1 _730_ (.CLK(clknet_3_3__leaf_clk),
    .D(net15),
    .Q(\aio_input_sync[3] ));
 sky130_fd_sc_hd__dfxtp_1 _731_ (.CLK(clknet_3_4__leaf_clk),
    .D(net16),
    .Q(\aio_input_sync[4] ));
 sky130_fd_sc_hd__dfxtp_1 _732_ (.CLK(clknet_3_1__leaf_clk),
    .D(net17),
    .Q(\aio_input_sync[5] ));
 sky130_fd_sc_hd__dfxtp_1 _733_ (.CLK(clknet_3_0__leaf_clk),
    .D(net18),
    .Q(\aio_input_sync[6] ));
 sky130_fd_sc_hd__dfxtp_1 _734_ (.CLK(clknet_3_5__leaf_clk),
    .D(net19),
    .Q(\aio_input_sync[7] ));
 sky130_fd_sc_hd__dfxtp_1 _735_ (.CLK(clknet_3_1__leaf_clk),
    .D(_073_),
    .Q(\clk_divider_I.compare[0] ));
 sky130_fd_sc_hd__dfxtp_1 _736_ (.CLK(clknet_3_1__leaf_clk),
    .D(_074_),
    .Q(\clk_divider_I.compare[1] ));
 sky130_fd_sc_hd__dfxtp_1 _737_ (.CLK(clknet_3_1__leaf_clk),
    .D(_075_),
    .Q(\clk_divider_I.compare[2] ));
 sky130_fd_sc_hd__dfxtp_1 _738_ (.CLK(clknet_3_1__leaf_clk),
    .D(_076_),
    .Q(\clk_divider_I.compare[3] ));
 sky130_fd_sc_hd__dfxtp_1 _739_ (.CLK(clknet_3_1__leaf_clk),
    .D(_077_),
    .Q(\clk_divider_I.compare[4] ));
 sky130_fd_sc_hd__dfxtp_1 _740_ (.CLK(clknet_3_0__leaf_clk),
    .D(_078_),
    .Q(\clk_divider_I.compare[5] ));
 sky130_fd_sc_hd__dfxtp_1 _741_ (.CLK(clknet_3_0__leaf_clk),
    .D(_079_),
    .Q(\clk_divider_I.compare[6] ));
 sky130_fd_sc_hd__dfxtp_1 _742_ (.CLK(clknet_3_1__leaf_clk),
    .D(_080_),
    .Q(\clk_divider_I.compare[7] ));
 sky130_fd_sc_hd__dfrtp_1 _743_ (.CLK(clknet_3_4__leaf_clk),
    .D(net11),
    .RESET_B(_043_),
    .Q(active));
 sky130_fd_sc_hd__dfxtp_1 _744_ (.CLK(clknet_3_7__leaf_clk),
    .D(_081_),
    .Q(\bit_cnt[0] ));
 sky130_fd_sc_hd__dfxtp_1 _745_ (.CLK(clknet_3_7__leaf_clk),
    .D(_082_),
    .Q(\bit_cnt[1] ));
 sky130_fd_sc_hd__dfxtp_1 _746_ (.CLK(clknet_3_7__leaf_clk),
    .D(_083_),
    .Q(\bit_cnt[2] ));
 sky130_fd_sc_hd__dfxtp_1 _747_ (.CLK(clknet_3_7__leaf_clk),
    .D(_084_),
    .Q(\proj_cnt[0] ));
 sky130_fd_sc_hd__dfxtp_1 _748_ (.CLK(clknet_3_7__leaf_clk),
    .D(_085_),
    .Q(\proj_cnt[1] ));
 sky130_fd_sc_hd__dfxtp_1 _749_ (.CLK(clknet_3_7__leaf_clk),
    .D(_086_),
    .Q(\proj_cnt[2] ));
 sky130_fd_sc_hd__dfxtp_1 _750_ (.CLK(clknet_3_7__leaf_clk),
    .D(_087_),
    .Q(\proj_cnt[3] ));
 sky130_fd_sc_hd__dfxtp_1 _751_ (.CLK(clknet_3_6__leaf_clk),
    .D(_088_),
    .Q(\proj_cnt[4] ));
 sky130_fd_sc_hd__dfxtp_1 _752_ (.CLK(clknet_3_6__leaf_clk),
    .D(_089_),
    .Q(\proj_cnt[5] ));
 sky130_fd_sc_hd__dfxtp_1 _753_ (.CLK(clknet_3_7__leaf_clk),
    .D(_090_),
    .Q(\proj_cnt[6] ));
 sky130_fd_sc_hd__dfxtp_1 _754_ (.CLK(clknet_3_7__leaf_clk),
    .D(_091_),
    .Q(\proj_cnt[7] ));
 sky130_fd_sc_hd__dfxtp_1 _755_ (.CLK(clknet_3_7__leaf_clk),
    .D(_092_),
    .Q(\proj_cnt[8] ));
 sky130_fd_sc_hd__dfxtp_1 _756_ (.CLK(clknet_3_6__leaf_clk),
    .D(_000_),
    .Q(int_scan_clk_out));
 sky130_fd_sc_hd__dfxtp_1 _757_ (.CLK(clknet_3_3__leaf_clk),
    .D(\aio_input_shift[7] ),
    .Q(int_scan_data_out));
 sky130_fd_sc_hd__dfxtp_1 _758_ (.CLK(clknet_3_6__leaf_clk),
    .D(_001_),
    .Q(int_scan_select));
 sky130_fd_sc_hd__dfxtp_1 _759_ (.CLK(clknet_3_6__leaf_clk),
    .D(\state[9] ),
    .Q(int_scan_latch_en));
 sky130_fd_sc_hd__dfxtp_1 _760_ (.CLK(clknet_3_1__leaf_clk),
    .D(_093_),
    .Q(\aio_input_reg[0] ));
 sky130_fd_sc_hd__dfxtp_1 _761_ (.CLK(clknet_3_1__leaf_clk),
    .D(_094_),
    .Q(\aio_input_reg[1] ));
 sky130_fd_sc_hd__dfxtp_1 _762_ (.CLK(clknet_3_3__leaf_clk),
    .D(_095_),
    .Q(\aio_input_reg[2] ));
 sky130_fd_sc_hd__dfxtp_1 _763_ (.CLK(clknet_3_3__leaf_clk),
    .D(_096_),
    .Q(\aio_input_reg[3] ));
 sky130_fd_sc_hd__dfxtp_1 _764_ (.CLK(clknet_3_4__leaf_clk),
    .D(_097_),
    .Q(\aio_input_reg[4] ));
 sky130_fd_sc_hd__dfxtp_1 _765_ (.CLK(clknet_3_4__leaf_clk),
    .D(_098_),
    .Q(\aio_input_reg[5] ));
 sky130_fd_sc_hd__dfxtp_1 _766_ (.CLK(clknet_3_5__leaf_clk),
    .D(_099_),
    .Q(\aio_input_reg[6] ));
 sky130_fd_sc_hd__dfxtp_1 _767_ (.CLK(clknet_3_5__leaf_clk),
    .D(_100_),
    .Q(\aio_input_reg[7] ));
 sky130_fd_sc_hd__dfxtp_1 _768_ (.CLK(clknet_1_0__leaf_scan_clk_in),
    .D(net25),
    .Q(\aio_output_shift[0] ));
 sky130_fd_sc_hd__dfxtp_1 _769_ (.CLK(clknet_1_0__leaf_scan_clk_in),
    .D(\aio_output_shift[0] ),
    .Q(\aio_output_shift[1] ));
 sky130_fd_sc_hd__dfxtp_1 _770_ (.CLK(clknet_1_1__leaf_scan_clk_in),
    .D(\aio_output_shift[1] ),
    .Q(\aio_output_shift[2] ));
 sky130_fd_sc_hd__dfxtp_1 _771_ (.CLK(clknet_1_1__leaf_scan_clk_in),
    .D(\aio_output_shift[2] ),
    .Q(\aio_output_shift[3] ));
 sky130_fd_sc_hd__dfxtp_1 _772_ (.CLK(clknet_1_1__leaf_scan_clk_in),
    .D(\aio_output_shift[3] ),
    .Q(\aio_output_shift[4] ));
 sky130_fd_sc_hd__dfxtp_1 _773_ (.CLK(clknet_1_0__leaf_scan_clk_in),
    .D(\aio_output_shift[4] ),
    .Q(\aio_output_shift[5] ));
 sky130_fd_sc_hd__dfxtp_1 _774_ (.CLK(clknet_1_0__leaf_scan_clk_in),
    .D(\aio_output_shift[5] ),
    .Q(\aio_output_shift[6] ));
 sky130_fd_sc_hd__dfxtp_1 _775_ (.CLK(clknet_1_0__leaf_scan_clk_in),
    .D(\aio_output_shift[6] ),
    .Q(\aio_output_shift[7] ));
 sky130_fd_sc_hd__dfxtp_1 _776_ (.CLK(clknet_3_2__leaf_clk),
    .D(_101_),
    .Q(\aio_output_reg[0] ));
 sky130_fd_sc_hd__dfxtp_1 _777_ (.CLK(clknet_3_2__leaf_clk),
    .D(_102_),
    .Q(\aio_output_reg[1] ));
 sky130_fd_sc_hd__dfxtp_1 _778_ (.CLK(clknet_3_0__leaf_clk),
    .D(_103_),
    .Q(\aio_output_reg[2] ));
 sky130_fd_sc_hd__dfxtp_1 _779_ (.CLK(clknet_3_2__leaf_clk),
    .D(_104_),
    .Q(\aio_output_reg[3] ));
 sky130_fd_sc_hd__dfxtp_1 _780_ (.CLK(clknet_3_0__leaf_clk),
    .D(_105_),
    .Q(\aio_output_reg[4] ));
 sky130_fd_sc_hd__dfxtp_1 _781_ (.CLK(clknet_3_0__leaf_clk),
    .D(_106_),
    .Q(\aio_output_reg[5] ));
 sky130_fd_sc_hd__dfxtp_1 _782_ (.CLK(clknet_3_0__leaf_clk),
    .D(_107_),
    .Q(\aio_output_reg[6] ));
 sky130_fd_sc_hd__dfxtp_1 _783_ (.CLK(clknet_3_0__leaf_clk),
    .D(_108_),
    .Q(\aio_output_reg[7] ));
 sky130_fd_sc_hd__dfrtp_1 _784_ (.CLK(clknet_3_0__leaf_clk),
    .D(_003_),
    .RESET_B(_044_),
    .Q(\ws_set_sync[0] ));
 sky130_fd_sc_hd__dfrtp_1 _785_ (.CLK(clknet_3_0__leaf_clk),
    .D(\ws_set_sync[0] ),
    .RESET_B(_045_),
    .Q(\ws_set_sync[1] ));
 sky130_fd_sc_hd__dfrtp_1 _786_ (.CLK(clknet_3_0__leaf_clk),
    .D(\ws_set_sync[1] ),
    .RESET_B(_046_),
    .Q(\ws_set_sync[2] ));
 sky130_fd_sc_hd__dfxtp_2 _787_ (.CLK(clknet_3_0__leaf_clk),
    .D(_002_),
    .Q(ws_set_now));
 sky130_fd_sc_hd__dfxtp_1 _788_ (.CLK(clknet_3_2__leaf_clk),
    .D(_109_),
    .Q(\ws_cnt[0] ));
 sky130_fd_sc_hd__dfxtp_1 _789_ (.CLK(clknet_3_2__leaf_clk),
    .D(_110_),
    .Q(\ws_cnt[1] ));
 sky130_fd_sc_hd__dfxtp_1 _790_ (.CLK(clknet_3_3__leaf_clk),
    .D(_111_),
    .Q(\ws_cnt[2] ));
 sky130_fd_sc_hd__dfxtp_1 _791_ (.CLK(clknet_3_3__leaf_clk),
    .D(_112_),
    .Q(\ws_cnt[3] ));
 sky130_fd_sc_hd__dfxtp_1 _792_ (.CLK(clknet_3_2__leaf_clk),
    .D(_113_),
    .Q(\ws_cnt[4] ));
 sky130_fd_sc_hd__dfxtp_1 _793_ (.CLK(clknet_3_2__leaf_clk),
    .D(_114_),
    .Q(\ws_cnt[5] ));
 sky130_fd_sc_hd__dfxtp_1 _794_ (.CLK(clknet_3_2__leaf_clk),
    .D(_115_),
    .Q(\ws_cnt[6] ));
 sky130_fd_sc_hd__dfxtp_1 _795_ (.CLK(clknet_3_2__leaf_clk),
    .D(_116_),
    .Q(\ws_cnt[7] ));
 sky130_fd_sc_hd__dfxtp_2 _796_ (.CLK(clknet_3_1__leaf_clk),
    .D(_014_),
    .Q(\clk_divider_I.set_now ));
 sky130_fd_sc_hd__dfxtp_1 _797_ (.CLK(clknet_3_2__leaf_clk),
    .D(net26),
    .Q(\clk_divider_I.set_sync[0] ));
 sky130_fd_sc_hd__dfxtp_1 _798_ (.CLK(clknet_3_2__leaf_clk),
    .D(\clk_divider_I.set_sync[0] ),
    .Q(\clk_divider_I.set_sync[1] ));
 sky130_fd_sc_hd__dfxtp_1 _799_ (.CLK(clknet_3_0__leaf_clk),
    .D(\clk_divider_I.set_sync[1] ),
    .Q(\clk_divider_I.active ));
 sky130_fd_sc_hd__dfrtp_4 _800_ (.CLK(clknet_3_5__leaf_clk),
    .D(_117_),
    .RESET_B(_047_),
    .Q(\clk_divider_I.counter[0] ));
 sky130_fd_sc_hd__dfrtp_2 _801_ (.CLK(clknet_3_5__leaf_clk),
    .D(_118_),
    .RESET_B(_048_),
    .Q(\clk_divider_I.counter[1] ));
 sky130_fd_sc_hd__dfrtp_1 _802_ (.CLK(clknet_3_5__leaf_clk),
    .D(_119_),
    .RESET_B(_049_),
    .Q(\clk_divider_I.counter[2] ));
 sky130_fd_sc_hd__dfrtp_1 _803_ (.CLK(clknet_3_4__leaf_clk),
    .D(_120_),
    .RESET_B(_050_),
    .Q(\clk_divider_I.counter[3] ));
 sky130_fd_sc_hd__dfrtp_1 _804_ (.CLK(clknet_3_4__leaf_clk),
    .D(_121_),
    .RESET_B(_051_),
    .Q(\clk_divider_I.counter[4] ));
 sky130_fd_sc_hd__dfrtp_1 _805_ (.CLK(clknet_3_4__leaf_clk),
    .D(_122_),
    .RESET_B(_052_),
    .Q(\clk_divider_I.counter[5] ));
 sky130_fd_sc_hd__dfrtp_1 _806_ (.CLK(clknet_3_4__leaf_clk),
    .D(_123_),
    .RESET_B(_053_),
    .Q(\clk_divider_I.counter[6] ));
 sky130_fd_sc_hd__dfrtp_1 _807_ (.CLK(clknet_3_4__leaf_clk),
    .D(_124_),
    .RESET_B(_054_),
    .Q(\clk_divider_I.counter[7] ));
 sky130_fd_sc_hd__dfrtp_2 _808_ (.CLK(clknet_3_4__leaf_clk),
    .D(_125_),
    .RESET_B(_055_),
    .Q(net41));
 sky130_fd_sc_hd__clkbuf_1 _848_ (.A(net25),
    .X(net27));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_scan_clk_in (.A(scan_clk_in),
    .X(clknet_0_scan_clk_in));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_scan_clk_in (.A(clknet_0_scan_clk_in),
    .X(clknet_1_0__leaf_scan_clk_in));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_scan_clk_in (.A(clknet_0_scan_clk_in),
    .X(clknet_1_1__leaf_scan_clk_in));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_0__f_clk (.A(clknet_0_clk),
    .X(clknet_3_0__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_1__f_clk (.A(clknet_0_clk),
    .X(clknet_3_1__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_2__f_clk (.A(clknet_0_clk),
    .X(clknet_3_2__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_3__f_clk (.A(clknet_0_clk),
    .X(clknet_3_3__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_4__f_clk (.A(clknet_0_clk),
    .X(clknet_3_4__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_5__f_clk (.A(clknet_0_clk),
    .X(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_6__f_clk (.A(clknet_0_clk),
    .X(clknet_3_6__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_7__f_clk (.A(clknet_0_clk),
    .X(clknet_3_7__leaf_clk));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1 (.A(\aio_output_shift[7] ),
    .X(net84));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2 (.A(\aio_output_shift[3] ),
    .X(net85));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3 (.A(\aio_output_shift[0] ),
    .X(net86));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4 (.A(\aio_output_shift[2] ),
    .X(net87));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5 (.A(\aio_output_shift[5] ),
    .X(net88));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6 (.A(\aio_output_shift[4] ),
    .X(net89));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7 (.A(\aio_output_shift[1] ),
    .X(net90));
 sky130_fd_sc_hd__dlygate4sd3_1 hold8 (.A(\aio_output_shift[6] ),
    .X(net91));
 sky130_fd_sc_hd__clkbuf_2 input1 (.A(active_select[0]),
    .X(net1));
 sky130_fd_sc_hd__buf_2 input10 (.A(driver_sel[0]),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_2 input11 (.A(driver_sel[1]),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_2 input12 (.A(inputs[0]),
    .X(net12));
 sky130_fd_sc_hd__dlymetal6s2s_1 input13 (.A(inputs[1]),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_2 input14 (.A(inputs[2]),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_2 input15 (.A(inputs[3]),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_2 input16 (.A(inputs[4]),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_1 input17 (.A(inputs[5]),
    .X(net17));
 sky130_fd_sc_hd__clkbuf_1 input18 (.A(inputs[6]),
    .X(net18));
 sky130_fd_sc_hd__clkbuf_2 input19 (.A(inputs[7]),
    .X(net19));
 sky130_fd_sc_hd__clkbuf_1 input2 (.A(active_select[1]),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_1 input20 (.A(la_scan_clk_in),
    .X(net20));
 sky130_fd_sc_hd__clkbuf_1 input21 (.A(la_scan_data_in),
    .X(net21));
 sky130_fd_sc_hd__clkbuf_1 input22 (.A(la_scan_latch_en),
    .X(net22));
 sky130_fd_sc_hd__clkbuf_1 input23 (.A(la_scan_select),
    .X(net23));
 sky130_fd_sc_hd__dlymetal6s2s_1 input24 (.A(reset),
    .X(net24));
 sky130_fd_sc_hd__clkbuf_2 input25 (.A(scan_data_in),
    .X(net25));
 sky130_fd_sc_hd__clkbuf_1 input26 (.A(set_clk_div),
    .X(net26));
 sky130_fd_sc_hd__clkbuf_1 input3 (.A(active_select[2]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_1 input4 (.A(active_select[3]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_1 input5 (.A(active_select[4]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_1 input6 (.A(active_select[5]),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_1 input7 (.A(active_select[6]),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_2 input8 (.A(active_select[7]),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_2 input9 (.A(active_select[8]),
    .X(net9));
 sky130_fd_sc_hd__buf_2 output27 (.A(net27),
    .X(la_scan_data_out));
 sky130_fd_sc_hd__clkbuf_1 output28 (.A(net28),
    .X(outputs[0]));
 sky130_fd_sc_hd__buf_2 output29 (.A(net29),
    .X(outputs[1]));
 sky130_fd_sc_hd__buf_2 output30 (.A(net30),
    .X(outputs[2]));
 sky130_fd_sc_hd__buf_2 output31 (.A(net31),
    .X(outputs[3]));
 sky130_fd_sc_hd__buf_2 output32 (.A(net32),
    .X(outputs[4]));
 sky130_fd_sc_hd__buf_2 output33 (.A(net33),
    .X(outputs[5]));
 sky130_fd_sc_hd__buf_2 output34 (.A(net34),
    .X(outputs[6]));
 sky130_fd_sc_hd__buf_2 output35 (.A(net35),
    .X(outputs[7]));
 sky130_fd_sc_hd__buf_2 output36 (.A(net36),
    .X(ready));
 sky130_fd_sc_hd__buf_2 output37 (.A(net37),
    .X(scan_clk_out));
 sky130_fd_sc_hd__buf_2 output38 (.A(net38),
    .X(scan_data_out));
 sky130_fd_sc_hd__buf_2 output39 (.A(net39),
    .X(scan_latch_en));
 sky130_fd_sc_hd__buf_2 output40 (.A(net40),
    .X(scan_select));
 sky130_fd_sc_hd__buf_2 output41 (.A(net41),
    .X(slow_clk));
 sky130_fd_sc_hd__conb_1 scan_controller_43 (.LO(net43));
 sky130_fd_sc_hd__conb_1 scan_controller_44 (.LO(net44));
 sky130_fd_sc_hd__conb_1 scan_controller_45 (.LO(net45));
 sky130_fd_sc_hd__conb_1 scan_controller_46 (.LO(net46));
 sky130_fd_sc_hd__conb_1 scan_controller_47 (.LO(net47));
 sky130_fd_sc_hd__conb_1 scan_controller_48 (.LO(net48));
 sky130_fd_sc_hd__conb_1 scan_controller_49 (.LO(net49));
 sky130_fd_sc_hd__conb_1 scan_controller_50 (.LO(net50));
 sky130_fd_sc_hd__conb_1 scan_controller_51 (.LO(net51));
 sky130_fd_sc_hd__conb_1 scan_controller_52 (.LO(net52));
 sky130_fd_sc_hd__conb_1 scan_controller_53 (.LO(net53));
 sky130_fd_sc_hd__conb_1 scan_controller_54 (.LO(net54));
 sky130_fd_sc_hd__conb_1 scan_controller_55 (.LO(net55));
 sky130_fd_sc_hd__conb_1 scan_controller_56 (.LO(net56));
 sky130_fd_sc_hd__conb_1 scan_controller_57 (.LO(net57));
 sky130_fd_sc_hd__conb_1 scan_controller_58 (.LO(net58));
 sky130_fd_sc_hd__conb_1 scan_controller_59 (.LO(net59));
 sky130_fd_sc_hd__conb_1 scan_controller_60 (.LO(net60));
 sky130_fd_sc_hd__conb_1 scan_controller_61 (.LO(net61));
 sky130_fd_sc_hd__conb_1 scan_controller_62 (.LO(net62));
 sky130_fd_sc_hd__conb_1 scan_controller_63 (.LO(net63));
 sky130_fd_sc_hd__conb_1 scan_controller_64 (.LO(net64));
 sky130_fd_sc_hd__conb_1 scan_controller_65 (.LO(net65));
 sky130_fd_sc_hd__conb_1 scan_controller_66 (.LO(net66));
 sky130_fd_sc_hd__conb_1 scan_controller_67 (.LO(net67));
 sky130_fd_sc_hd__conb_1 scan_controller_68 (.LO(net68));
 sky130_fd_sc_hd__conb_1 scan_controller_69 (.LO(net69));
 sky130_fd_sc_hd__conb_1 scan_controller_70 (.LO(net70));
 sky130_fd_sc_hd__conb_1 scan_controller_71 (.LO(net71));
 sky130_fd_sc_hd__conb_1 scan_controller_72 (.LO(net72));
 sky130_fd_sc_hd__conb_1 scan_controller_73 (.LO(net73));
 sky130_fd_sc_hd__conb_1 scan_controller_74 (.LO(net74));
 sky130_fd_sc_hd__conb_1 scan_controller_75 (.LO(net75));
 sky130_fd_sc_hd__conb_1 scan_controller_76 (.LO(net76));
 sky130_fd_sc_hd__conb_1 scan_controller_77 (.LO(net77));
 sky130_fd_sc_hd__conb_1 scan_controller_78 (.LO(net78));
 sky130_fd_sc_hd__conb_1 scan_controller_79 (.LO(net79));
 sky130_fd_sc_hd__conb_1 scan_controller_80 (.LO(net80));
 assign oeb[0] = net43;
 assign oeb[10] = net53;
 assign oeb[11] = net54;
 assign oeb[12] = net55;
 assign oeb[13] = net56;
 assign oeb[14] = net57;
 assign oeb[15] = net58;
 assign oeb[16] = net59;
 assign oeb[17] = net60;
 assign oeb[18] = net61;
 assign oeb[19] = net62;
 assign oeb[1] = net44;
 assign oeb[20] = net63;
 assign oeb[21] = net64;
 assign oeb[22] = net65;
 assign oeb[23] = net66;
 assign oeb[24] = net67;
 assign oeb[25] = net68;
 assign oeb[26] = net69;
 assign oeb[27] = net70;
 assign oeb[28] = net71;
 assign oeb[29] = net72;
 assign oeb[2] = net45;
 assign oeb[30] = net73;
 assign oeb[31] = net74;
 assign oeb[32] = net75;
 assign oeb[33] = net76;
 assign oeb[34] = net77;
 assign oeb[35] = net78;
 assign oeb[36] = net79;
 assign oeb[37] = net80;
 assign oeb[3] = net46;
 assign oeb[4] = net47;
 assign oeb[5] = net48;
 assign oeb[6] = net49;
 assign oeb[7] = net50;
 assign oeb[8] = net51;
 assign oeb[9] = net52;
endmodule

