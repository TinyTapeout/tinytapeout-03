magic
tech sky130A
magscale 1 2
timestamp 1682077834
<< viali >>
rect 3886 11849 3920 11883
rect 3617 11713 3651 11747
rect 3890 11645 3924 11679
rect 4353 11645 4387 11679
rect 2513 11509 2547 11543
rect 3433 11237 3467 11271
rect 2421 11101 2455 11135
rect 2697 11101 2731 11135
rect 3886 10761 3920 10795
rect 3617 10625 3651 10659
rect 3890 10557 3924 10591
rect 4353 10557 4387 10591
rect 2513 10421 2547 10455
rect 2056 10081 2090 10115
rect 2329 10081 2363 10115
rect 1593 10013 1627 10047
rect 2059 9877 2093 9911
rect 3433 9877 3467 9911
rect 3886 9673 3920 9707
rect 3617 9469 3651 9503
rect 3847 9469 3881 9503
rect 4353 9469 4387 9503
rect 2513 9333 2547 9367
rect 2056 8993 2090 9027
rect 2329 8993 2363 9027
rect 1593 8925 1627 8959
rect 2059 8789 2093 8823
rect 3433 8789 3467 8823
rect 3886 8585 3920 8619
rect 3617 8449 3651 8483
rect 3874 8383 3908 8417
rect 4353 8381 4387 8415
rect 2513 8245 2547 8279
rect 2056 7887 2090 7921
rect 2329 7905 2363 7939
rect 1593 7837 1627 7871
rect 2059 7701 2093 7735
rect 3433 7701 3467 7735
rect 2513 7497 2547 7531
rect 3886 7497 3920 7531
rect 3617 7361 3651 7395
rect 3847 7293 3881 7327
rect 4353 7293 4387 7327
rect 3433 6953 3467 6987
rect 2421 6817 2455 6851
rect 2697 6749 2731 6783
rect 3985 6613 4019 6647
rect 2605 6341 2639 6375
rect 2329 6205 2363 6239
rect 4353 6205 4387 6239
rect 3433 5865 3467 5899
rect 2421 5729 2455 5763
rect 2697 5661 2731 5695
rect 4353 5321 4387 5355
rect 2145 5185 2179 5219
rect 3617 5185 3651 5219
rect 1869 5117 1903 5151
rect 3341 5117 3375 5151
rect 2881 4981 2915 5015
rect 4261 4777 4295 4811
rect 2421 4573 2455 4607
rect 2697 4573 2731 4607
rect 4169 4573 4203 4607
rect 3433 4437 3467 4471
rect 4353 4233 4387 4267
rect 3617 4097 3651 4131
rect 3341 4029 3375 4063
rect 3617 3009 3651 3043
rect 3341 2941 3375 2975
rect 4353 2805 4387 2839
rect 2513 1989 2547 2023
rect 2053 1921 2087 1955
rect 3709 1921 3743 1955
rect 3985 1853 4019 1887
rect 2973 1309 3007 1343
rect 3249 1241 3283 1275
<< metal1 >>
rect 1104 22874 5035 22896
rect 1104 22822 1892 22874
rect 1944 22822 1956 22874
rect 2008 22822 2020 22874
rect 2072 22822 2084 22874
rect 2136 22822 2148 22874
rect 2200 22822 2835 22874
rect 2887 22822 2899 22874
rect 2951 22822 2963 22874
rect 3015 22822 3027 22874
rect 3079 22822 3091 22874
rect 3143 22822 3778 22874
rect 3830 22822 3842 22874
rect 3894 22822 3906 22874
rect 3958 22822 3970 22874
rect 4022 22822 4034 22874
rect 4086 22822 4721 22874
rect 4773 22822 4785 22874
rect 4837 22822 4849 22874
rect 4901 22822 4913 22874
rect 4965 22822 4977 22874
rect 5029 22822 5035 22874
rect 1104 22800 5035 22822
rect 1104 22330 4876 22352
rect 1104 22278 1421 22330
rect 1473 22278 1485 22330
rect 1537 22278 1549 22330
rect 1601 22278 1613 22330
rect 1665 22278 1677 22330
rect 1729 22278 2364 22330
rect 2416 22278 2428 22330
rect 2480 22278 2492 22330
rect 2544 22278 2556 22330
rect 2608 22278 2620 22330
rect 2672 22278 3307 22330
rect 3359 22278 3371 22330
rect 3423 22278 3435 22330
rect 3487 22278 3499 22330
rect 3551 22278 3563 22330
rect 3615 22278 4250 22330
rect 4302 22278 4314 22330
rect 4366 22278 4378 22330
rect 4430 22278 4442 22330
rect 4494 22278 4506 22330
rect 4558 22278 4876 22330
rect 1104 22256 4876 22278
rect 1104 21786 5035 21808
rect 1104 21734 1892 21786
rect 1944 21734 1956 21786
rect 2008 21734 2020 21786
rect 2072 21734 2084 21786
rect 2136 21734 2148 21786
rect 2200 21734 2835 21786
rect 2887 21734 2899 21786
rect 2951 21734 2963 21786
rect 3015 21734 3027 21786
rect 3079 21734 3091 21786
rect 3143 21734 3778 21786
rect 3830 21734 3842 21786
rect 3894 21734 3906 21786
rect 3958 21734 3970 21786
rect 4022 21734 4034 21786
rect 4086 21734 4721 21786
rect 4773 21734 4785 21786
rect 4837 21734 4849 21786
rect 4901 21734 4913 21786
rect 4965 21734 4977 21786
rect 5029 21734 5035 21786
rect 1104 21712 5035 21734
rect 1104 21242 4876 21264
rect 1104 21190 1421 21242
rect 1473 21190 1485 21242
rect 1537 21190 1549 21242
rect 1601 21190 1613 21242
rect 1665 21190 1677 21242
rect 1729 21190 2364 21242
rect 2416 21190 2428 21242
rect 2480 21190 2492 21242
rect 2544 21190 2556 21242
rect 2608 21190 2620 21242
rect 2672 21190 3307 21242
rect 3359 21190 3371 21242
rect 3423 21190 3435 21242
rect 3487 21190 3499 21242
rect 3551 21190 3563 21242
rect 3615 21190 4250 21242
rect 4302 21190 4314 21242
rect 4366 21190 4378 21242
rect 4430 21190 4442 21242
rect 4494 21190 4506 21242
rect 4558 21190 4876 21242
rect 1104 21168 4876 21190
rect 1104 20698 5035 20720
rect 1104 20646 1892 20698
rect 1944 20646 1956 20698
rect 2008 20646 2020 20698
rect 2072 20646 2084 20698
rect 2136 20646 2148 20698
rect 2200 20646 2835 20698
rect 2887 20646 2899 20698
rect 2951 20646 2963 20698
rect 3015 20646 3027 20698
rect 3079 20646 3091 20698
rect 3143 20646 3778 20698
rect 3830 20646 3842 20698
rect 3894 20646 3906 20698
rect 3958 20646 3970 20698
rect 4022 20646 4034 20698
rect 4086 20646 4721 20698
rect 4773 20646 4785 20698
rect 4837 20646 4849 20698
rect 4901 20646 4913 20698
rect 4965 20646 4977 20698
rect 5029 20646 5035 20698
rect 1104 20624 5035 20646
rect 1104 20154 4876 20176
rect 1104 20102 1421 20154
rect 1473 20102 1485 20154
rect 1537 20102 1549 20154
rect 1601 20102 1613 20154
rect 1665 20102 1677 20154
rect 1729 20102 2364 20154
rect 2416 20102 2428 20154
rect 2480 20102 2492 20154
rect 2544 20102 2556 20154
rect 2608 20102 2620 20154
rect 2672 20102 3307 20154
rect 3359 20102 3371 20154
rect 3423 20102 3435 20154
rect 3487 20102 3499 20154
rect 3551 20102 3563 20154
rect 3615 20102 4250 20154
rect 4302 20102 4314 20154
rect 4366 20102 4378 20154
rect 4430 20102 4442 20154
rect 4494 20102 4506 20154
rect 4558 20102 4876 20154
rect 1104 20080 4876 20102
rect 1104 19610 5035 19632
rect 1104 19558 1892 19610
rect 1944 19558 1956 19610
rect 2008 19558 2020 19610
rect 2072 19558 2084 19610
rect 2136 19558 2148 19610
rect 2200 19558 2835 19610
rect 2887 19558 2899 19610
rect 2951 19558 2963 19610
rect 3015 19558 3027 19610
rect 3079 19558 3091 19610
rect 3143 19558 3778 19610
rect 3830 19558 3842 19610
rect 3894 19558 3906 19610
rect 3958 19558 3970 19610
rect 4022 19558 4034 19610
rect 4086 19558 4721 19610
rect 4773 19558 4785 19610
rect 4837 19558 4849 19610
rect 4901 19558 4913 19610
rect 4965 19558 4977 19610
rect 5029 19558 5035 19610
rect 1104 19536 5035 19558
rect 1104 19066 4876 19088
rect 1104 19014 1421 19066
rect 1473 19014 1485 19066
rect 1537 19014 1549 19066
rect 1601 19014 1613 19066
rect 1665 19014 1677 19066
rect 1729 19014 2364 19066
rect 2416 19014 2428 19066
rect 2480 19014 2492 19066
rect 2544 19014 2556 19066
rect 2608 19014 2620 19066
rect 2672 19014 3307 19066
rect 3359 19014 3371 19066
rect 3423 19014 3435 19066
rect 3487 19014 3499 19066
rect 3551 19014 3563 19066
rect 3615 19014 4250 19066
rect 4302 19014 4314 19066
rect 4366 19014 4378 19066
rect 4430 19014 4442 19066
rect 4494 19014 4506 19066
rect 4558 19014 4876 19066
rect 1104 18992 4876 19014
rect 1104 18522 5035 18544
rect 1104 18470 1892 18522
rect 1944 18470 1956 18522
rect 2008 18470 2020 18522
rect 2072 18470 2084 18522
rect 2136 18470 2148 18522
rect 2200 18470 2835 18522
rect 2887 18470 2899 18522
rect 2951 18470 2963 18522
rect 3015 18470 3027 18522
rect 3079 18470 3091 18522
rect 3143 18470 3778 18522
rect 3830 18470 3842 18522
rect 3894 18470 3906 18522
rect 3958 18470 3970 18522
rect 4022 18470 4034 18522
rect 4086 18470 4721 18522
rect 4773 18470 4785 18522
rect 4837 18470 4849 18522
rect 4901 18470 4913 18522
rect 4965 18470 4977 18522
rect 5029 18470 5035 18522
rect 1104 18448 5035 18470
rect 1104 17978 4876 18000
rect 1104 17926 1421 17978
rect 1473 17926 1485 17978
rect 1537 17926 1549 17978
rect 1601 17926 1613 17978
rect 1665 17926 1677 17978
rect 1729 17926 2364 17978
rect 2416 17926 2428 17978
rect 2480 17926 2492 17978
rect 2544 17926 2556 17978
rect 2608 17926 2620 17978
rect 2672 17926 3307 17978
rect 3359 17926 3371 17978
rect 3423 17926 3435 17978
rect 3487 17926 3499 17978
rect 3551 17926 3563 17978
rect 3615 17926 4250 17978
rect 4302 17926 4314 17978
rect 4366 17926 4378 17978
rect 4430 17926 4442 17978
rect 4494 17926 4506 17978
rect 4558 17926 4876 17978
rect 1104 17904 4876 17926
rect 1104 17434 5035 17456
rect 1104 17382 1892 17434
rect 1944 17382 1956 17434
rect 2008 17382 2020 17434
rect 2072 17382 2084 17434
rect 2136 17382 2148 17434
rect 2200 17382 2835 17434
rect 2887 17382 2899 17434
rect 2951 17382 2963 17434
rect 3015 17382 3027 17434
rect 3079 17382 3091 17434
rect 3143 17382 3778 17434
rect 3830 17382 3842 17434
rect 3894 17382 3906 17434
rect 3958 17382 3970 17434
rect 4022 17382 4034 17434
rect 4086 17382 4721 17434
rect 4773 17382 4785 17434
rect 4837 17382 4849 17434
rect 4901 17382 4913 17434
rect 4965 17382 4977 17434
rect 5029 17382 5035 17434
rect 1104 17360 5035 17382
rect 1104 16890 4876 16912
rect 1104 16838 1421 16890
rect 1473 16838 1485 16890
rect 1537 16838 1549 16890
rect 1601 16838 1613 16890
rect 1665 16838 1677 16890
rect 1729 16838 2364 16890
rect 2416 16838 2428 16890
rect 2480 16838 2492 16890
rect 2544 16838 2556 16890
rect 2608 16838 2620 16890
rect 2672 16838 3307 16890
rect 3359 16838 3371 16890
rect 3423 16838 3435 16890
rect 3487 16838 3499 16890
rect 3551 16838 3563 16890
rect 3615 16838 4250 16890
rect 4302 16838 4314 16890
rect 4366 16838 4378 16890
rect 4430 16838 4442 16890
rect 4494 16838 4506 16890
rect 4558 16838 4876 16890
rect 1104 16816 4876 16838
rect 1104 16346 5035 16368
rect 1104 16294 1892 16346
rect 1944 16294 1956 16346
rect 2008 16294 2020 16346
rect 2072 16294 2084 16346
rect 2136 16294 2148 16346
rect 2200 16294 2835 16346
rect 2887 16294 2899 16346
rect 2951 16294 2963 16346
rect 3015 16294 3027 16346
rect 3079 16294 3091 16346
rect 3143 16294 3778 16346
rect 3830 16294 3842 16346
rect 3894 16294 3906 16346
rect 3958 16294 3970 16346
rect 4022 16294 4034 16346
rect 4086 16294 4721 16346
rect 4773 16294 4785 16346
rect 4837 16294 4849 16346
rect 4901 16294 4913 16346
rect 4965 16294 4977 16346
rect 5029 16294 5035 16346
rect 1104 16272 5035 16294
rect 1104 15802 4876 15824
rect 1104 15750 1421 15802
rect 1473 15750 1485 15802
rect 1537 15750 1549 15802
rect 1601 15750 1613 15802
rect 1665 15750 1677 15802
rect 1729 15750 2364 15802
rect 2416 15750 2428 15802
rect 2480 15750 2492 15802
rect 2544 15750 2556 15802
rect 2608 15750 2620 15802
rect 2672 15750 3307 15802
rect 3359 15750 3371 15802
rect 3423 15750 3435 15802
rect 3487 15750 3499 15802
rect 3551 15750 3563 15802
rect 3615 15750 4250 15802
rect 4302 15750 4314 15802
rect 4366 15750 4378 15802
rect 4430 15750 4442 15802
rect 4494 15750 4506 15802
rect 4558 15750 4876 15802
rect 1104 15728 4876 15750
rect 1104 15258 5035 15280
rect 1104 15206 1892 15258
rect 1944 15206 1956 15258
rect 2008 15206 2020 15258
rect 2072 15206 2084 15258
rect 2136 15206 2148 15258
rect 2200 15206 2835 15258
rect 2887 15206 2899 15258
rect 2951 15206 2963 15258
rect 3015 15206 3027 15258
rect 3079 15206 3091 15258
rect 3143 15206 3778 15258
rect 3830 15206 3842 15258
rect 3894 15206 3906 15258
rect 3958 15206 3970 15258
rect 4022 15206 4034 15258
rect 4086 15206 4721 15258
rect 4773 15206 4785 15258
rect 4837 15206 4849 15258
rect 4901 15206 4913 15258
rect 4965 15206 4977 15258
rect 5029 15206 5035 15258
rect 1104 15184 5035 15206
rect 1104 14714 4876 14736
rect 1104 14662 1421 14714
rect 1473 14662 1485 14714
rect 1537 14662 1549 14714
rect 1601 14662 1613 14714
rect 1665 14662 1677 14714
rect 1729 14662 2364 14714
rect 2416 14662 2428 14714
rect 2480 14662 2492 14714
rect 2544 14662 2556 14714
rect 2608 14662 2620 14714
rect 2672 14662 3307 14714
rect 3359 14662 3371 14714
rect 3423 14662 3435 14714
rect 3487 14662 3499 14714
rect 3551 14662 3563 14714
rect 3615 14662 4250 14714
rect 4302 14662 4314 14714
rect 4366 14662 4378 14714
rect 4430 14662 4442 14714
rect 4494 14662 4506 14714
rect 4558 14662 4876 14714
rect 1104 14640 4876 14662
rect 1104 14170 5035 14192
rect 1104 14118 1892 14170
rect 1944 14118 1956 14170
rect 2008 14118 2020 14170
rect 2072 14118 2084 14170
rect 2136 14118 2148 14170
rect 2200 14118 2835 14170
rect 2887 14118 2899 14170
rect 2951 14118 2963 14170
rect 3015 14118 3027 14170
rect 3079 14118 3091 14170
rect 3143 14118 3778 14170
rect 3830 14118 3842 14170
rect 3894 14118 3906 14170
rect 3958 14118 3970 14170
rect 4022 14118 4034 14170
rect 4086 14118 4721 14170
rect 4773 14118 4785 14170
rect 4837 14118 4849 14170
rect 4901 14118 4913 14170
rect 4965 14118 4977 14170
rect 5029 14118 5035 14170
rect 1104 14096 5035 14118
rect 1104 13626 4876 13648
rect 1104 13574 1421 13626
rect 1473 13574 1485 13626
rect 1537 13574 1549 13626
rect 1601 13574 1613 13626
rect 1665 13574 1677 13626
rect 1729 13574 2364 13626
rect 2416 13574 2428 13626
rect 2480 13574 2492 13626
rect 2544 13574 2556 13626
rect 2608 13574 2620 13626
rect 2672 13574 3307 13626
rect 3359 13574 3371 13626
rect 3423 13574 3435 13626
rect 3487 13574 3499 13626
rect 3551 13574 3563 13626
rect 3615 13574 4250 13626
rect 4302 13574 4314 13626
rect 4366 13574 4378 13626
rect 4430 13574 4442 13626
rect 4494 13574 4506 13626
rect 4558 13574 4876 13626
rect 1104 13552 4876 13574
rect 1104 13082 5035 13104
rect 1104 13030 1892 13082
rect 1944 13030 1956 13082
rect 2008 13030 2020 13082
rect 2072 13030 2084 13082
rect 2136 13030 2148 13082
rect 2200 13030 2835 13082
rect 2887 13030 2899 13082
rect 2951 13030 2963 13082
rect 3015 13030 3027 13082
rect 3079 13030 3091 13082
rect 3143 13030 3778 13082
rect 3830 13030 3842 13082
rect 3894 13030 3906 13082
rect 3958 13030 3970 13082
rect 4022 13030 4034 13082
rect 4086 13030 4721 13082
rect 4773 13030 4785 13082
rect 4837 13030 4849 13082
rect 4901 13030 4913 13082
rect 4965 13030 4977 13082
rect 5029 13030 5035 13082
rect 1104 13008 5035 13030
rect 1104 12538 4876 12560
rect 1104 12486 1421 12538
rect 1473 12486 1485 12538
rect 1537 12486 1549 12538
rect 1601 12486 1613 12538
rect 1665 12486 1677 12538
rect 1729 12486 2364 12538
rect 2416 12486 2428 12538
rect 2480 12486 2492 12538
rect 2544 12486 2556 12538
rect 2608 12486 2620 12538
rect 2672 12486 3307 12538
rect 3359 12486 3371 12538
rect 3423 12486 3435 12538
rect 3487 12486 3499 12538
rect 3551 12486 3563 12538
rect 3615 12486 4250 12538
rect 4302 12486 4314 12538
rect 4366 12486 4378 12538
rect 4430 12486 4442 12538
rect 4494 12486 4506 12538
rect 4558 12486 4876 12538
rect 1104 12464 4876 12486
rect 1104 11994 5035 12016
rect 1104 11942 1892 11994
rect 1944 11942 1956 11994
rect 2008 11942 2020 11994
rect 2072 11942 2084 11994
rect 2136 11942 2148 11994
rect 2200 11942 2835 11994
rect 2887 11942 2899 11994
rect 2951 11942 2963 11994
rect 3015 11942 3027 11994
rect 3079 11942 3091 11994
rect 3143 11942 3778 11994
rect 3830 11942 3842 11994
rect 3894 11942 3906 11994
rect 3958 11942 3970 11994
rect 4022 11942 4034 11994
rect 4086 11942 4721 11994
rect 4773 11942 4785 11994
rect 4837 11942 4849 11994
rect 4901 11942 4913 11994
rect 4965 11942 4977 11994
rect 5029 11942 5035 11994
rect 1104 11920 5035 11942
rect 3142 11840 3148 11892
rect 3200 11880 3206 11892
rect 3874 11883 3932 11889
rect 3874 11880 3886 11883
rect 3200 11852 3886 11880
rect 3200 11840 3206 11852
rect 3874 11849 3886 11852
rect 3920 11849 3932 11883
rect 3874 11843 3932 11849
rect 3605 11747 3663 11753
rect 3605 11713 3617 11747
rect 3651 11744 3663 11747
rect 5074 11744 5080 11756
rect 3651 11716 5080 11744
rect 3651 11713 3663 11716
rect 3605 11707 3663 11713
rect 5074 11704 5080 11716
rect 5132 11704 5138 11756
rect 3878 11676 3884 11688
rect 3839 11648 3884 11676
rect 3878 11636 3884 11648
rect 3936 11636 3942 11688
rect 4154 11636 4160 11688
rect 4212 11676 4218 11688
rect 4341 11679 4399 11685
rect 4341 11676 4353 11679
rect 4212 11648 4353 11676
rect 4212 11636 4218 11648
rect 4341 11645 4353 11648
rect 4387 11645 4399 11679
rect 4341 11639 4399 11645
rect 1762 11500 1768 11552
rect 1820 11540 1826 11552
rect 2501 11543 2559 11549
rect 2501 11540 2513 11543
rect 1820 11512 2513 11540
rect 1820 11500 1826 11512
rect 2501 11509 2513 11512
rect 2547 11509 2559 11543
rect 2501 11503 2559 11509
rect 3878 11500 3884 11552
rect 3936 11540 3942 11552
rect 5074 11540 5080 11552
rect 3936 11512 5080 11540
rect 3936 11500 3942 11512
rect 5074 11500 5080 11512
rect 5132 11500 5138 11552
rect 1104 11450 4876 11472
rect 1104 11398 1421 11450
rect 1473 11398 1485 11450
rect 1537 11398 1549 11450
rect 1601 11398 1613 11450
rect 1665 11398 1677 11450
rect 1729 11398 2364 11450
rect 2416 11398 2428 11450
rect 2480 11398 2492 11450
rect 2544 11398 2556 11450
rect 2608 11398 2620 11450
rect 2672 11398 3307 11450
rect 3359 11398 3371 11450
rect 3423 11398 3435 11450
rect 3487 11398 3499 11450
rect 3551 11398 3563 11450
rect 3615 11398 4250 11450
rect 4302 11398 4314 11450
rect 4366 11398 4378 11450
rect 4430 11398 4442 11450
rect 4494 11398 4506 11450
rect 4558 11398 4876 11450
rect 1104 11376 4876 11398
rect 3418 11228 3424 11280
rect 3476 11228 3482 11280
rect 1210 11092 1216 11144
rect 1268 11132 1274 11144
rect 2409 11135 2467 11141
rect 2409 11132 2421 11135
rect 1268 11104 2421 11132
rect 1268 11092 1274 11104
rect 2409 11101 2421 11104
rect 2455 11101 2467 11135
rect 2409 11095 2467 11101
rect 2682 11092 2688 11144
rect 2740 11092 2746 11144
rect 1104 10906 5035 10928
rect 1104 10854 1892 10906
rect 1944 10854 1956 10906
rect 2008 10854 2020 10906
rect 2072 10854 2084 10906
rect 2136 10854 2148 10906
rect 2200 10854 2835 10906
rect 2887 10854 2899 10906
rect 2951 10854 2963 10906
rect 3015 10854 3027 10906
rect 3079 10854 3091 10906
rect 3143 10854 3778 10906
rect 3830 10854 3842 10906
rect 3894 10854 3906 10906
rect 3958 10854 3970 10906
rect 4022 10854 4034 10906
rect 4086 10854 4721 10906
rect 4773 10854 4785 10906
rect 4837 10854 4849 10906
rect 4901 10854 4913 10906
rect 4965 10854 4977 10906
rect 5029 10854 5035 10906
rect 1104 10832 5035 10854
rect 2222 10752 2228 10804
rect 2280 10792 2286 10804
rect 3234 10792 3240 10804
rect 2280 10764 3240 10792
rect 2280 10752 2286 10764
rect 3234 10752 3240 10764
rect 3292 10792 3298 10804
rect 3874 10795 3932 10801
rect 3874 10792 3886 10795
rect 3292 10764 3886 10792
rect 3292 10752 3298 10764
rect 3874 10761 3886 10764
rect 3920 10761 3932 10795
rect 3874 10755 3932 10761
rect 3605 10659 3663 10665
rect 3605 10625 3617 10659
rect 3651 10656 3663 10659
rect 5166 10656 5172 10668
rect 3651 10628 5172 10656
rect 3651 10625 3663 10628
rect 3605 10619 3663 10625
rect 5166 10616 5172 10628
rect 5224 10616 5230 10668
rect 3878 10588 3884 10600
rect 3839 10560 3884 10588
rect 3878 10548 3884 10560
rect 3936 10548 3942 10600
rect 4154 10548 4160 10600
rect 4212 10588 4218 10600
rect 4341 10591 4399 10597
rect 4341 10588 4353 10591
rect 4212 10560 4353 10588
rect 4212 10548 4218 10560
rect 4341 10557 4353 10560
rect 4387 10557 4399 10591
rect 4341 10551 4399 10557
rect 2501 10455 2559 10461
rect 2501 10421 2513 10455
rect 2547 10452 2559 10455
rect 3142 10452 3148 10464
rect 2547 10424 3148 10452
rect 2547 10421 2559 10424
rect 2501 10415 2559 10421
rect 3142 10412 3148 10424
rect 3200 10412 3206 10464
rect 1104 10362 4876 10384
rect 1104 10310 1421 10362
rect 1473 10310 1485 10362
rect 1537 10310 1549 10362
rect 1601 10310 1613 10362
rect 1665 10310 1677 10362
rect 1729 10310 2364 10362
rect 2416 10310 2428 10362
rect 2480 10310 2492 10362
rect 2544 10310 2556 10362
rect 2608 10310 2620 10362
rect 2672 10310 3307 10362
rect 3359 10310 3371 10362
rect 3423 10310 3435 10362
rect 3487 10310 3499 10362
rect 3551 10310 3563 10362
rect 3615 10310 4250 10362
rect 4302 10310 4314 10362
rect 4366 10310 4378 10362
rect 4430 10310 4442 10362
rect 4494 10310 4506 10362
rect 4558 10310 4876 10362
rect 1104 10288 4876 10310
rect 1302 10072 1308 10124
rect 1360 10112 1366 10124
rect 2044 10115 2102 10121
rect 2044 10112 2056 10115
rect 1360 10084 2056 10112
rect 1360 10072 1366 10084
rect 2044 10081 2056 10084
rect 2090 10081 2102 10115
rect 2044 10075 2102 10081
rect 2317 10115 2375 10121
rect 2317 10081 2329 10115
rect 2363 10112 2375 10115
rect 5534 10112 5540 10124
rect 2363 10084 5540 10112
rect 2363 10081 2375 10084
rect 2317 10075 2375 10081
rect 5534 10072 5540 10084
rect 5592 10072 5598 10124
rect 1118 10004 1124 10056
rect 1176 10044 1182 10056
rect 1581 10047 1639 10053
rect 1581 10044 1593 10047
rect 1176 10016 1593 10044
rect 1176 10004 1182 10016
rect 1581 10013 1593 10016
rect 1627 10013 1639 10047
rect 1581 10007 1639 10013
rect 3602 9936 3608 9988
rect 3660 9976 3666 9988
rect 5258 9976 5264 9988
rect 3660 9948 5264 9976
rect 3660 9936 3666 9948
rect 5258 9936 5264 9948
rect 5316 9936 5322 9988
rect 2047 9911 2105 9917
rect 2047 9877 2059 9911
rect 2093 9908 2105 9911
rect 2222 9908 2228 9920
rect 2093 9880 2228 9908
rect 2093 9877 2105 9880
rect 2047 9871 2105 9877
rect 2222 9868 2228 9880
rect 2280 9868 2286 9920
rect 3421 9911 3479 9917
rect 3421 9877 3433 9911
rect 3467 9908 3479 9911
rect 3878 9908 3884 9920
rect 3467 9880 3884 9908
rect 3467 9877 3479 9880
rect 3421 9871 3479 9877
rect 3878 9868 3884 9880
rect 3936 9908 3942 9920
rect 4614 9908 4620 9920
rect 3936 9880 4620 9908
rect 3936 9868 3942 9880
rect 4614 9868 4620 9880
rect 4672 9868 4678 9920
rect 1104 9818 5035 9840
rect 1104 9766 1892 9818
rect 1944 9766 1956 9818
rect 2008 9766 2020 9818
rect 2072 9766 2084 9818
rect 2136 9766 2148 9818
rect 2200 9766 2835 9818
rect 2887 9766 2899 9818
rect 2951 9766 2963 9818
rect 3015 9766 3027 9818
rect 3079 9766 3091 9818
rect 3143 9766 3778 9818
rect 3830 9766 3842 9818
rect 3894 9766 3906 9818
rect 3958 9766 3970 9818
rect 4022 9766 4034 9818
rect 4086 9766 4721 9818
rect 4773 9766 4785 9818
rect 4837 9766 4849 9818
rect 4901 9766 4913 9818
rect 4965 9766 4977 9818
rect 5029 9766 5035 9818
rect 1104 9744 5035 9766
rect 3878 9713 3884 9716
rect 3874 9667 3884 9713
rect 3936 9704 3942 9716
rect 3936 9676 3974 9704
rect 3878 9664 3884 9667
rect 3936 9664 3942 9676
rect 3234 9528 3240 9580
rect 3292 9568 3298 9580
rect 3292 9540 3740 9568
rect 3292 9528 3298 9540
rect 3602 9460 3608 9512
rect 3660 9460 3666 9512
rect 3712 9500 3740 9540
rect 3835 9503 3893 9509
rect 3835 9500 3847 9503
rect 3712 9472 3847 9500
rect 3835 9469 3847 9472
rect 3881 9469 3893 9503
rect 3835 9463 3893 9469
rect 4154 9460 4160 9512
rect 4212 9500 4218 9512
rect 4341 9503 4399 9509
rect 4341 9500 4353 9503
rect 4212 9472 4353 9500
rect 4212 9460 4218 9472
rect 4341 9469 4353 9472
rect 4387 9469 4399 9503
rect 4341 9463 4399 9469
rect 2501 9367 2559 9373
rect 2501 9333 2513 9367
rect 2547 9364 2559 9367
rect 2682 9364 2688 9376
rect 2547 9336 2688 9364
rect 2547 9333 2559 9336
rect 2501 9327 2559 9333
rect 2682 9324 2688 9336
rect 2740 9324 2746 9376
rect 3786 9324 3792 9376
rect 3844 9364 3850 9376
rect 4522 9364 4528 9376
rect 3844 9336 4528 9364
rect 3844 9324 3850 9336
rect 4522 9324 4528 9336
rect 4580 9324 4586 9376
rect 1104 9274 4876 9296
rect 1104 9222 1421 9274
rect 1473 9222 1485 9274
rect 1537 9222 1549 9274
rect 1601 9222 1613 9274
rect 1665 9222 1677 9274
rect 1729 9222 2364 9274
rect 2416 9222 2428 9274
rect 2480 9222 2492 9274
rect 2544 9222 2556 9274
rect 2608 9222 2620 9274
rect 2672 9222 3307 9274
rect 3359 9222 3371 9274
rect 3423 9222 3435 9274
rect 3487 9222 3499 9274
rect 3551 9222 3563 9274
rect 3615 9222 4250 9274
rect 4302 9222 4314 9274
rect 4366 9222 4378 9274
rect 4430 9222 4442 9274
rect 4494 9222 4506 9274
rect 4558 9222 4876 9274
rect 1104 9200 4876 9222
rect 1762 9120 1768 9172
rect 1820 9160 1826 9172
rect 3510 9160 3516 9172
rect 1820 9132 3516 9160
rect 1820 9120 1826 9132
rect 3510 9120 3516 9132
rect 3568 9120 3574 9172
rect 3602 9120 3608 9172
rect 3660 9160 3666 9172
rect 3878 9160 3884 9172
rect 3660 9132 3884 9160
rect 3660 9120 3666 9132
rect 3878 9120 3884 9132
rect 3936 9120 3942 9172
rect 2038 8984 2044 9036
rect 2096 8984 2102 9036
rect 2317 9027 2375 9033
rect 2317 8993 2329 9027
rect 2363 9024 2375 9027
rect 3694 9024 3700 9036
rect 2363 8996 3700 9024
rect 2363 8993 2375 8996
rect 2317 8987 2375 8993
rect 3694 8984 3700 8996
rect 3752 8984 3758 9036
rect 1118 8916 1124 8968
rect 1176 8956 1182 8968
rect 1581 8959 1639 8965
rect 1581 8956 1593 8959
rect 1176 8928 1593 8956
rect 1176 8916 1182 8928
rect 1581 8925 1593 8928
rect 1627 8925 1639 8959
rect 1581 8919 1639 8925
rect 1670 8780 1676 8832
rect 1728 8820 1734 8832
rect 2047 8823 2105 8829
rect 2047 8820 2059 8823
rect 1728 8792 2059 8820
rect 1728 8780 1734 8792
rect 2047 8789 2059 8792
rect 2093 8789 2105 8823
rect 2047 8783 2105 8789
rect 3421 8823 3479 8829
rect 3421 8789 3433 8823
rect 3467 8820 3479 8823
rect 5074 8820 5080 8832
rect 3467 8792 5080 8820
rect 3467 8789 3479 8792
rect 3421 8783 3479 8789
rect 5074 8780 5080 8792
rect 5132 8820 5138 8832
rect 5258 8820 5264 8832
rect 5132 8792 5264 8820
rect 5132 8780 5138 8792
rect 5258 8780 5264 8792
rect 5316 8780 5322 8832
rect 1104 8730 5035 8752
rect 1104 8678 1892 8730
rect 1944 8678 1956 8730
rect 2008 8678 2020 8730
rect 2072 8678 2084 8730
rect 2136 8678 2148 8730
rect 2200 8678 2835 8730
rect 2887 8678 2899 8730
rect 2951 8678 2963 8730
rect 3015 8678 3027 8730
rect 3079 8678 3091 8730
rect 3143 8678 3778 8730
rect 3830 8678 3842 8730
rect 3894 8678 3906 8730
rect 3958 8678 3970 8730
rect 4022 8678 4034 8730
rect 4086 8678 4721 8730
rect 4773 8678 4785 8730
rect 4837 8678 4849 8730
rect 4901 8678 4913 8730
rect 4965 8678 4977 8730
rect 5029 8678 5035 8730
rect 1104 8656 5035 8678
rect 1670 8576 1676 8628
rect 1728 8616 1734 8628
rect 2130 8616 2136 8628
rect 1728 8588 2136 8616
rect 1728 8576 1734 8588
rect 2130 8576 2136 8588
rect 2188 8616 2194 8628
rect 3602 8616 3608 8628
rect 2188 8588 3608 8616
rect 2188 8576 2194 8588
rect 3602 8576 3608 8588
rect 3660 8616 3666 8628
rect 3874 8619 3932 8625
rect 3874 8616 3886 8619
rect 3660 8588 3886 8616
rect 3660 8576 3666 8588
rect 3874 8585 3886 8588
rect 3920 8585 3932 8619
rect 3874 8579 3932 8585
rect 3605 8483 3663 8489
rect 3605 8449 3617 8483
rect 3651 8480 3663 8483
rect 3694 8480 3700 8492
rect 3651 8452 3700 8480
rect 3651 8449 3663 8452
rect 3605 8443 3663 8449
rect 3694 8440 3700 8452
rect 3752 8440 3758 8492
rect 5534 8480 5540 8492
rect 3804 8452 5540 8480
rect 3510 8372 3516 8424
rect 3568 8412 3574 8424
rect 3804 8414 3832 8452
rect 5534 8440 5540 8452
rect 5592 8440 5598 8492
rect 3862 8417 3920 8423
rect 3862 8414 3874 8417
rect 3804 8412 3874 8414
rect 3568 8386 3874 8412
rect 3568 8384 3832 8386
rect 3568 8372 3574 8384
rect 3862 8383 3874 8386
rect 3908 8383 3920 8417
rect 3862 8377 3920 8383
rect 4154 8372 4160 8424
rect 4212 8412 4218 8424
rect 4341 8415 4399 8421
rect 4341 8412 4353 8415
rect 4212 8384 4353 8412
rect 4212 8372 4218 8384
rect 4341 8381 4353 8384
rect 4387 8381 4399 8415
rect 4341 8375 4399 8381
rect 1302 8236 1308 8288
rect 1360 8276 1366 8288
rect 2501 8279 2559 8285
rect 2501 8276 2513 8279
rect 1360 8248 2513 8276
rect 1360 8236 1366 8248
rect 2501 8245 2513 8248
rect 2547 8245 2559 8279
rect 2501 8239 2559 8245
rect 1104 8186 4876 8208
rect 1104 8134 1421 8186
rect 1473 8134 1485 8186
rect 1537 8134 1549 8186
rect 1601 8134 1613 8186
rect 1665 8134 1677 8186
rect 1729 8134 2364 8186
rect 2416 8134 2428 8186
rect 2480 8134 2492 8186
rect 2544 8134 2556 8186
rect 2608 8134 2620 8186
rect 2672 8134 3307 8186
rect 3359 8134 3371 8186
rect 3423 8134 3435 8186
rect 3487 8134 3499 8186
rect 3551 8134 3563 8186
rect 3615 8134 4250 8186
rect 4302 8134 4314 8186
rect 4366 8134 4378 8186
rect 4430 8134 4442 8186
rect 4494 8134 4506 8186
rect 4558 8134 4876 8186
rect 1104 8112 4876 8134
rect 1854 7896 1860 7948
rect 1912 7918 1918 7948
rect 2317 7939 2375 7945
rect 2044 7921 2102 7927
rect 2044 7918 2056 7921
rect 1912 7896 2056 7918
rect 1872 7890 2056 7896
rect 2044 7887 2056 7890
rect 2090 7887 2102 7921
rect 2317 7905 2329 7939
rect 2363 7936 2375 7939
rect 5442 7936 5448 7948
rect 2363 7908 5448 7936
rect 2363 7905 2375 7908
rect 2317 7899 2375 7905
rect 5442 7896 5448 7908
rect 5500 7896 5506 7948
rect 2044 7881 2102 7887
rect 1118 7828 1124 7880
rect 1176 7868 1182 7880
rect 1578 7868 1584 7880
rect 1176 7840 1584 7868
rect 1176 7828 1182 7840
rect 1578 7828 1584 7840
rect 1636 7828 1642 7880
rect 1118 7692 1124 7744
rect 1176 7732 1182 7744
rect 1854 7732 1860 7744
rect 1176 7704 1860 7732
rect 1176 7692 1182 7704
rect 1854 7692 1860 7704
rect 1912 7692 1918 7744
rect 2038 7732 2044 7744
rect 2096 7741 2102 7744
rect 2005 7704 2044 7732
rect 2038 7692 2044 7704
rect 2096 7695 2105 7741
rect 3421 7735 3479 7741
rect 3421 7701 3433 7735
rect 3467 7732 3479 7735
rect 3694 7732 3700 7744
rect 3467 7704 3700 7732
rect 3467 7701 3479 7704
rect 3421 7695 3479 7701
rect 2096 7692 2102 7695
rect 3694 7692 3700 7704
rect 3752 7692 3758 7744
rect 1104 7642 5035 7664
rect 1104 7590 1892 7642
rect 1944 7590 1956 7642
rect 2008 7590 2020 7642
rect 2072 7590 2084 7642
rect 2136 7590 2148 7642
rect 2200 7590 2835 7642
rect 2887 7590 2899 7642
rect 2951 7590 2963 7642
rect 3015 7590 3027 7642
rect 3079 7590 3091 7642
rect 3143 7590 3778 7642
rect 3830 7590 3842 7642
rect 3894 7590 3906 7642
rect 3958 7590 3970 7642
rect 4022 7590 4034 7642
rect 4086 7590 4721 7642
rect 4773 7590 4785 7642
rect 4837 7590 4849 7642
rect 4901 7590 4913 7642
rect 4965 7590 4977 7642
rect 5029 7590 5035 7642
rect 1104 7568 5035 7590
rect 1762 7488 1768 7540
rect 1820 7528 1826 7540
rect 2501 7531 2559 7537
rect 2501 7528 2513 7531
rect 1820 7500 2513 7528
rect 1820 7488 1826 7500
rect 2501 7497 2513 7500
rect 2547 7497 2559 7531
rect 3874 7531 3932 7537
rect 3874 7528 3886 7531
rect 2501 7491 2559 7497
rect 2792 7500 3886 7528
rect 2792 7472 2820 7500
rect 3874 7497 3886 7500
rect 3920 7497 3932 7531
rect 3874 7491 3932 7497
rect 1578 7420 1584 7472
rect 1636 7460 1642 7472
rect 2222 7460 2228 7472
rect 1636 7432 2228 7460
rect 1636 7420 1642 7432
rect 2222 7420 2228 7432
rect 2280 7420 2286 7472
rect 2314 7420 2320 7472
rect 2372 7460 2378 7472
rect 2774 7460 2780 7472
rect 2372 7432 2780 7460
rect 2372 7420 2378 7432
rect 2774 7420 2780 7432
rect 2832 7420 2838 7472
rect 3605 7395 3663 7401
rect 3605 7361 3617 7395
rect 3651 7392 3663 7395
rect 5350 7392 5356 7404
rect 3651 7364 5356 7392
rect 3651 7361 3663 7364
rect 3605 7355 3663 7361
rect 5350 7352 5356 7364
rect 5408 7352 5414 7404
rect 3694 7284 3700 7336
rect 3752 7324 3758 7336
rect 3835 7327 3893 7333
rect 3835 7324 3847 7327
rect 3752 7296 3847 7324
rect 3752 7284 3758 7296
rect 3835 7293 3847 7296
rect 3881 7293 3893 7327
rect 3835 7287 3893 7293
rect 4154 7284 4160 7336
rect 4212 7324 4218 7336
rect 4341 7327 4399 7333
rect 4341 7324 4353 7327
rect 4212 7296 4353 7324
rect 4212 7284 4218 7296
rect 4341 7293 4353 7296
rect 4387 7293 4399 7327
rect 4341 7287 4399 7293
rect 1104 7098 4876 7120
rect 1104 7046 1421 7098
rect 1473 7046 1485 7098
rect 1537 7046 1549 7098
rect 1601 7046 1613 7098
rect 1665 7046 1677 7098
rect 1729 7046 2364 7098
rect 2416 7046 2428 7098
rect 2480 7046 2492 7098
rect 2544 7046 2556 7098
rect 2608 7046 2620 7098
rect 2672 7046 3307 7098
rect 3359 7046 3371 7098
rect 3423 7046 3435 7098
rect 3487 7046 3499 7098
rect 3551 7046 3563 7098
rect 3615 7046 4250 7098
rect 4302 7046 4314 7098
rect 4366 7046 4378 7098
rect 4430 7046 4442 7098
rect 4494 7046 4506 7098
rect 4558 7046 4876 7098
rect 1104 7024 4876 7046
rect 3421 6987 3479 6993
rect 3421 6953 3433 6987
rect 3467 6984 3479 6987
rect 5166 6984 5172 6996
rect 3467 6956 5172 6984
rect 3467 6953 3479 6956
rect 3421 6947 3479 6953
rect 5166 6944 5172 6956
rect 5224 6944 5230 6996
rect 1210 6808 1216 6860
rect 1268 6848 1274 6860
rect 2409 6851 2467 6857
rect 2409 6848 2421 6851
rect 1268 6820 2421 6848
rect 1268 6808 1274 6820
rect 2409 6817 2421 6820
rect 2455 6817 2467 6851
rect 2409 6811 2467 6817
rect 2685 6783 2743 6789
rect 2685 6749 2697 6783
rect 2731 6780 2743 6783
rect 3142 6780 3148 6792
rect 2731 6752 3148 6780
rect 2731 6749 2743 6752
rect 2685 6743 2743 6749
rect 3142 6740 3148 6752
rect 3200 6740 3206 6792
rect 2590 6672 2596 6724
rect 2648 6712 2654 6724
rect 2774 6712 2780 6724
rect 2648 6684 2780 6712
rect 2648 6672 2654 6684
rect 2774 6672 2780 6684
rect 2832 6672 2838 6724
rect 3694 6604 3700 6656
rect 3752 6644 3758 6656
rect 3973 6647 4031 6653
rect 3973 6644 3985 6647
rect 3752 6616 3985 6644
rect 3752 6604 3758 6616
rect 3973 6613 3985 6616
rect 4019 6613 4031 6647
rect 3973 6607 4031 6613
rect 1104 6554 5035 6576
rect 1104 6502 1892 6554
rect 1944 6502 1956 6554
rect 2008 6502 2020 6554
rect 2072 6502 2084 6554
rect 2136 6502 2148 6554
rect 2200 6502 2835 6554
rect 2887 6502 2899 6554
rect 2951 6502 2963 6554
rect 3015 6502 3027 6554
rect 3079 6502 3091 6554
rect 3143 6502 3778 6554
rect 3830 6502 3842 6554
rect 3894 6502 3906 6554
rect 3958 6502 3970 6554
rect 4022 6502 4034 6554
rect 4086 6502 4721 6554
rect 4773 6502 4785 6554
rect 4837 6502 4849 6554
rect 4901 6502 4913 6554
rect 4965 6502 4977 6554
rect 5029 6502 5035 6554
rect 1104 6480 5035 6502
rect 2593 6375 2651 6381
rect 2593 6341 2605 6375
rect 2639 6372 2651 6375
rect 2682 6372 2688 6384
rect 2639 6344 2688 6372
rect 2639 6341 2651 6344
rect 2593 6335 2651 6341
rect 2682 6332 2688 6344
rect 2740 6332 2746 6384
rect 3694 6264 3700 6316
rect 3752 6264 3758 6316
rect 2222 6196 2228 6248
rect 2280 6236 2286 6248
rect 2317 6239 2375 6245
rect 2317 6236 2329 6239
rect 2280 6208 2329 6236
rect 2280 6196 2286 6208
rect 2317 6205 2329 6208
rect 2363 6236 2375 6239
rect 4154 6236 4160 6248
rect 2363 6208 4160 6236
rect 2363 6205 2375 6208
rect 2317 6199 2375 6205
rect 4154 6196 4160 6208
rect 4212 6196 4218 6248
rect 4341 6239 4399 6245
rect 4341 6205 4353 6239
rect 4387 6236 4399 6239
rect 4614 6236 4620 6248
rect 4387 6208 4620 6236
rect 4387 6205 4399 6208
rect 4341 6199 4399 6205
rect 4614 6196 4620 6208
rect 4672 6196 4678 6248
rect 1762 6060 1768 6112
rect 1820 6100 1826 6112
rect 2222 6100 2228 6112
rect 1820 6072 2228 6100
rect 1820 6060 1826 6072
rect 2222 6060 2228 6072
rect 2280 6060 2286 6112
rect 1104 6010 4876 6032
rect 1104 5958 1421 6010
rect 1473 5958 1485 6010
rect 1537 5958 1549 6010
rect 1601 5958 1613 6010
rect 1665 5958 1677 6010
rect 1729 5958 2364 6010
rect 2416 5958 2428 6010
rect 2480 5958 2492 6010
rect 2544 5958 2556 6010
rect 2608 5958 2620 6010
rect 2672 5958 3307 6010
rect 3359 5958 3371 6010
rect 3423 5958 3435 6010
rect 3487 5958 3499 6010
rect 3551 5958 3563 6010
rect 3615 5958 4250 6010
rect 4302 5958 4314 6010
rect 4366 5958 4378 6010
rect 4430 5958 4442 6010
rect 4494 5958 4506 6010
rect 4558 5958 4876 6010
rect 1104 5936 4876 5958
rect 3421 5899 3479 5905
rect 3421 5865 3433 5899
rect 3467 5896 3479 5899
rect 3694 5896 3700 5908
rect 3467 5868 3700 5896
rect 3467 5865 3479 5868
rect 3421 5859 3479 5865
rect 3694 5856 3700 5868
rect 3752 5856 3758 5908
rect 3234 5788 3240 5840
rect 3292 5828 3298 5840
rect 4706 5828 4712 5840
rect 3292 5800 4712 5828
rect 3292 5788 3298 5800
rect 4706 5788 4712 5800
rect 4764 5788 4770 5840
rect 1210 5720 1216 5772
rect 1268 5760 1274 5772
rect 1762 5760 1768 5772
rect 1268 5732 1768 5760
rect 1268 5720 1274 5732
rect 1762 5720 1768 5732
rect 1820 5760 1826 5772
rect 2409 5763 2467 5769
rect 2409 5760 2421 5763
rect 1820 5732 2421 5760
rect 1820 5720 1826 5732
rect 2409 5729 2421 5732
rect 2455 5729 2467 5763
rect 2409 5723 2467 5729
rect 2685 5695 2743 5701
rect 2685 5661 2697 5695
rect 2731 5661 2743 5695
rect 2685 5655 2743 5661
rect 1302 5584 1308 5636
rect 1360 5624 1366 5636
rect 2700 5624 2728 5655
rect 1360 5596 2728 5624
rect 1360 5584 1366 5596
rect 1104 5466 5035 5488
rect 1104 5414 1892 5466
rect 1944 5414 1956 5466
rect 2008 5414 2020 5466
rect 2072 5414 2084 5466
rect 2136 5414 2148 5466
rect 2200 5414 2835 5466
rect 2887 5414 2899 5466
rect 2951 5414 2963 5466
rect 3015 5414 3027 5466
rect 3079 5414 3091 5466
rect 3143 5414 3778 5466
rect 3830 5414 3842 5466
rect 3894 5414 3906 5466
rect 3958 5414 3970 5466
rect 4022 5414 4034 5466
rect 4086 5414 4721 5466
rect 4773 5414 4785 5466
rect 4837 5414 4849 5466
rect 4901 5414 4913 5466
rect 4965 5414 4977 5466
rect 5029 5414 5035 5466
rect 1104 5392 5035 5414
rect 4341 5355 4399 5361
rect 4341 5321 4353 5355
rect 4387 5352 4399 5355
rect 5166 5352 5172 5364
rect 4387 5324 5172 5352
rect 4387 5321 4399 5324
rect 4341 5315 4399 5321
rect 5166 5312 5172 5324
rect 5224 5312 5230 5364
rect 2133 5219 2191 5225
rect 2133 5185 2145 5219
rect 2179 5216 2191 5219
rect 2222 5216 2228 5228
rect 2179 5188 2228 5216
rect 2179 5185 2191 5188
rect 2133 5179 2191 5185
rect 2222 5176 2228 5188
rect 2280 5176 2286 5228
rect 3234 5176 3240 5228
rect 3292 5216 3298 5228
rect 3605 5219 3663 5225
rect 3605 5216 3617 5219
rect 3292 5188 3617 5216
rect 3292 5176 3298 5188
rect 3605 5185 3617 5188
rect 3651 5185 3663 5219
rect 3605 5179 3663 5185
rect 1854 5108 1860 5160
rect 1912 5108 1918 5160
rect 3142 5108 3148 5160
rect 3200 5148 3206 5160
rect 3329 5151 3387 5157
rect 3329 5148 3341 5151
rect 3200 5120 3341 5148
rect 3200 5108 3206 5120
rect 3329 5117 3341 5120
rect 3375 5117 3387 5151
rect 3329 5111 3387 5117
rect 2682 4972 2688 5024
rect 2740 5012 2746 5024
rect 2869 5015 2927 5021
rect 2869 5012 2881 5015
rect 2740 4984 2881 5012
rect 2740 4972 2746 4984
rect 2869 4981 2881 4984
rect 2915 4981 2927 5015
rect 2869 4975 2927 4981
rect 1104 4922 4876 4944
rect 1104 4870 1421 4922
rect 1473 4870 1485 4922
rect 1537 4870 1549 4922
rect 1601 4870 1613 4922
rect 1665 4870 1677 4922
rect 1729 4870 2364 4922
rect 2416 4870 2428 4922
rect 2480 4870 2492 4922
rect 2544 4870 2556 4922
rect 2608 4870 2620 4922
rect 2672 4870 3307 4922
rect 3359 4870 3371 4922
rect 3423 4870 3435 4922
rect 3487 4870 3499 4922
rect 3551 4870 3563 4922
rect 3615 4870 4250 4922
rect 4302 4870 4314 4922
rect 4366 4870 4378 4922
rect 4430 4870 4442 4922
rect 4494 4870 4506 4922
rect 4558 4870 4876 4922
rect 1104 4848 4876 4870
rect 4154 4768 4160 4820
rect 4212 4808 4218 4820
rect 4249 4811 4307 4817
rect 4249 4808 4261 4811
rect 4212 4780 4261 4808
rect 4212 4768 4218 4780
rect 4249 4777 4261 4780
rect 4295 4777 4307 4811
rect 4249 4771 4307 4777
rect 5258 4672 5264 4684
rect 3988 4644 5264 4672
rect 1854 4564 1860 4616
rect 1912 4604 1918 4616
rect 2406 4604 2412 4616
rect 1912 4576 2412 4604
rect 1912 4564 1918 4576
rect 2406 4564 2412 4576
rect 2464 4564 2470 4616
rect 2685 4607 2743 4613
rect 2685 4573 2697 4607
rect 2731 4604 2743 4607
rect 3988 4604 4016 4644
rect 5258 4632 5264 4644
rect 5316 4632 5322 4684
rect 2731 4576 4016 4604
rect 2731 4573 2743 4576
rect 2685 4567 2743 4573
rect 4154 4564 4160 4616
rect 4212 4564 4218 4616
rect 3421 4471 3479 4477
rect 3421 4437 3433 4471
rect 3467 4468 3479 4471
rect 5166 4468 5172 4480
rect 3467 4440 5172 4468
rect 3467 4437 3479 4440
rect 3421 4431 3479 4437
rect 5166 4428 5172 4440
rect 5224 4428 5230 4480
rect 1104 4378 5035 4400
rect 1104 4326 1892 4378
rect 1944 4326 1956 4378
rect 2008 4326 2020 4378
rect 2072 4326 2084 4378
rect 2136 4326 2148 4378
rect 2200 4326 2835 4378
rect 2887 4326 2899 4378
rect 2951 4326 2963 4378
rect 3015 4326 3027 4378
rect 3079 4326 3091 4378
rect 3143 4326 3778 4378
rect 3830 4326 3842 4378
rect 3894 4326 3906 4378
rect 3958 4326 3970 4378
rect 4022 4326 4034 4378
rect 4086 4326 4721 4378
rect 4773 4326 4785 4378
rect 4837 4326 4849 4378
rect 4901 4326 4913 4378
rect 4965 4326 4977 4378
rect 5029 4326 5035 4378
rect 1104 4304 5035 4326
rect 4341 4267 4399 4273
rect 4341 4233 4353 4267
rect 4387 4264 4399 4267
rect 5074 4264 5080 4276
rect 4387 4236 5080 4264
rect 4387 4233 4399 4236
rect 4341 4227 4399 4233
rect 5074 4224 5080 4236
rect 5132 4224 5138 4276
rect 3605 4131 3663 4137
rect 3605 4097 3617 4131
rect 3651 4128 3663 4131
rect 5442 4128 5448 4140
rect 3651 4100 5448 4128
rect 3651 4097 3663 4100
rect 3605 4091 3663 4097
rect 5442 4088 5448 4100
rect 5500 4088 5506 4140
rect 2406 4020 2412 4072
rect 2464 4060 2470 4072
rect 3142 4060 3148 4072
rect 2464 4032 3148 4060
rect 2464 4020 2470 4032
rect 3142 4020 3148 4032
rect 3200 4060 3206 4072
rect 3329 4063 3387 4069
rect 3329 4060 3341 4063
rect 3200 4032 3341 4060
rect 3200 4020 3206 4032
rect 3329 4029 3341 4032
rect 3375 4029 3387 4063
rect 3329 4023 3387 4029
rect 1104 3834 4876 3856
rect 1104 3782 1421 3834
rect 1473 3782 1485 3834
rect 1537 3782 1549 3834
rect 1601 3782 1613 3834
rect 1665 3782 1677 3834
rect 1729 3782 2364 3834
rect 2416 3782 2428 3834
rect 2480 3782 2492 3834
rect 2544 3782 2556 3834
rect 2608 3782 2620 3834
rect 2672 3782 3307 3834
rect 3359 3782 3371 3834
rect 3423 3782 3435 3834
rect 3487 3782 3499 3834
rect 3551 3782 3563 3834
rect 3615 3782 4250 3834
rect 4302 3782 4314 3834
rect 4366 3782 4378 3834
rect 4430 3782 4442 3834
rect 4494 3782 4506 3834
rect 4558 3782 4876 3834
rect 1104 3760 4876 3782
rect 1104 3290 5035 3312
rect 1104 3238 1892 3290
rect 1944 3238 1956 3290
rect 2008 3238 2020 3290
rect 2072 3238 2084 3290
rect 2136 3238 2148 3290
rect 2200 3238 2835 3290
rect 2887 3238 2899 3290
rect 2951 3238 2963 3290
rect 3015 3238 3027 3290
rect 3079 3238 3091 3290
rect 3143 3238 3778 3290
rect 3830 3238 3842 3290
rect 3894 3238 3906 3290
rect 3958 3238 3970 3290
rect 4022 3238 4034 3290
rect 4086 3238 4721 3290
rect 4773 3238 4785 3290
rect 4837 3238 4849 3290
rect 4901 3238 4913 3290
rect 4965 3238 4977 3290
rect 5029 3238 5035 3290
rect 1104 3216 5035 3238
rect 3605 3043 3663 3049
rect 3605 3009 3617 3043
rect 3651 3040 3663 3043
rect 3694 3040 3700 3052
rect 3651 3012 3700 3040
rect 3651 3009 3663 3012
rect 3605 3003 3663 3009
rect 3694 3000 3700 3012
rect 3752 3000 3758 3052
rect 3142 2932 3148 2984
rect 3200 2972 3206 2984
rect 3329 2975 3387 2981
rect 3329 2972 3341 2975
rect 3200 2944 3341 2972
rect 3200 2932 3206 2944
rect 3329 2941 3341 2944
rect 3375 2941 3387 2975
rect 3329 2935 3387 2941
rect 4341 2839 4399 2845
rect 4341 2805 4353 2839
rect 4387 2836 4399 2839
rect 5074 2836 5080 2848
rect 4387 2808 5080 2836
rect 4387 2805 4399 2808
rect 4341 2799 4399 2805
rect 5074 2796 5080 2808
rect 5132 2796 5138 2848
rect 1104 2746 4876 2768
rect 1104 2694 1421 2746
rect 1473 2694 1485 2746
rect 1537 2694 1549 2746
rect 1601 2694 1613 2746
rect 1665 2694 1677 2746
rect 1729 2694 2364 2746
rect 2416 2694 2428 2746
rect 2480 2694 2492 2746
rect 2544 2694 2556 2746
rect 2608 2694 2620 2746
rect 2672 2694 3307 2746
rect 3359 2694 3371 2746
rect 3423 2694 3435 2746
rect 3487 2694 3499 2746
rect 3551 2694 3563 2746
rect 3615 2694 4250 2746
rect 4302 2694 4314 2746
rect 4366 2694 4378 2746
rect 4430 2694 4442 2746
rect 4494 2694 4506 2746
rect 4558 2694 4876 2746
rect 1104 2672 4876 2694
rect 1104 2202 5035 2224
rect 1104 2150 1892 2202
rect 1944 2150 1956 2202
rect 2008 2150 2020 2202
rect 2072 2150 2084 2202
rect 2136 2150 2148 2202
rect 2200 2150 2835 2202
rect 2887 2150 2899 2202
rect 2951 2150 2963 2202
rect 3015 2150 3027 2202
rect 3079 2150 3091 2202
rect 3143 2150 3778 2202
rect 3830 2150 3842 2202
rect 3894 2150 3906 2202
rect 3958 2150 3970 2202
rect 4022 2150 4034 2202
rect 4086 2150 4721 2202
rect 4773 2150 4785 2202
rect 4837 2150 4849 2202
rect 4901 2150 4913 2202
rect 4965 2150 4977 2202
rect 5029 2150 5035 2202
rect 1104 2128 5035 2150
rect 2501 2023 2559 2029
rect 2501 1989 2513 2023
rect 2547 2020 2559 2023
rect 4154 2020 4160 2032
rect 2547 1992 4160 2020
rect 2547 1989 2559 1992
rect 2501 1983 2559 1989
rect 4154 1980 4160 1992
rect 4212 2020 4218 2032
rect 5534 2020 5540 2032
rect 4212 1992 5540 2020
rect 4212 1980 4218 1992
rect 5534 1980 5540 1992
rect 5592 1980 5598 2032
rect 382 1912 388 1964
rect 440 1952 446 1964
rect 2041 1955 2099 1961
rect 2041 1952 2053 1955
rect 440 1924 2053 1952
rect 440 1912 446 1924
rect 2041 1921 2053 1924
rect 2087 1921 2099 1955
rect 2041 1915 2099 1921
rect 3697 1955 3755 1961
rect 3697 1921 3709 1955
rect 3743 1921 3755 1955
rect 3697 1915 3755 1921
rect 1762 1844 1768 1896
rect 1820 1884 1826 1896
rect 2222 1884 2228 1896
rect 1820 1856 2228 1884
rect 1820 1844 1826 1856
rect 2222 1844 2228 1856
rect 2280 1884 2286 1896
rect 3712 1884 3740 1915
rect 2280 1856 3740 1884
rect 3973 1887 4031 1893
rect 2280 1844 2286 1856
rect 3973 1853 3985 1887
rect 4019 1884 4031 1887
rect 4154 1884 4160 1896
rect 4019 1856 4160 1884
rect 4019 1853 4031 1856
rect 3973 1847 4031 1853
rect 4154 1844 4160 1856
rect 4212 1844 4218 1896
rect 1104 1658 4876 1680
rect 1104 1606 1421 1658
rect 1473 1606 1485 1658
rect 1537 1606 1549 1658
rect 1601 1606 1613 1658
rect 1665 1606 1677 1658
rect 1729 1606 2364 1658
rect 2416 1606 2428 1658
rect 2480 1606 2492 1658
rect 2544 1606 2556 1658
rect 2608 1606 2620 1658
rect 2672 1606 3307 1658
rect 3359 1606 3371 1658
rect 3423 1606 3435 1658
rect 3487 1606 3499 1658
rect 3551 1606 3563 1658
rect 3615 1606 4250 1658
rect 4302 1606 4314 1658
rect 4366 1606 4378 1658
rect 4430 1606 4442 1658
rect 4494 1606 4506 1658
rect 4558 1606 4876 1658
rect 1104 1584 4876 1606
rect 2590 1300 2596 1352
rect 2648 1340 2654 1352
rect 2961 1343 3019 1349
rect 2961 1340 2973 1343
rect 2648 1312 2973 1340
rect 2648 1300 2654 1312
rect 2961 1309 2973 1312
rect 3007 1340 3019 1343
rect 3142 1340 3148 1352
rect 3007 1312 3148 1340
rect 3007 1309 3019 1312
rect 2961 1303 3019 1309
rect 3142 1300 3148 1312
rect 3200 1300 3206 1352
rect 3237 1275 3295 1281
rect 3237 1241 3249 1275
rect 3283 1272 3295 1275
rect 3326 1272 3332 1284
rect 3283 1244 3332 1272
rect 3283 1241 3295 1244
rect 3237 1235 3295 1241
rect 3326 1232 3332 1244
rect 3384 1232 3390 1284
rect 1104 1114 5035 1136
rect 1104 1062 1892 1114
rect 1944 1062 1956 1114
rect 2008 1062 2020 1114
rect 2072 1062 2084 1114
rect 2136 1062 2148 1114
rect 2200 1062 2835 1114
rect 2887 1062 2899 1114
rect 2951 1062 2963 1114
rect 3015 1062 3027 1114
rect 3079 1062 3091 1114
rect 3143 1062 3778 1114
rect 3830 1062 3842 1114
rect 3894 1062 3906 1114
rect 3958 1062 3970 1114
rect 4022 1062 4034 1114
rect 4086 1062 4721 1114
rect 4773 1062 4785 1114
rect 4837 1062 4849 1114
rect 4901 1062 4913 1114
rect 4965 1062 4977 1114
rect 5029 1062 5035 1114
rect 1104 1040 5035 1062
<< via1 >>
rect 1892 22822 1944 22874
rect 1956 22822 2008 22874
rect 2020 22822 2072 22874
rect 2084 22822 2136 22874
rect 2148 22822 2200 22874
rect 2835 22822 2887 22874
rect 2899 22822 2951 22874
rect 2963 22822 3015 22874
rect 3027 22822 3079 22874
rect 3091 22822 3143 22874
rect 3778 22822 3830 22874
rect 3842 22822 3894 22874
rect 3906 22822 3958 22874
rect 3970 22822 4022 22874
rect 4034 22822 4086 22874
rect 4721 22822 4773 22874
rect 4785 22822 4837 22874
rect 4849 22822 4901 22874
rect 4913 22822 4965 22874
rect 4977 22822 5029 22874
rect 1421 22278 1473 22330
rect 1485 22278 1537 22330
rect 1549 22278 1601 22330
rect 1613 22278 1665 22330
rect 1677 22278 1729 22330
rect 2364 22278 2416 22330
rect 2428 22278 2480 22330
rect 2492 22278 2544 22330
rect 2556 22278 2608 22330
rect 2620 22278 2672 22330
rect 3307 22278 3359 22330
rect 3371 22278 3423 22330
rect 3435 22278 3487 22330
rect 3499 22278 3551 22330
rect 3563 22278 3615 22330
rect 4250 22278 4302 22330
rect 4314 22278 4366 22330
rect 4378 22278 4430 22330
rect 4442 22278 4494 22330
rect 4506 22278 4558 22330
rect 1892 21734 1944 21786
rect 1956 21734 2008 21786
rect 2020 21734 2072 21786
rect 2084 21734 2136 21786
rect 2148 21734 2200 21786
rect 2835 21734 2887 21786
rect 2899 21734 2951 21786
rect 2963 21734 3015 21786
rect 3027 21734 3079 21786
rect 3091 21734 3143 21786
rect 3778 21734 3830 21786
rect 3842 21734 3894 21786
rect 3906 21734 3958 21786
rect 3970 21734 4022 21786
rect 4034 21734 4086 21786
rect 4721 21734 4773 21786
rect 4785 21734 4837 21786
rect 4849 21734 4901 21786
rect 4913 21734 4965 21786
rect 4977 21734 5029 21786
rect 1421 21190 1473 21242
rect 1485 21190 1537 21242
rect 1549 21190 1601 21242
rect 1613 21190 1665 21242
rect 1677 21190 1729 21242
rect 2364 21190 2416 21242
rect 2428 21190 2480 21242
rect 2492 21190 2544 21242
rect 2556 21190 2608 21242
rect 2620 21190 2672 21242
rect 3307 21190 3359 21242
rect 3371 21190 3423 21242
rect 3435 21190 3487 21242
rect 3499 21190 3551 21242
rect 3563 21190 3615 21242
rect 4250 21190 4302 21242
rect 4314 21190 4366 21242
rect 4378 21190 4430 21242
rect 4442 21190 4494 21242
rect 4506 21190 4558 21242
rect 1892 20646 1944 20698
rect 1956 20646 2008 20698
rect 2020 20646 2072 20698
rect 2084 20646 2136 20698
rect 2148 20646 2200 20698
rect 2835 20646 2887 20698
rect 2899 20646 2951 20698
rect 2963 20646 3015 20698
rect 3027 20646 3079 20698
rect 3091 20646 3143 20698
rect 3778 20646 3830 20698
rect 3842 20646 3894 20698
rect 3906 20646 3958 20698
rect 3970 20646 4022 20698
rect 4034 20646 4086 20698
rect 4721 20646 4773 20698
rect 4785 20646 4837 20698
rect 4849 20646 4901 20698
rect 4913 20646 4965 20698
rect 4977 20646 5029 20698
rect 1421 20102 1473 20154
rect 1485 20102 1537 20154
rect 1549 20102 1601 20154
rect 1613 20102 1665 20154
rect 1677 20102 1729 20154
rect 2364 20102 2416 20154
rect 2428 20102 2480 20154
rect 2492 20102 2544 20154
rect 2556 20102 2608 20154
rect 2620 20102 2672 20154
rect 3307 20102 3359 20154
rect 3371 20102 3423 20154
rect 3435 20102 3487 20154
rect 3499 20102 3551 20154
rect 3563 20102 3615 20154
rect 4250 20102 4302 20154
rect 4314 20102 4366 20154
rect 4378 20102 4430 20154
rect 4442 20102 4494 20154
rect 4506 20102 4558 20154
rect 1892 19558 1944 19610
rect 1956 19558 2008 19610
rect 2020 19558 2072 19610
rect 2084 19558 2136 19610
rect 2148 19558 2200 19610
rect 2835 19558 2887 19610
rect 2899 19558 2951 19610
rect 2963 19558 3015 19610
rect 3027 19558 3079 19610
rect 3091 19558 3143 19610
rect 3778 19558 3830 19610
rect 3842 19558 3894 19610
rect 3906 19558 3958 19610
rect 3970 19558 4022 19610
rect 4034 19558 4086 19610
rect 4721 19558 4773 19610
rect 4785 19558 4837 19610
rect 4849 19558 4901 19610
rect 4913 19558 4965 19610
rect 4977 19558 5029 19610
rect 1421 19014 1473 19066
rect 1485 19014 1537 19066
rect 1549 19014 1601 19066
rect 1613 19014 1665 19066
rect 1677 19014 1729 19066
rect 2364 19014 2416 19066
rect 2428 19014 2480 19066
rect 2492 19014 2544 19066
rect 2556 19014 2608 19066
rect 2620 19014 2672 19066
rect 3307 19014 3359 19066
rect 3371 19014 3423 19066
rect 3435 19014 3487 19066
rect 3499 19014 3551 19066
rect 3563 19014 3615 19066
rect 4250 19014 4302 19066
rect 4314 19014 4366 19066
rect 4378 19014 4430 19066
rect 4442 19014 4494 19066
rect 4506 19014 4558 19066
rect 1892 18470 1944 18522
rect 1956 18470 2008 18522
rect 2020 18470 2072 18522
rect 2084 18470 2136 18522
rect 2148 18470 2200 18522
rect 2835 18470 2887 18522
rect 2899 18470 2951 18522
rect 2963 18470 3015 18522
rect 3027 18470 3079 18522
rect 3091 18470 3143 18522
rect 3778 18470 3830 18522
rect 3842 18470 3894 18522
rect 3906 18470 3958 18522
rect 3970 18470 4022 18522
rect 4034 18470 4086 18522
rect 4721 18470 4773 18522
rect 4785 18470 4837 18522
rect 4849 18470 4901 18522
rect 4913 18470 4965 18522
rect 4977 18470 5029 18522
rect 1421 17926 1473 17978
rect 1485 17926 1537 17978
rect 1549 17926 1601 17978
rect 1613 17926 1665 17978
rect 1677 17926 1729 17978
rect 2364 17926 2416 17978
rect 2428 17926 2480 17978
rect 2492 17926 2544 17978
rect 2556 17926 2608 17978
rect 2620 17926 2672 17978
rect 3307 17926 3359 17978
rect 3371 17926 3423 17978
rect 3435 17926 3487 17978
rect 3499 17926 3551 17978
rect 3563 17926 3615 17978
rect 4250 17926 4302 17978
rect 4314 17926 4366 17978
rect 4378 17926 4430 17978
rect 4442 17926 4494 17978
rect 4506 17926 4558 17978
rect 1892 17382 1944 17434
rect 1956 17382 2008 17434
rect 2020 17382 2072 17434
rect 2084 17382 2136 17434
rect 2148 17382 2200 17434
rect 2835 17382 2887 17434
rect 2899 17382 2951 17434
rect 2963 17382 3015 17434
rect 3027 17382 3079 17434
rect 3091 17382 3143 17434
rect 3778 17382 3830 17434
rect 3842 17382 3894 17434
rect 3906 17382 3958 17434
rect 3970 17382 4022 17434
rect 4034 17382 4086 17434
rect 4721 17382 4773 17434
rect 4785 17382 4837 17434
rect 4849 17382 4901 17434
rect 4913 17382 4965 17434
rect 4977 17382 5029 17434
rect 1421 16838 1473 16890
rect 1485 16838 1537 16890
rect 1549 16838 1601 16890
rect 1613 16838 1665 16890
rect 1677 16838 1729 16890
rect 2364 16838 2416 16890
rect 2428 16838 2480 16890
rect 2492 16838 2544 16890
rect 2556 16838 2608 16890
rect 2620 16838 2672 16890
rect 3307 16838 3359 16890
rect 3371 16838 3423 16890
rect 3435 16838 3487 16890
rect 3499 16838 3551 16890
rect 3563 16838 3615 16890
rect 4250 16838 4302 16890
rect 4314 16838 4366 16890
rect 4378 16838 4430 16890
rect 4442 16838 4494 16890
rect 4506 16838 4558 16890
rect 1892 16294 1944 16346
rect 1956 16294 2008 16346
rect 2020 16294 2072 16346
rect 2084 16294 2136 16346
rect 2148 16294 2200 16346
rect 2835 16294 2887 16346
rect 2899 16294 2951 16346
rect 2963 16294 3015 16346
rect 3027 16294 3079 16346
rect 3091 16294 3143 16346
rect 3778 16294 3830 16346
rect 3842 16294 3894 16346
rect 3906 16294 3958 16346
rect 3970 16294 4022 16346
rect 4034 16294 4086 16346
rect 4721 16294 4773 16346
rect 4785 16294 4837 16346
rect 4849 16294 4901 16346
rect 4913 16294 4965 16346
rect 4977 16294 5029 16346
rect 1421 15750 1473 15802
rect 1485 15750 1537 15802
rect 1549 15750 1601 15802
rect 1613 15750 1665 15802
rect 1677 15750 1729 15802
rect 2364 15750 2416 15802
rect 2428 15750 2480 15802
rect 2492 15750 2544 15802
rect 2556 15750 2608 15802
rect 2620 15750 2672 15802
rect 3307 15750 3359 15802
rect 3371 15750 3423 15802
rect 3435 15750 3487 15802
rect 3499 15750 3551 15802
rect 3563 15750 3615 15802
rect 4250 15750 4302 15802
rect 4314 15750 4366 15802
rect 4378 15750 4430 15802
rect 4442 15750 4494 15802
rect 4506 15750 4558 15802
rect 1892 15206 1944 15258
rect 1956 15206 2008 15258
rect 2020 15206 2072 15258
rect 2084 15206 2136 15258
rect 2148 15206 2200 15258
rect 2835 15206 2887 15258
rect 2899 15206 2951 15258
rect 2963 15206 3015 15258
rect 3027 15206 3079 15258
rect 3091 15206 3143 15258
rect 3778 15206 3830 15258
rect 3842 15206 3894 15258
rect 3906 15206 3958 15258
rect 3970 15206 4022 15258
rect 4034 15206 4086 15258
rect 4721 15206 4773 15258
rect 4785 15206 4837 15258
rect 4849 15206 4901 15258
rect 4913 15206 4965 15258
rect 4977 15206 5029 15258
rect 1421 14662 1473 14714
rect 1485 14662 1537 14714
rect 1549 14662 1601 14714
rect 1613 14662 1665 14714
rect 1677 14662 1729 14714
rect 2364 14662 2416 14714
rect 2428 14662 2480 14714
rect 2492 14662 2544 14714
rect 2556 14662 2608 14714
rect 2620 14662 2672 14714
rect 3307 14662 3359 14714
rect 3371 14662 3423 14714
rect 3435 14662 3487 14714
rect 3499 14662 3551 14714
rect 3563 14662 3615 14714
rect 4250 14662 4302 14714
rect 4314 14662 4366 14714
rect 4378 14662 4430 14714
rect 4442 14662 4494 14714
rect 4506 14662 4558 14714
rect 1892 14118 1944 14170
rect 1956 14118 2008 14170
rect 2020 14118 2072 14170
rect 2084 14118 2136 14170
rect 2148 14118 2200 14170
rect 2835 14118 2887 14170
rect 2899 14118 2951 14170
rect 2963 14118 3015 14170
rect 3027 14118 3079 14170
rect 3091 14118 3143 14170
rect 3778 14118 3830 14170
rect 3842 14118 3894 14170
rect 3906 14118 3958 14170
rect 3970 14118 4022 14170
rect 4034 14118 4086 14170
rect 4721 14118 4773 14170
rect 4785 14118 4837 14170
rect 4849 14118 4901 14170
rect 4913 14118 4965 14170
rect 4977 14118 5029 14170
rect 1421 13574 1473 13626
rect 1485 13574 1537 13626
rect 1549 13574 1601 13626
rect 1613 13574 1665 13626
rect 1677 13574 1729 13626
rect 2364 13574 2416 13626
rect 2428 13574 2480 13626
rect 2492 13574 2544 13626
rect 2556 13574 2608 13626
rect 2620 13574 2672 13626
rect 3307 13574 3359 13626
rect 3371 13574 3423 13626
rect 3435 13574 3487 13626
rect 3499 13574 3551 13626
rect 3563 13574 3615 13626
rect 4250 13574 4302 13626
rect 4314 13574 4366 13626
rect 4378 13574 4430 13626
rect 4442 13574 4494 13626
rect 4506 13574 4558 13626
rect 1892 13030 1944 13082
rect 1956 13030 2008 13082
rect 2020 13030 2072 13082
rect 2084 13030 2136 13082
rect 2148 13030 2200 13082
rect 2835 13030 2887 13082
rect 2899 13030 2951 13082
rect 2963 13030 3015 13082
rect 3027 13030 3079 13082
rect 3091 13030 3143 13082
rect 3778 13030 3830 13082
rect 3842 13030 3894 13082
rect 3906 13030 3958 13082
rect 3970 13030 4022 13082
rect 4034 13030 4086 13082
rect 4721 13030 4773 13082
rect 4785 13030 4837 13082
rect 4849 13030 4901 13082
rect 4913 13030 4965 13082
rect 4977 13030 5029 13082
rect 1421 12486 1473 12538
rect 1485 12486 1537 12538
rect 1549 12486 1601 12538
rect 1613 12486 1665 12538
rect 1677 12486 1729 12538
rect 2364 12486 2416 12538
rect 2428 12486 2480 12538
rect 2492 12486 2544 12538
rect 2556 12486 2608 12538
rect 2620 12486 2672 12538
rect 3307 12486 3359 12538
rect 3371 12486 3423 12538
rect 3435 12486 3487 12538
rect 3499 12486 3551 12538
rect 3563 12486 3615 12538
rect 4250 12486 4302 12538
rect 4314 12486 4366 12538
rect 4378 12486 4430 12538
rect 4442 12486 4494 12538
rect 4506 12486 4558 12538
rect 1892 11942 1944 11994
rect 1956 11942 2008 11994
rect 2020 11942 2072 11994
rect 2084 11942 2136 11994
rect 2148 11942 2200 11994
rect 2835 11942 2887 11994
rect 2899 11942 2951 11994
rect 2963 11942 3015 11994
rect 3027 11942 3079 11994
rect 3091 11942 3143 11994
rect 3778 11942 3830 11994
rect 3842 11942 3894 11994
rect 3906 11942 3958 11994
rect 3970 11942 4022 11994
rect 4034 11942 4086 11994
rect 4721 11942 4773 11994
rect 4785 11942 4837 11994
rect 4849 11942 4901 11994
rect 4913 11942 4965 11994
rect 4977 11942 5029 11994
rect 3148 11840 3200 11892
rect 5080 11704 5132 11756
rect 3884 11679 3936 11688
rect 3884 11645 3890 11679
rect 3890 11645 3924 11679
rect 3924 11645 3936 11679
rect 3884 11636 3936 11645
rect 4160 11636 4212 11688
rect 1768 11500 1820 11552
rect 3884 11500 3936 11552
rect 5080 11500 5132 11552
rect 1421 11398 1473 11450
rect 1485 11398 1537 11450
rect 1549 11398 1601 11450
rect 1613 11398 1665 11450
rect 1677 11398 1729 11450
rect 2364 11398 2416 11450
rect 2428 11398 2480 11450
rect 2492 11398 2544 11450
rect 2556 11398 2608 11450
rect 2620 11398 2672 11450
rect 3307 11398 3359 11450
rect 3371 11398 3423 11450
rect 3435 11398 3487 11450
rect 3499 11398 3551 11450
rect 3563 11398 3615 11450
rect 4250 11398 4302 11450
rect 4314 11398 4366 11450
rect 4378 11398 4430 11450
rect 4442 11398 4494 11450
rect 4506 11398 4558 11450
rect 3424 11271 3476 11280
rect 3424 11237 3433 11271
rect 3433 11237 3467 11271
rect 3467 11237 3476 11271
rect 3424 11228 3476 11237
rect 1216 11092 1268 11144
rect 2688 11135 2740 11144
rect 2688 11101 2697 11135
rect 2697 11101 2731 11135
rect 2731 11101 2740 11135
rect 2688 11092 2740 11101
rect 1892 10854 1944 10906
rect 1956 10854 2008 10906
rect 2020 10854 2072 10906
rect 2084 10854 2136 10906
rect 2148 10854 2200 10906
rect 2835 10854 2887 10906
rect 2899 10854 2951 10906
rect 2963 10854 3015 10906
rect 3027 10854 3079 10906
rect 3091 10854 3143 10906
rect 3778 10854 3830 10906
rect 3842 10854 3894 10906
rect 3906 10854 3958 10906
rect 3970 10854 4022 10906
rect 4034 10854 4086 10906
rect 4721 10854 4773 10906
rect 4785 10854 4837 10906
rect 4849 10854 4901 10906
rect 4913 10854 4965 10906
rect 4977 10854 5029 10906
rect 2228 10752 2280 10804
rect 3240 10752 3292 10804
rect 5172 10616 5224 10668
rect 3884 10591 3936 10600
rect 3884 10557 3890 10591
rect 3890 10557 3924 10591
rect 3924 10557 3936 10591
rect 3884 10548 3936 10557
rect 4160 10548 4212 10600
rect 3148 10412 3200 10464
rect 1421 10310 1473 10362
rect 1485 10310 1537 10362
rect 1549 10310 1601 10362
rect 1613 10310 1665 10362
rect 1677 10310 1729 10362
rect 2364 10310 2416 10362
rect 2428 10310 2480 10362
rect 2492 10310 2544 10362
rect 2556 10310 2608 10362
rect 2620 10310 2672 10362
rect 3307 10310 3359 10362
rect 3371 10310 3423 10362
rect 3435 10310 3487 10362
rect 3499 10310 3551 10362
rect 3563 10310 3615 10362
rect 4250 10310 4302 10362
rect 4314 10310 4366 10362
rect 4378 10310 4430 10362
rect 4442 10310 4494 10362
rect 4506 10310 4558 10362
rect 1308 10072 1360 10124
rect 5540 10072 5592 10124
rect 1124 10004 1176 10056
rect 3608 9936 3660 9988
rect 5264 9936 5316 9988
rect 2228 9868 2280 9920
rect 3884 9868 3936 9920
rect 4620 9868 4672 9920
rect 1892 9766 1944 9818
rect 1956 9766 2008 9818
rect 2020 9766 2072 9818
rect 2084 9766 2136 9818
rect 2148 9766 2200 9818
rect 2835 9766 2887 9818
rect 2899 9766 2951 9818
rect 2963 9766 3015 9818
rect 3027 9766 3079 9818
rect 3091 9766 3143 9818
rect 3778 9766 3830 9818
rect 3842 9766 3894 9818
rect 3906 9766 3958 9818
rect 3970 9766 4022 9818
rect 4034 9766 4086 9818
rect 4721 9766 4773 9818
rect 4785 9766 4837 9818
rect 4849 9766 4901 9818
rect 4913 9766 4965 9818
rect 4977 9766 5029 9818
rect 3884 9707 3936 9716
rect 3884 9673 3886 9707
rect 3886 9673 3920 9707
rect 3920 9673 3936 9707
rect 3884 9664 3936 9673
rect 3240 9528 3292 9580
rect 3608 9503 3660 9512
rect 3608 9469 3617 9503
rect 3617 9469 3651 9503
rect 3651 9469 3660 9503
rect 3608 9460 3660 9469
rect 4160 9460 4212 9512
rect 2688 9324 2740 9376
rect 3792 9324 3844 9376
rect 4528 9324 4580 9376
rect 1421 9222 1473 9274
rect 1485 9222 1537 9274
rect 1549 9222 1601 9274
rect 1613 9222 1665 9274
rect 1677 9222 1729 9274
rect 2364 9222 2416 9274
rect 2428 9222 2480 9274
rect 2492 9222 2544 9274
rect 2556 9222 2608 9274
rect 2620 9222 2672 9274
rect 3307 9222 3359 9274
rect 3371 9222 3423 9274
rect 3435 9222 3487 9274
rect 3499 9222 3551 9274
rect 3563 9222 3615 9274
rect 4250 9222 4302 9274
rect 4314 9222 4366 9274
rect 4378 9222 4430 9274
rect 4442 9222 4494 9274
rect 4506 9222 4558 9274
rect 1768 9120 1820 9172
rect 3516 9120 3568 9172
rect 3608 9120 3660 9172
rect 3884 9120 3936 9172
rect 2044 9027 2096 9036
rect 2044 8993 2056 9027
rect 2056 8993 2090 9027
rect 2090 8993 2096 9027
rect 2044 8984 2096 8993
rect 3700 8984 3752 9036
rect 1124 8916 1176 8968
rect 1676 8780 1728 8832
rect 5080 8780 5132 8832
rect 5264 8780 5316 8832
rect 1892 8678 1944 8730
rect 1956 8678 2008 8730
rect 2020 8678 2072 8730
rect 2084 8678 2136 8730
rect 2148 8678 2200 8730
rect 2835 8678 2887 8730
rect 2899 8678 2951 8730
rect 2963 8678 3015 8730
rect 3027 8678 3079 8730
rect 3091 8678 3143 8730
rect 3778 8678 3830 8730
rect 3842 8678 3894 8730
rect 3906 8678 3958 8730
rect 3970 8678 4022 8730
rect 4034 8678 4086 8730
rect 4721 8678 4773 8730
rect 4785 8678 4837 8730
rect 4849 8678 4901 8730
rect 4913 8678 4965 8730
rect 4977 8678 5029 8730
rect 1676 8576 1728 8628
rect 2136 8576 2188 8628
rect 3608 8576 3660 8628
rect 3700 8440 3752 8492
rect 3516 8372 3568 8424
rect 5540 8440 5592 8492
rect 4160 8372 4212 8424
rect 1308 8236 1360 8288
rect 1421 8134 1473 8186
rect 1485 8134 1537 8186
rect 1549 8134 1601 8186
rect 1613 8134 1665 8186
rect 1677 8134 1729 8186
rect 2364 8134 2416 8186
rect 2428 8134 2480 8186
rect 2492 8134 2544 8186
rect 2556 8134 2608 8186
rect 2620 8134 2672 8186
rect 3307 8134 3359 8186
rect 3371 8134 3423 8186
rect 3435 8134 3487 8186
rect 3499 8134 3551 8186
rect 3563 8134 3615 8186
rect 4250 8134 4302 8186
rect 4314 8134 4366 8186
rect 4378 8134 4430 8186
rect 4442 8134 4494 8186
rect 4506 8134 4558 8186
rect 1860 7896 1912 7948
rect 5448 7896 5500 7948
rect 1124 7828 1176 7880
rect 1584 7871 1636 7880
rect 1584 7837 1593 7871
rect 1593 7837 1627 7871
rect 1627 7837 1636 7871
rect 1584 7828 1636 7837
rect 1124 7692 1176 7744
rect 1860 7692 1912 7744
rect 2044 7735 2096 7744
rect 2044 7701 2059 7735
rect 2059 7701 2093 7735
rect 2093 7701 2096 7735
rect 2044 7692 2096 7701
rect 3700 7692 3752 7744
rect 1892 7590 1944 7642
rect 1956 7590 2008 7642
rect 2020 7590 2072 7642
rect 2084 7590 2136 7642
rect 2148 7590 2200 7642
rect 2835 7590 2887 7642
rect 2899 7590 2951 7642
rect 2963 7590 3015 7642
rect 3027 7590 3079 7642
rect 3091 7590 3143 7642
rect 3778 7590 3830 7642
rect 3842 7590 3894 7642
rect 3906 7590 3958 7642
rect 3970 7590 4022 7642
rect 4034 7590 4086 7642
rect 4721 7590 4773 7642
rect 4785 7590 4837 7642
rect 4849 7590 4901 7642
rect 4913 7590 4965 7642
rect 4977 7590 5029 7642
rect 1768 7488 1820 7540
rect 1584 7420 1636 7472
rect 2228 7420 2280 7472
rect 2320 7420 2372 7472
rect 2780 7420 2832 7472
rect 5356 7352 5408 7404
rect 3700 7284 3752 7336
rect 4160 7284 4212 7336
rect 1421 7046 1473 7098
rect 1485 7046 1537 7098
rect 1549 7046 1601 7098
rect 1613 7046 1665 7098
rect 1677 7046 1729 7098
rect 2364 7046 2416 7098
rect 2428 7046 2480 7098
rect 2492 7046 2544 7098
rect 2556 7046 2608 7098
rect 2620 7046 2672 7098
rect 3307 7046 3359 7098
rect 3371 7046 3423 7098
rect 3435 7046 3487 7098
rect 3499 7046 3551 7098
rect 3563 7046 3615 7098
rect 4250 7046 4302 7098
rect 4314 7046 4366 7098
rect 4378 7046 4430 7098
rect 4442 7046 4494 7098
rect 4506 7046 4558 7098
rect 5172 6944 5224 6996
rect 1216 6808 1268 6860
rect 3148 6740 3200 6792
rect 2596 6672 2648 6724
rect 2780 6672 2832 6724
rect 3700 6604 3752 6656
rect 1892 6502 1944 6554
rect 1956 6502 2008 6554
rect 2020 6502 2072 6554
rect 2084 6502 2136 6554
rect 2148 6502 2200 6554
rect 2835 6502 2887 6554
rect 2899 6502 2951 6554
rect 2963 6502 3015 6554
rect 3027 6502 3079 6554
rect 3091 6502 3143 6554
rect 3778 6502 3830 6554
rect 3842 6502 3894 6554
rect 3906 6502 3958 6554
rect 3970 6502 4022 6554
rect 4034 6502 4086 6554
rect 4721 6502 4773 6554
rect 4785 6502 4837 6554
rect 4849 6502 4901 6554
rect 4913 6502 4965 6554
rect 4977 6502 5029 6554
rect 2688 6332 2740 6384
rect 3700 6264 3752 6316
rect 2228 6196 2280 6248
rect 4160 6196 4212 6248
rect 4620 6196 4672 6248
rect 1768 6060 1820 6112
rect 2228 6060 2280 6112
rect 1421 5958 1473 6010
rect 1485 5958 1537 6010
rect 1549 5958 1601 6010
rect 1613 5958 1665 6010
rect 1677 5958 1729 6010
rect 2364 5958 2416 6010
rect 2428 5958 2480 6010
rect 2492 5958 2544 6010
rect 2556 5958 2608 6010
rect 2620 5958 2672 6010
rect 3307 5958 3359 6010
rect 3371 5958 3423 6010
rect 3435 5958 3487 6010
rect 3499 5958 3551 6010
rect 3563 5958 3615 6010
rect 4250 5958 4302 6010
rect 4314 5958 4366 6010
rect 4378 5958 4430 6010
rect 4442 5958 4494 6010
rect 4506 5958 4558 6010
rect 3700 5856 3752 5908
rect 3240 5788 3292 5840
rect 4712 5788 4764 5840
rect 1216 5720 1268 5772
rect 1768 5720 1820 5772
rect 1308 5584 1360 5636
rect 1892 5414 1944 5466
rect 1956 5414 2008 5466
rect 2020 5414 2072 5466
rect 2084 5414 2136 5466
rect 2148 5414 2200 5466
rect 2835 5414 2887 5466
rect 2899 5414 2951 5466
rect 2963 5414 3015 5466
rect 3027 5414 3079 5466
rect 3091 5414 3143 5466
rect 3778 5414 3830 5466
rect 3842 5414 3894 5466
rect 3906 5414 3958 5466
rect 3970 5414 4022 5466
rect 4034 5414 4086 5466
rect 4721 5414 4773 5466
rect 4785 5414 4837 5466
rect 4849 5414 4901 5466
rect 4913 5414 4965 5466
rect 4977 5414 5029 5466
rect 5172 5312 5224 5364
rect 2228 5176 2280 5228
rect 3240 5176 3292 5228
rect 1860 5151 1912 5160
rect 1860 5117 1869 5151
rect 1869 5117 1903 5151
rect 1903 5117 1912 5151
rect 1860 5108 1912 5117
rect 3148 5108 3200 5160
rect 2688 4972 2740 5024
rect 1421 4870 1473 4922
rect 1485 4870 1537 4922
rect 1549 4870 1601 4922
rect 1613 4870 1665 4922
rect 1677 4870 1729 4922
rect 2364 4870 2416 4922
rect 2428 4870 2480 4922
rect 2492 4870 2544 4922
rect 2556 4870 2608 4922
rect 2620 4870 2672 4922
rect 3307 4870 3359 4922
rect 3371 4870 3423 4922
rect 3435 4870 3487 4922
rect 3499 4870 3551 4922
rect 3563 4870 3615 4922
rect 4250 4870 4302 4922
rect 4314 4870 4366 4922
rect 4378 4870 4430 4922
rect 4442 4870 4494 4922
rect 4506 4870 4558 4922
rect 4160 4768 4212 4820
rect 1860 4564 1912 4616
rect 2412 4607 2464 4616
rect 2412 4573 2421 4607
rect 2421 4573 2455 4607
rect 2455 4573 2464 4607
rect 2412 4564 2464 4573
rect 5264 4632 5316 4684
rect 4160 4607 4212 4616
rect 4160 4573 4169 4607
rect 4169 4573 4203 4607
rect 4203 4573 4212 4607
rect 4160 4564 4212 4573
rect 5172 4428 5224 4480
rect 1892 4326 1944 4378
rect 1956 4326 2008 4378
rect 2020 4326 2072 4378
rect 2084 4326 2136 4378
rect 2148 4326 2200 4378
rect 2835 4326 2887 4378
rect 2899 4326 2951 4378
rect 2963 4326 3015 4378
rect 3027 4326 3079 4378
rect 3091 4326 3143 4378
rect 3778 4326 3830 4378
rect 3842 4326 3894 4378
rect 3906 4326 3958 4378
rect 3970 4326 4022 4378
rect 4034 4326 4086 4378
rect 4721 4326 4773 4378
rect 4785 4326 4837 4378
rect 4849 4326 4901 4378
rect 4913 4326 4965 4378
rect 4977 4326 5029 4378
rect 5080 4224 5132 4276
rect 5448 4088 5500 4140
rect 2412 4020 2464 4072
rect 3148 4020 3200 4072
rect 1421 3782 1473 3834
rect 1485 3782 1537 3834
rect 1549 3782 1601 3834
rect 1613 3782 1665 3834
rect 1677 3782 1729 3834
rect 2364 3782 2416 3834
rect 2428 3782 2480 3834
rect 2492 3782 2544 3834
rect 2556 3782 2608 3834
rect 2620 3782 2672 3834
rect 3307 3782 3359 3834
rect 3371 3782 3423 3834
rect 3435 3782 3487 3834
rect 3499 3782 3551 3834
rect 3563 3782 3615 3834
rect 4250 3782 4302 3834
rect 4314 3782 4366 3834
rect 4378 3782 4430 3834
rect 4442 3782 4494 3834
rect 4506 3782 4558 3834
rect 1892 3238 1944 3290
rect 1956 3238 2008 3290
rect 2020 3238 2072 3290
rect 2084 3238 2136 3290
rect 2148 3238 2200 3290
rect 2835 3238 2887 3290
rect 2899 3238 2951 3290
rect 2963 3238 3015 3290
rect 3027 3238 3079 3290
rect 3091 3238 3143 3290
rect 3778 3238 3830 3290
rect 3842 3238 3894 3290
rect 3906 3238 3958 3290
rect 3970 3238 4022 3290
rect 4034 3238 4086 3290
rect 4721 3238 4773 3290
rect 4785 3238 4837 3290
rect 4849 3238 4901 3290
rect 4913 3238 4965 3290
rect 4977 3238 5029 3290
rect 3700 3000 3752 3052
rect 3148 2932 3200 2984
rect 5080 2796 5132 2848
rect 1421 2694 1473 2746
rect 1485 2694 1537 2746
rect 1549 2694 1601 2746
rect 1613 2694 1665 2746
rect 1677 2694 1729 2746
rect 2364 2694 2416 2746
rect 2428 2694 2480 2746
rect 2492 2694 2544 2746
rect 2556 2694 2608 2746
rect 2620 2694 2672 2746
rect 3307 2694 3359 2746
rect 3371 2694 3423 2746
rect 3435 2694 3487 2746
rect 3499 2694 3551 2746
rect 3563 2694 3615 2746
rect 4250 2694 4302 2746
rect 4314 2694 4366 2746
rect 4378 2694 4430 2746
rect 4442 2694 4494 2746
rect 4506 2694 4558 2746
rect 1892 2150 1944 2202
rect 1956 2150 2008 2202
rect 2020 2150 2072 2202
rect 2084 2150 2136 2202
rect 2148 2150 2200 2202
rect 2835 2150 2887 2202
rect 2899 2150 2951 2202
rect 2963 2150 3015 2202
rect 3027 2150 3079 2202
rect 3091 2150 3143 2202
rect 3778 2150 3830 2202
rect 3842 2150 3894 2202
rect 3906 2150 3958 2202
rect 3970 2150 4022 2202
rect 4034 2150 4086 2202
rect 4721 2150 4773 2202
rect 4785 2150 4837 2202
rect 4849 2150 4901 2202
rect 4913 2150 4965 2202
rect 4977 2150 5029 2202
rect 4160 1980 4212 2032
rect 5540 1980 5592 2032
rect 388 1912 440 1964
rect 1768 1844 1820 1896
rect 2228 1844 2280 1896
rect 4160 1844 4212 1896
rect 1421 1606 1473 1658
rect 1485 1606 1537 1658
rect 1549 1606 1601 1658
rect 1613 1606 1665 1658
rect 1677 1606 1729 1658
rect 2364 1606 2416 1658
rect 2428 1606 2480 1658
rect 2492 1606 2544 1658
rect 2556 1606 2608 1658
rect 2620 1606 2672 1658
rect 3307 1606 3359 1658
rect 3371 1606 3423 1658
rect 3435 1606 3487 1658
rect 3499 1606 3551 1658
rect 3563 1606 3615 1658
rect 4250 1606 4302 1658
rect 4314 1606 4366 1658
rect 4378 1606 4430 1658
rect 4442 1606 4494 1658
rect 4506 1606 4558 1658
rect 2596 1300 2648 1352
rect 3148 1300 3200 1352
rect 3332 1232 3384 1284
rect 1892 1062 1944 1114
rect 1956 1062 2008 1114
rect 2020 1062 2072 1114
rect 2084 1062 2136 1114
rect 2148 1062 2200 1114
rect 2835 1062 2887 1114
rect 2899 1062 2951 1114
rect 2963 1062 3015 1114
rect 3027 1062 3079 1114
rect 3091 1062 3143 1114
rect 3778 1062 3830 1114
rect 3842 1062 3894 1114
rect 3906 1062 3958 1114
rect 3970 1062 4022 1114
rect 4034 1062 4086 1114
rect 4721 1062 4773 1114
rect 4785 1062 4837 1114
rect 4849 1062 4901 1114
rect 4913 1062 4965 1114
rect 4977 1062 5029 1114
<< metal2 >>
rect 5078 23216 5134 23225
rect 5134 23174 5304 23202
rect 5078 23151 5134 23160
rect 1892 22876 2200 22885
rect 1892 22874 1898 22876
rect 1954 22874 1978 22876
rect 2034 22874 2058 22876
rect 2114 22874 2138 22876
rect 2194 22874 2200 22876
rect 1954 22822 1956 22874
rect 2136 22822 2138 22874
rect 1892 22820 1898 22822
rect 1954 22820 1978 22822
rect 2034 22820 2058 22822
rect 2114 22820 2138 22822
rect 2194 22820 2200 22822
rect 1892 22811 2200 22820
rect 2835 22876 3143 22885
rect 2835 22874 2841 22876
rect 2897 22874 2921 22876
rect 2977 22874 3001 22876
rect 3057 22874 3081 22876
rect 3137 22874 3143 22876
rect 2897 22822 2899 22874
rect 3079 22822 3081 22874
rect 2835 22820 2841 22822
rect 2897 22820 2921 22822
rect 2977 22820 3001 22822
rect 3057 22820 3081 22822
rect 3137 22820 3143 22822
rect 2835 22811 3143 22820
rect 3778 22876 4086 22885
rect 3778 22874 3784 22876
rect 3840 22874 3864 22876
rect 3920 22874 3944 22876
rect 4000 22874 4024 22876
rect 4080 22874 4086 22876
rect 3840 22822 3842 22874
rect 4022 22822 4024 22874
rect 3778 22820 3784 22822
rect 3840 22820 3864 22822
rect 3920 22820 3944 22822
rect 4000 22820 4024 22822
rect 4080 22820 4086 22822
rect 3778 22811 4086 22820
rect 4721 22876 5029 22885
rect 4721 22874 4727 22876
rect 4783 22874 4807 22876
rect 4863 22874 4887 22876
rect 4943 22874 4967 22876
rect 5023 22874 5029 22876
rect 4783 22822 4785 22874
rect 4965 22822 4967 22874
rect 4721 22820 4727 22822
rect 4783 22820 4807 22822
rect 4863 22820 4887 22822
rect 4943 22820 4967 22822
rect 5023 22820 5029 22822
rect 4721 22811 5029 22820
rect 1421 22332 1729 22341
rect 1421 22330 1427 22332
rect 1483 22330 1507 22332
rect 1563 22330 1587 22332
rect 1643 22330 1667 22332
rect 1723 22330 1729 22332
rect 1483 22278 1485 22330
rect 1665 22278 1667 22330
rect 1421 22276 1427 22278
rect 1483 22276 1507 22278
rect 1563 22276 1587 22278
rect 1643 22276 1667 22278
rect 1723 22276 1729 22278
rect 1421 22267 1729 22276
rect 2364 22332 2672 22341
rect 2364 22330 2370 22332
rect 2426 22330 2450 22332
rect 2506 22330 2530 22332
rect 2586 22330 2610 22332
rect 2666 22330 2672 22332
rect 2426 22278 2428 22330
rect 2608 22278 2610 22330
rect 2364 22276 2370 22278
rect 2426 22276 2450 22278
rect 2506 22276 2530 22278
rect 2586 22276 2610 22278
rect 2666 22276 2672 22278
rect 2364 22267 2672 22276
rect 3307 22332 3615 22341
rect 3307 22330 3313 22332
rect 3369 22330 3393 22332
rect 3449 22330 3473 22332
rect 3529 22330 3553 22332
rect 3609 22330 3615 22332
rect 3369 22278 3371 22330
rect 3551 22278 3553 22330
rect 3307 22276 3313 22278
rect 3369 22276 3393 22278
rect 3449 22276 3473 22278
rect 3529 22276 3553 22278
rect 3609 22276 3615 22278
rect 3307 22267 3615 22276
rect 4250 22332 4558 22341
rect 4250 22330 4256 22332
rect 4312 22330 4336 22332
rect 4392 22330 4416 22332
rect 4472 22330 4496 22332
rect 4552 22330 4558 22332
rect 4312 22278 4314 22330
rect 4494 22278 4496 22330
rect 4250 22276 4256 22278
rect 4312 22276 4336 22278
rect 4392 22276 4416 22278
rect 4472 22276 4496 22278
rect 4552 22276 4558 22278
rect 4250 22267 4558 22276
rect 1892 21788 2200 21797
rect 1892 21786 1898 21788
rect 1954 21786 1978 21788
rect 2034 21786 2058 21788
rect 2114 21786 2138 21788
rect 2194 21786 2200 21788
rect 1954 21734 1956 21786
rect 2136 21734 2138 21786
rect 1892 21732 1898 21734
rect 1954 21732 1978 21734
rect 2034 21732 2058 21734
rect 2114 21732 2138 21734
rect 2194 21732 2200 21734
rect 1892 21723 2200 21732
rect 2835 21788 3143 21797
rect 2835 21786 2841 21788
rect 2897 21786 2921 21788
rect 2977 21786 3001 21788
rect 3057 21786 3081 21788
rect 3137 21786 3143 21788
rect 2897 21734 2899 21786
rect 3079 21734 3081 21786
rect 2835 21732 2841 21734
rect 2897 21732 2921 21734
rect 2977 21732 3001 21734
rect 3057 21732 3081 21734
rect 3137 21732 3143 21734
rect 2835 21723 3143 21732
rect 3778 21788 4086 21797
rect 3778 21786 3784 21788
rect 3840 21786 3864 21788
rect 3920 21786 3944 21788
rect 4000 21786 4024 21788
rect 4080 21786 4086 21788
rect 3840 21734 3842 21786
rect 4022 21734 4024 21786
rect 3778 21732 3784 21734
rect 3840 21732 3864 21734
rect 3920 21732 3944 21734
rect 4000 21732 4024 21734
rect 4080 21732 4086 21734
rect 3778 21723 4086 21732
rect 4721 21788 5029 21797
rect 4721 21786 4727 21788
rect 4783 21786 4807 21788
rect 4863 21786 4887 21788
rect 4943 21786 4967 21788
rect 5023 21786 5029 21788
rect 4783 21734 4785 21786
rect 4965 21734 4967 21786
rect 4721 21732 4727 21734
rect 4783 21732 4807 21734
rect 4863 21732 4887 21734
rect 4943 21732 4967 21734
rect 5023 21732 5029 21734
rect 4721 21723 5029 21732
rect 5170 21448 5226 21457
rect 5170 21383 5226 21392
rect 1421 21244 1729 21253
rect 1421 21242 1427 21244
rect 1483 21242 1507 21244
rect 1563 21242 1587 21244
rect 1643 21242 1667 21244
rect 1723 21242 1729 21244
rect 1483 21190 1485 21242
rect 1665 21190 1667 21242
rect 1421 21188 1427 21190
rect 1483 21188 1507 21190
rect 1563 21188 1587 21190
rect 1643 21188 1667 21190
rect 1723 21188 1729 21190
rect 1421 21179 1729 21188
rect 2364 21244 2672 21253
rect 2364 21242 2370 21244
rect 2426 21242 2450 21244
rect 2506 21242 2530 21244
rect 2586 21242 2610 21244
rect 2666 21242 2672 21244
rect 2426 21190 2428 21242
rect 2608 21190 2610 21242
rect 2364 21188 2370 21190
rect 2426 21188 2450 21190
rect 2506 21188 2530 21190
rect 2586 21188 2610 21190
rect 2666 21188 2672 21190
rect 2364 21179 2672 21188
rect 3307 21244 3615 21253
rect 3307 21242 3313 21244
rect 3369 21242 3393 21244
rect 3449 21242 3473 21244
rect 3529 21242 3553 21244
rect 3609 21242 3615 21244
rect 3369 21190 3371 21242
rect 3551 21190 3553 21242
rect 3307 21188 3313 21190
rect 3369 21188 3393 21190
rect 3449 21188 3473 21190
rect 3529 21188 3553 21190
rect 3609 21188 3615 21190
rect 3307 21179 3615 21188
rect 4250 21244 4558 21253
rect 4250 21242 4256 21244
rect 4312 21242 4336 21244
rect 4392 21242 4416 21244
rect 4472 21242 4496 21244
rect 4552 21242 4558 21244
rect 4312 21190 4314 21242
rect 4494 21190 4496 21242
rect 4250 21188 4256 21190
rect 4312 21188 4336 21190
rect 4392 21188 4416 21190
rect 4472 21188 4496 21190
rect 4552 21188 4558 21190
rect 4250 21179 4558 21188
rect 1892 20700 2200 20709
rect 1892 20698 1898 20700
rect 1954 20698 1978 20700
rect 2034 20698 2058 20700
rect 2114 20698 2138 20700
rect 2194 20698 2200 20700
rect 1954 20646 1956 20698
rect 2136 20646 2138 20698
rect 1892 20644 1898 20646
rect 1954 20644 1978 20646
rect 2034 20644 2058 20646
rect 2114 20644 2138 20646
rect 2194 20644 2200 20646
rect 1892 20635 2200 20644
rect 2835 20700 3143 20709
rect 2835 20698 2841 20700
rect 2897 20698 2921 20700
rect 2977 20698 3001 20700
rect 3057 20698 3081 20700
rect 3137 20698 3143 20700
rect 2897 20646 2899 20698
rect 3079 20646 3081 20698
rect 2835 20644 2841 20646
rect 2897 20644 2921 20646
rect 2977 20644 3001 20646
rect 3057 20644 3081 20646
rect 3137 20644 3143 20646
rect 2835 20635 3143 20644
rect 3778 20700 4086 20709
rect 3778 20698 3784 20700
rect 3840 20698 3864 20700
rect 3920 20698 3944 20700
rect 4000 20698 4024 20700
rect 4080 20698 4086 20700
rect 3840 20646 3842 20698
rect 4022 20646 4024 20698
rect 3778 20644 3784 20646
rect 3840 20644 3864 20646
rect 3920 20644 3944 20646
rect 4000 20644 4024 20646
rect 4080 20644 4086 20646
rect 3778 20635 4086 20644
rect 4721 20700 5029 20709
rect 4721 20698 4727 20700
rect 4783 20698 4807 20700
rect 4863 20698 4887 20700
rect 4943 20698 4967 20700
rect 5023 20698 5029 20700
rect 4783 20646 4785 20698
rect 4965 20646 4967 20698
rect 4721 20644 4727 20646
rect 4783 20644 4807 20646
rect 4863 20644 4887 20646
rect 4943 20644 4967 20646
rect 5023 20644 5029 20646
rect 4721 20635 5029 20644
rect 1421 20156 1729 20165
rect 1421 20154 1427 20156
rect 1483 20154 1507 20156
rect 1563 20154 1587 20156
rect 1643 20154 1667 20156
rect 1723 20154 1729 20156
rect 1483 20102 1485 20154
rect 1665 20102 1667 20154
rect 1421 20100 1427 20102
rect 1483 20100 1507 20102
rect 1563 20100 1587 20102
rect 1643 20100 1667 20102
rect 1723 20100 1729 20102
rect 1421 20091 1729 20100
rect 2364 20156 2672 20165
rect 2364 20154 2370 20156
rect 2426 20154 2450 20156
rect 2506 20154 2530 20156
rect 2586 20154 2610 20156
rect 2666 20154 2672 20156
rect 2426 20102 2428 20154
rect 2608 20102 2610 20154
rect 2364 20100 2370 20102
rect 2426 20100 2450 20102
rect 2506 20100 2530 20102
rect 2586 20100 2610 20102
rect 2666 20100 2672 20102
rect 2364 20091 2672 20100
rect 3307 20156 3615 20165
rect 3307 20154 3313 20156
rect 3369 20154 3393 20156
rect 3449 20154 3473 20156
rect 3529 20154 3553 20156
rect 3609 20154 3615 20156
rect 3369 20102 3371 20154
rect 3551 20102 3553 20154
rect 3307 20100 3313 20102
rect 3369 20100 3393 20102
rect 3449 20100 3473 20102
rect 3529 20100 3553 20102
rect 3609 20100 3615 20102
rect 3307 20091 3615 20100
rect 4250 20156 4558 20165
rect 4250 20154 4256 20156
rect 4312 20154 4336 20156
rect 4392 20154 4416 20156
rect 4472 20154 4496 20156
rect 4552 20154 4558 20156
rect 4312 20102 4314 20154
rect 4494 20102 4496 20154
rect 4250 20100 4256 20102
rect 4312 20100 4336 20102
rect 4392 20100 4416 20102
rect 4472 20100 4496 20102
rect 4552 20100 4558 20102
rect 4250 20091 4558 20100
rect 1892 19612 2200 19621
rect 1892 19610 1898 19612
rect 1954 19610 1978 19612
rect 2034 19610 2058 19612
rect 2114 19610 2138 19612
rect 2194 19610 2200 19612
rect 1954 19558 1956 19610
rect 2136 19558 2138 19610
rect 1892 19556 1898 19558
rect 1954 19556 1978 19558
rect 2034 19556 2058 19558
rect 2114 19556 2138 19558
rect 2194 19556 2200 19558
rect 1892 19547 2200 19556
rect 2835 19612 3143 19621
rect 2835 19610 2841 19612
rect 2897 19610 2921 19612
rect 2977 19610 3001 19612
rect 3057 19610 3081 19612
rect 3137 19610 3143 19612
rect 2897 19558 2899 19610
rect 3079 19558 3081 19610
rect 2835 19556 2841 19558
rect 2897 19556 2921 19558
rect 2977 19556 3001 19558
rect 3057 19556 3081 19558
rect 3137 19556 3143 19558
rect 2835 19547 3143 19556
rect 3778 19612 4086 19621
rect 3778 19610 3784 19612
rect 3840 19610 3864 19612
rect 3920 19610 3944 19612
rect 4000 19610 4024 19612
rect 4080 19610 4086 19612
rect 3840 19558 3842 19610
rect 4022 19558 4024 19610
rect 3778 19556 3784 19558
rect 3840 19556 3864 19558
rect 3920 19556 3944 19558
rect 4000 19556 4024 19558
rect 4080 19556 4086 19558
rect 3778 19547 4086 19556
rect 4721 19612 5029 19621
rect 4721 19610 4727 19612
rect 4783 19610 4807 19612
rect 4863 19610 4887 19612
rect 4943 19610 4967 19612
rect 5023 19610 5029 19612
rect 4783 19558 4785 19610
rect 4965 19558 4967 19610
rect 4721 19556 4727 19558
rect 4783 19556 4807 19558
rect 4863 19556 4887 19558
rect 4943 19556 4967 19558
rect 5023 19556 5029 19558
rect 4721 19547 5029 19556
rect 1421 19068 1729 19077
rect 1421 19066 1427 19068
rect 1483 19066 1507 19068
rect 1563 19066 1587 19068
rect 1643 19066 1667 19068
rect 1723 19066 1729 19068
rect 1483 19014 1485 19066
rect 1665 19014 1667 19066
rect 1421 19012 1427 19014
rect 1483 19012 1507 19014
rect 1563 19012 1587 19014
rect 1643 19012 1667 19014
rect 1723 19012 1729 19014
rect 1421 19003 1729 19012
rect 2364 19068 2672 19077
rect 2364 19066 2370 19068
rect 2426 19066 2450 19068
rect 2506 19066 2530 19068
rect 2586 19066 2610 19068
rect 2666 19066 2672 19068
rect 2426 19014 2428 19066
rect 2608 19014 2610 19066
rect 2364 19012 2370 19014
rect 2426 19012 2450 19014
rect 2506 19012 2530 19014
rect 2586 19012 2610 19014
rect 2666 19012 2672 19014
rect 2364 19003 2672 19012
rect 3307 19068 3615 19077
rect 3307 19066 3313 19068
rect 3369 19066 3393 19068
rect 3449 19066 3473 19068
rect 3529 19066 3553 19068
rect 3609 19066 3615 19068
rect 3369 19014 3371 19066
rect 3551 19014 3553 19066
rect 3307 19012 3313 19014
rect 3369 19012 3393 19014
rect 3449 19012 3473 19014
rect 3529 19012 3553 19014
rect 3609 19012 3615 19014
rect 3307 19003 3615 19012
rect 4250 19068 4558 19077
rect 4250 19066 4256 19068
rect 4312 19066 4336 19068
rect 4392 19066 4416 19068
rect 4472 19066 4496 19068
rect 4552 19066 4558 19068
rect 4312 19014 4314 19066
rect 4494 19014 4496 19066
rect 4250 19012 4256 19014
rect 4312 19012 4336 19014
rect 4392 19012 4416 19014
rect 4472 19012 4496 19014
rect 4552 19012 4558 19014
rect 4250 19003 4558 19012
rect 4618 18728 4674 18737
rect 4618 18663 4674 18672
rect 1892 18524 2200 18533
rect 1892 18522 1898 18524
rect 1954 18522 1978 18524
rect 2034 18522 2058 18524
rect 2114 18522 2138 18524
rect 2194 18522 2200 18524
rect 1954 18470 1956 18522
rect 2136 18470 2138 18522
rect 1892 18468 1898 18470
rect 1954 18468 1978 18470
rect 2034 18468 2058 18470
rect 2114 18468 2138 18470
rect 2194 18468 2200 18470
rect 1892 18459 2200 18468
rect 2835 18524 3143 18533
rect 2835 18522 2841 18524
rect 2897 18522 2921 18524
rect 2977 18522 3001 18524
rect 3057 18522 3081 18524
rect 3137 18522 3143 18524
rect 2897 18470 2899 18522
rect 3079 18470 3081 18522
rect 2835 18468 2841 18470
rect 2897 18468 2921 18470
rect 2977 18468 3001 18470
rect 3057 18468 3081 18470
rect 3137 18468 3143 18470
rect 2835 18459 3143 18468
rect 3778 18524 4086 18533
rect 3778 18522 3784 18524
rect 3840 18522 3864 18524
rect 3920 18522 3944 18524
rect 4000 18522 4024 18524
rect 4080 18522 4086 18524
rect 3840 18470 3842 18522
rect 4022 18470 4024 18522
rect 3778 18468 3784 18470
rect 3840 18468 3864 18470
rect 3920 18468 3944 18470
rect 4000 18468 4024 18470
rect 4080 18468 4086 18470
rect 3778 18459 4086 18468
rect 1421 17980 1729 17989
rect 1421 17978 1427 17980
rect 1483 17978 1507 17980
rect 1563 17978 1587 17980
rect 1643 17978 1667 17980
rect 1723 17978 1729 17980
rect 1483 17926 1485 17978
rect 1665 17926 1667 17978
rect 1421 17924 1427 17926
rect 1483 17924 1507 17926
rect 1563 17924 1587 17926
rect 1643 17924 1667 17926
rect 1723 17924 1729 17926
rect 1421 17915 1729 17924
rect 2364 17980 2672 17989
rect 2364 17978 2370 17980
rect 2426 17978 2450 17980
rect 2506 17978 2530 17980
rect 2586 17978 2610 17980
rect 2666 17978 2672 17980
rect 2426 17926 2428 17978
rect 2608 17926 2610 17978
rect 2364 17924 2370 17926
rect 2426 17924 2450 17926
rect 2506 17924 2530 17926
rect 2586 17924 2610 17926
rect 2666 17924 2672 17926
rect 2364 17915 2672 17924
rect 3307 17980 3615 17989
rect 3307 17978 3313 17980
rect 3369 17978 3393 17980
rect 3449 17978 3473 17980
rect 3529 17978 3553 17980
rect 3609 17978 3615 17980
rect 3369 17926 3371 17978
rect 3551 17926 3553 17978
rect 3307 17924 3313 17926
rect 3369 17924 3393 17926
rect 3449 17924 3473 17926
rect 3529 17924 3553 17926
rect 3609 17924 3615 17926
rect 3307 17915 3615 17924
rect 4250 17980 4558 17989
rect 4250 17978 4256 17980
rect 4312 17978 4336 17980
rect 4392 17978 4416 17980
rect 4472 17978 4496 17980
rect 4552 17978 4558 17980
rect 4312 17926 4314 17978
rect 4494 17926 4496 17978
rect 4250 17924 4256 17926
rect 4312 17924 4336 17926
rect 4392 17924 4416 17926
rect 4472 17924 4496 17926
rect 4552 17924 4558 17926
rect 4250 17915 4558 17924
rect 1892 17436 2200 17445
rect 1892 17434 1898 17436
rect 1954 17434 1978 17436
rect 2034 17434 2058 17436
rect 2114 17434 2138 17436
rect 2194 17434 2200 17436
rect 1954 17382 1956 17434
rect 2136 17382 2138 17434
rect 1892 17380 1898 17382
rect 1954 17380 1978 17382
rect 2034 17380 2058 17382
rect 2114 17380 2138 17382
rect 2194 17380 2200 17382
rect 1892 17371 2200 17380
rect 2835 17436 3143 17445
rect 2835 17434 2841 17436
rect 2897 17434 2921 17436
rect 2977 17434 3001 17436
rect 3057 17434 3081 17436
rect 3137 17434 3143 17436
rect 2897 17382 2899 17434
rect 3079 17382 3081 17434
rect 2835 17380 2841 17382
rect 2897 17380 2921 17382
rect 2977 17380 3001 17382
rect 3057 17380 3081 17382
rect 3137 17380 3143 17382
rect 2835 17371 3143 17380
rect 3778 17436 4086 17445
rect 3778 17434 3784 17436
rect 3840 17434 3864 17436
rect 3920 17434 3944 17436
rect 4000 17434 4024 17436
rect 4080 17434 4086 17436
rect 3840 17382 3842 17434
rect 4022 17382 4024 17434
rect 3778 17380 3784 17382
rect 3840 17380 3864 17382
rect 3920 17380 3944 17382
rect 4000 17380 4024 17382
rect 4080 17380 4086 17382
rect 3778 17371 4086 17380
rect 1421 16892 1729 16901
rect 1421 16890 1427 16892
rect 1483 16890 1507 16892
rect 1563 16890 1587 16892
rect 1643 16890 1667 16892
rect 1723 16890 1729 16892
rect 1483 16838 1485 16890
rect 1665 16838 1667 16890
rect 1421 16836 1427 16838
rect 1483 16836 1507 16838
rect 1563 16836 1587 16838
rect 1643 16836 1667 16838
rect 1723 16836 1729 16838
rect 1421 16827 1729 16836
rect 2364 16892 2672 16901
rect 2364 16890 2370 16892
rect 2426 16890 2450 16892
rect 2506 16890 2530 16892
rect 2586 16890 2610 16892
rect 2666 16890 2672 16892
rect 2426 16838 2428 16890
rect 2608 16838 2610 16890
rect 2364 16836 2370 16838
rect 2426 16836 2450 16838
rect 2506 16836 2530 16838
rect 2586 16836 2610 16838
rect 2666 16836 2672 16838
rect 2364 16827 2672 16836
rect 3307 16892 3615 16901
rect 3307 16890 3313 16892
rect 3369 16890 3393 16892
rect 3449 16890 3473 16892
rect 3529 16890 3553 16892
rect 3609 16890 3615 16892
rect 3369 16838 3371 16890
rect 3551 16838 3553 16890
rect 3307 16836 3313 16838
rect 3369 16836 3393 16838
rect 3449 16836 3473 16838
rect 3529 16836 3553 16838
rect 3609 16836 3615 16838
rect 3307 16827 3615 16836
rect 4250 16892 4558 16901
rect 4250 16890 4256 16892
rect 4312 16890 4336 16892
rect 4392 16890 4416 16892
rect 4472 16890 4496 16892
rect 4552 16890 4558 16892
rect 4312 16838 4314 16890
rect 4494 16838 4496 16890
rect 4250 16836 4256 16838
rect 4312 16836 4336 16838
rect 4392 16836 4416 16838
rect 4472 16836 4496 16838
rect 4552 16836 4558 16838
rect 4250 16827 4558 16836
rect 1892 16348 2200 16357
rect 1892 16346 1898 16348
rect 1954 16346 1978 16348
rect 2034 16346 2058 16348
rect 2114 16346 2138 16348
rect 2194 16346 2200 16348
rect 1954 16294 1956 16346
rect 2136 16294 2138 16346
rect 1892 16292 1898 16294
rect 1954 16292 1978 16294
rect 2034 16292 2058 16294
rect 2114 16292 2138 16294
rect 2194 16292 2200 16294
rect 1892 16283 2200 16292
rect 2835 16348 3143 16357
rect 2835 16346 2841 16348
rect 2897 16346 2921 16348
rect 2977 16346 3001 16348
rect 3057 16346 3081 16348
rect 3137 16346 3143 16348
rect 2897 16294 2899 16346
rect 3079 16294 3081 16346
rect 2835 16292 2841 16294
rect 2897 16292 2921 16294
rect 2977 16292 3001 16294
rect 3057 16292 3081 16294
rect 3137 16292 3143 16294
rect 2835 16283 3143 16292
rect 3778 16348 4086 16357
rect 3778 16346 3784 16348
rect 3840 16346 3864 16348
rect 3920 16346 3944 16348
rect 4000 16346 4024 16348
rect 4080 16346 4086 16348
rect 3840 16294 3842 16346
rect 4022 16294 4024 16346
rect 3778 16292 3784 16294
rect 3840 16292 3864 16294
rect 3920 16292 3944 16294
rect 4000 16292 4024 16294
rect 4080 16292 4086 16294
rect 3778 16283 4086 16292
rect 1421 15804 1729 15813
rect 1421 15802 1427 15804
rect 1483 15802 1507 15804
rect 1563 15802 1587 15804
rect 1643 15802 1667 15804
rect 1723 15802 1729 15804
rect 1483 15750 1485 15802
rect 1665 15750 1667 15802
rect 1421 15748 1427 15750
rect 1483 15748 1507 15750
rect 1563 15748 1587 15750
rect 1643 15748 1667 15750
rect 1723 15748 1729 15750
rect 1421 15739 1729 15748
rect 2364 15804 2672 15813
rect 2364 15802 2370 15804
rect 2426 15802 2450 15804
rect 2506 15802 2530 15804
rect 2586 15802 2610 15804
rect 2666 15802 2672 15804
rect 2426 15750 2428 15802
rect 2608 15750 2610 15802
rect 2364 15748 2370 15750
rect 2426 15748 2450 15750
rect 2506 15748 2530 15750
rect 2586 15748 2610 15750
rect 2666 15748 2672 15750
rect 2364 15739 2672 15748
rect 3307 15804 3615 15813
rect 3307 15802 3313 15804
rect 3369 15802 3393 15804
rect 3449 15802 3473 15804
rect 3529 15802 3553 15804
rect 3609 15802 3615 15804
rect 3369 15750 3371 15802
rect 3551 15750 3553 15802
rect 3307 15748 3313 15750
rect 3369 15748 3393 15750
rect 3449 15748 3473 15750
rect 3529 15748 3553 15750
rect 3609 15748 3615 15750
rect 3307 15739 3615 15748
rect 4250 15804 4558 15813
rect 4250 15802 4256 15804
rect 4312 15802 4336 15804
rect 4392 15802 4416 15804
rect 4472 15802 4496 15804
rect 4552 15802 4558 15804
rect 4312 15750 4314 15802
rect 4494 15750 4496 15802
rect 4250 15748 4256 15750
rect 4312 15748 4336 15750
rect 4392 15748 4416 15750
rect 4472 15748 4496 15750
rect 4552 15748 4558 15750
rect 4250 15739 4558 15748
rect 3698 15600 3754 15609
rect 3698 15535 3754 15544
rect 1892 15260 2200 15269
rect 1892 15258 1898 15260
rect 1954 15258 1978 15260
rect 2034 15258 2058 15260
rect 2114 15258 2138 15260
rect 2194 15258 2200 15260
rect 1954 15206 1956 15258
rect 2136 15206 2138 15258
rect 1892 15204 1898 15206
rect 1954 15204 1978 15206
rect 2034 15204 2058 15206
rect 2114 15204 2138 15206
rect 2194 15204 2200 15206
rect 1892 15195 2200 15204
rect 2835 15260 3143 15269
rect 2835 15258 2841 15260
rect 2897 15258 2921 15260
rect 2977 15258 3001 15260
rect 3057 15258 3081 15260
rect 3137 15258 3143 15260
rect 2897 15206 2899 15258
rect 3079 15206 3081 15258
rect 2835 15204 2841 15206
rect 2897 15204 2921 15206
rect 2977 15204 3001 15206
rect 3057 15204 3081 15206
rect 3137 15204 3143 15206
rect 2835 15195 3143 15204
rect 1421 14716 1729 14725
rect 1421 14714 1427 14716
rect 1483 14714 1507 14716
rect 1563 14714 1587 14716
rect 1643 14714 1667 14716
rect 1723 14714 1729 14716
rect 1483 14662 1485 14714
rect 1665 14662 1667 14714
rect 1421 14660 1427 14662
rect 1483 14660 1507 14662
rect 1563 14660 1587 14662
rect 1643 14660 1667 14662
rect 1723 14660 1729 14662
rect 1421 14651 1729 14660
rect 2364 14716 2672 14725
rect 2364 14714 2370 14716
rect 2426 14714 2450 14716
rect 2506 14714 2530 14716
rect 2586 14714 2610 14716
rect 2666 14714 2672 14716
rect 2426 14662 2428 14714
rect 2608 14662 2610 14714
rect 2364 14660 2370 14662
rect 2426 14660 2450 14662
rect 2506 14660 2530 14662
rect 2586 14660 2610 14662
rect 2666 14660 2672 14662
rect 2364 14651 2672 14660
rect 3307 14716 3615 14725
rect 3307 14714 3313 14716
rect 3369 14714 3393 14716
rect 3449 14714 3473 14716
rect 3529 14714 3553 14716
rect 3609 14714 3615 14716
rect 3369 14662 3371 14714
rect 3551 14662 3553 14714
rect 3307 14660 3313 14662
rect 3369 14660 3393 14662
rect 3449 14660 3473 14662
rect 3529 14660 3553 14662
rect 3609 14660 3615 14662
rect 3307 14651 3615 14660
rect 1892 14172 2200 14181
rect 1892 14170 1898 14172
rect 1954 14170 1978 14172
rect 2034 14170 2058 14172
rect 2114 14170 2138 14172
rect 2194 14170 2200 14172
rect 1954 14118 1956 14170
rect 2136 14118 2138 14170
rect 1892 14116 1898 14118
rect 1954 14116 1978 14118
rect 2034 14116 2058 14118
rect 2114 14116 2138 14118
rect 2194 14116 2200 14118
rect 1892 14107 2200 14116
rect 2835 14172 3143 14181
rect 2835 14170 2841 14172
rect 2897 14170 2921 14172
rect 2977 14170 3001 14172
rect 3057 14170 3081 14172
rect 3137 14170 3143 14172
rect 2897 14118 2899 14170
rect 3079 14118 3081 14170
rect 2835 14116 2841 14118
rect 2897 14116 2921 14118
rect 2977 14116 3001 14118
rect 3057 14116 3081 14118
rect 3137 14116 3143 14118
rect 2835 14107 3143 14116
rect 1421 13628 1729 13637
rect 1421 13626 1427 13628
rect 1483 13626 1507 13628
rect 1563 13626 1587 13628
rect 1643 13626 1667 13628
rect 1723 13626 1729 13628
rect 1483 13574 1485 13626
rect 1665 13574 1667 13626
rect 1421 13572 1427 13574
rect 1483 13572 1507 13574
rect 1563 13572 1587 13574
rect 1643 13572 1667 13574
rect 1723 13572 1729 13574
rect 1421 13563 1729 13572
rect 2364 13628 2672 13637
rect 2364 13626 2370 13628
rect 2426 13626 2450 13628
rect 2506 13626 2530 13628
rect 2586 13626 2610 13628
rect 2666 13626 2672 13628
rect 2426 13574 2428 13626
rect 2608 13574 2610 13626
rect 2364 13572 2370 13574
rect 2426 13572 2450 13574
rect 2506 13572 2530 13574
rect 2586 13572 2610 13574
rect 2666 13572 2672 13574
rect 2364 13563 2672 13572
rect 3307 13628 3615 13637
rect 3307 13626 3313 13628
rect 3369 13626 3393 13628
rect 3449 13626 3473 13628
rect 3529 13626 3553 13628
rect 3609 13626 3615 13628
rect 3369 13574 3371 13626
rect 3551 13574 3553 13626
rect 3307 13572 3313 13574
rect 3369 13572 3393 13574
rect 3449 13572 3473 13574
rect 3529 13572 3553 13574
rect 3609 13572 3615 13574
rect 3307 13563 3615 13572
rect 1892 13084 2200 13093
rect 1892 13082 1898 13084
rect 1954 13082 1978 13084
rect 2034 13082 2058 13084
rect 2114 13082 2138 13084
rect 2194 13082 2200 13084
rect 1954 13030 1956 13082
rect 2136 13030 2138 13082
rect 1892 13028 1898 13030
rect 1954 13028 1978 13030
rect 2034 13028 2058 13030
rect 2114 13028 2138 13030
rect 2194 13028 2200 13030
rect 1892 13019 2200 13028
rect 2835 13084 3143 13093
rect 2835 13082 2841 13084
rect 2897 13082 2921 13084
rect 2977 13082 3001 13084
rect 3057 13082 3081 13084
rect 3137 13082 3143 13084
rect 2897 13030 2899 13082
rect 3079 13030 3081 13082
rect 2835 13028 2841 13030
rect 2897 13028 2921 13030
rect 2977 13028 3001 13030
rect 3057 13028 3081 13030
rect 3137 13028 3143 13030
rect 2835 13019 3143 13028
rect 1421 12540 1729 12549
rect 1421 12538 1427 12540
rect 1483 12538 1507 12540
rect 1563 12538 1587 12540
rect 1643 12538 1667 12540
rect 1723 12538 1729 12540
rect 1483 12486 1485 12538
rect 1665 12486 1667 12538
rect 1421 12484 1427 12486
rect 1483 12484 1507 12486
rect 1563 12484 1587 12486
rect 1643 12484 1667 12486
rect 1723 12484 1729 12486
rect 1421 12475 1729 12484
rect 2364 12540 2672 12549
rect 2364 12538 2370 12540
rect 2426 12538 2450 12540
rect 2506 12538 2530 12540
rect 2586 12538 2610 12540
rect 2666 12538 2672 12540
rect 2426 12486 2428 12538
rect 2608 12486 2610 12538
rect 2364 12484 2370 12486
rect 2426 12484 2450 12486
rect 2506 12484 2530 12486
rect 2586 12484 2610 12486
rect 2666 12484 2672 12486
rect 2364 12475 2672 12484
rect 3307 12540 3615 12549
rect 3307 12538 3313 12540
rect 3369 12538 3393 12540
rect 3449 12538 3473 12540
rect 3529 12538 3553 12540
rect 3609 12538 3615 12540
rect 3369 12486 3371 12538
rect 3551 12486 3553 12538
rect 3307 12484 3313 12486
rect 3369 12484 3393 12486
rect 3449 12484 3473 12486
rect 3529 12484 3553 12486
rect 3609 12484 3615 12486
rect 3307 12475 3615 12484
rect 1892 11996 2200 12005
rect 1892 11994 1898 11996
rect 1954 11994 1978 11996
rect 2034 11994 2058 11996
rect 2114 11994 2138 11996
rect 2194 11994 2200 11996
rect 1954 11942 1956 11994
rect 2136 11942 2138 11994
rect 1892 11940 1898 11942
rect 1954 11940 1978 11942
rect 2034 11940 2058 11942
rect 2114 11940 2138 11942
rect 2194 11940 2200 11942
rect 1892 11931 2200 11940
rect 2835 11996 3143 12005
rect 2835 11994 2841 11996
rect 2897 11994 2921 11996
rect 2977 11994 3001 11996
rect 3057 11994 3081 11996
rect 3137 11994 3143 11996
rect 2897 11942 2899 11994
rect 3079 11942 3081 11994
rect 2835 11940 2841 11942
rect 2897 11940 2921 11942
rect 2977 11940 3001 11942
rect 3057 11940 3081 11942
rect 3137 11940 3143 11942
rect 2835 11931 3143 11940
rect 3148 11892 3200 11898
rect 3148 11834 3200 11840
rect 1768 11552 1820 11558
rect 1768 11494 1820 11500
rect 1421 11452 1729 11461
rect 1421 11450 1427 11452
rect 1483 11450 1507 11452
rect 1563 11450 1587 11452
rect 1643 11450 1667 11452
rect 1723 11450 1729 11452
rect 1483 11398 1485 11450
rect 1665 11398 1667 11450
rect 1421 11396 1427 11398
rect 1483 11396 1507 11398
rect 1563 11396 1587 11398
rect 1643 11396 1667 11398
rect 1723 11396 1729 11398
rect 1421 11387 1729 11396
rect 1216 11144 1268 11150
rect 1216 11086 1268 11092
rect 1124 10056 1176 10062
rect 1124 9998 1176 10004
rect 1136 8974 1164 9998
rect 1124 8968 1176 8974
rect 1124 8910 1176 8916
rect 1136 7886 1164 8910
rect 1124 7880 1176 7886
rect 1124 7822 1176 7828
rect 1124 7744 1176 7750
rect 1124 7686 1176 7692
rect 388 1964 440 1970
rect 388 1906 440 1912
rect 400 800 428 1906
rect 1136 800 1164 7686
rect 1228 6866 1256 11086
rect 1421 10364 1729 10373
rect 1421 10362 1427 10364
rect 1483 10362 1507 10364
rect 1563 10362 1587 10364
rect 1643 10362 1667 10364
rect 1723 10362 1729 10364
rect 1483 10310 1485 10362
rect 1665 10310 1667 10362
rect 1421 10308 1427 10310
rect 1483 10308 1507 10310
rect 1563 10308 1587 10310
rect 1643 10308 1667 10310
rect 1723 10308 1729 10310
rect 1421 10299 1729 10308
rect 1308 10124 1360 10130
rect 1308 10066 1360 10072
rect 1320 8294 1348 10066
rect 1421 9276 1729 9285
rect 1421 9274 1427 9276
rect 1483 9274 1507 9276
rect 1563 9274 1587 9276
rect 1643 9274 1667 9276
rect 1723 9274 1729 9276
rect 1483 9222 1485 9274
rect 1665 9222 1667 9274
rect 1421 9220 1427 9222
rect 1483 9220 1507 9222
rect 1563 9220 1587 9222
rect 1643 9220 1667 9222
rect 1723 9220 1729 9222
rect 1421 9211 1729 9220
rect 1780 9178 1808 11494
rect 2364 11452 2672 11461
rect 2364 11450 2370 11452
rect 2426 11450 2450 11452
rect 2506 11450 2530 11452
rect 2586 11450 2610 11452
rect 2666 11450 2672 11452
rect 2426 11398 2428 11450
rect 2608 11398 2610 11450
rect 2364 11396 2370 11398
rect 2426 11396 2450 11398
rect 2506 11396 2530 11398
rect 2586 11396 2610 11398
rect 2666 11396 2672 11398
rect 2364 11387 2672 11396
rect 3160 11370 3188 11834
rect 3307 11452 3615 11461
rect 3307 11450 3313 11452
rect 3369 11450 3393 11452
rect 3449 11450 3473 11452
rect 3529 11450 3553 11452
rect 3609 11450 3615 11452
rect 3369 11398 3371 11450
rect 3551 11398 3553 11450
rect 3307 11396 3313 11398
rect 3369 11396 3393 11398
rect 3449 11396 3473 11398
rect 3529 11396 3553 11398
rect 3609 11396 3615 11398
rect 3307 11387 3615 11396
rect 3160 11342 3280 11370
rect 2688 11144 2740 11150
rect 2688 11086 2740 11092
rect 1892 10908 2200 10917
rect 1892 10906 1898 10908
rect 1954 10906 1978 10908
rect 2034 10906 2058 10908
rect 2114 10906 2138 10908
rect 2194 10906 2200 10908
rect 1954 10854 1956 10906
rect 2136 10854 2138 10906
rect 1892 10852 1898 10854
rect 1954 10852 1978 10854
rect 2034 10852 2058 10854
rect 2114 10852 2138 10854
rect 2194 10852 2200 10854
rect 1892 10843 2200 10852
rect 2228 10804 2280 10810
rect 2228 10746 2280 10752
rect 2240 9926 2268 10746
rect 2364 10364 2672 10373
rect 2364 10362 2370 10364
rect 2426 10362 2450 10364
rect 2506 10362 2530 10364
rect 2586 10362 2610 10364
rect 2666 10362 2672 10364
rect 2426 10310 2428 10362
rect 2608 10310 2610 10362
rect 2364 10308 2370 10310
rect 2426 10308 2450 10310
rect 2506 10308 2530 10310
rect 2586 10308 2610 10310
rect 2666 10308 2672 10310
rect 2364 10299 2672 10308
rect 2228 9920 2280 9926
rect 2228 9862 2280 9868
rect 1892 9820 2200 9829
rect 1892 9818 1898 9820
rect 1954 9818 1978 9820
rect 2034 9818 2058 9820
rect 2114 9818 2138 9820
rect 2194 9818 2200 9820
rect 1954 9766 1956 9818
rect 2136 9766 2138 9818
rect 1892 9764 1898 9766
rect 1954 9764 1978 9766
rect 2034 9764 2058 9766
rect 2114 9764 2138 9766
rect 2194 9764 2200 9766
rect 1892 9755 2200 9764
rect 1768 9172 1820 9178
rect 1768 9114 1820 9120
rect 2044 9036 2096 9042
rect 2044 8978 2096 8984
rect 2056 8922 2084 8978
rect 1780 8894 2084 8922
rect 1676 8832 1728 8838
rect 1676 8774 1728 8780
rect 1688 8634 1716 8774
rect 1676 8628 1728 8634
rect 1676 8570 1728 8576
rect 1308 8288 1360 8294
rect 1308 8230 1360 8236
rect 1216 6860 1268 6866
rect 1216 6802 1268 6808
rect 1228 5778 1256 6802
rect 1216 5772 1268 5778
rect 1216 5714 1268 5720
rect 1320 5642 1348 8230
rect 1421 8188 1729 8197
rect 1421 8186 1427 8188
rect 1483 8186 1507 8188
rect 1563 8186 1587 8188
rect 1643 8186 1667 8188
rect 1723 8186 1729 8188
rect 1483 8134 1485 8186
rect 1665 8134 1667 8186
rect 1421 8132 1427 8134
rect 1483 8132 1507 8134
rect 1563 8132 1587 8134
rect 1643 8132 1667 8134
rect 1723 8132 1729 8134
rect 1421 8123 1729 8132
rect 1584 7880 1636 7886
rect 1584 7822 1636 7828
rect 1596 7478 1624 7822
rect 1780 7546 1808 8894
rect 1892 8732 2200 8741
rect 1892 8730 1898 8732
rect 1954 8730 1978 8732
rect 2034 8730 2058 8732
rect 2114 8730 2138 8732
rect 2194 8730 2200 8732
rect 1954 8678 1956 8730
rect 2136 8678 2138 8730
rect 1892 8676 1898 8678
rect 1954 8676 1978 8678
rect 2034 8676 2058 8678
rect 2114 8676 2138 8678
rect 2194 8676 2200 8678
rect 1892 8667 2200 8676
rect 2136 8628 2188 8634
rect 2136 8570 2188 8576
rect 2148 8514 2176 8570
rect 2240 8514 2268 9862
rect 2700 9382 2728 11086
rect 2835 10908 3143 10917
rect 2835 10906 2841 10908
rect 2897 10906 2921 10908
rect 2977 10906 3001 10908
rect 3057 10906 3081 10908
rect 3137 10906 3143 10908
rect 2897 10854 2899 10906
rect 3079 10854 3081 10906
rect 2835 10852 2841 10854
rect 2897 10852 2921 10854
rect 2977 10852 3001 10854
rect 3057 10852 3081 10854
rect 3137 10852 3143 10854
rect 2835 10843 3143 10852
rect 3252 10810 3280 11342
rect 3424 11280 3476 11286
rect 3422 11248 3424 11257
rect 3476 11248 3478 11257
rect 3422 11183 3478 11192
rect 3240 10804 3292 10810
rect 3240 10746 3292 10752
rect 3148 10464 3200 10470
rect 3148 10406 3200 10412
rect 3160 10282 3188 10406
rect 3307 10364 3615 10373
rect 3307 10362 3313 10364
rect 3369 10362 3393 10364
rect 3449 10362 3473 10364
rect 3529 10362 3553 10364
rect 3609 10362 3615 10364
rect 3369 10310 3371 10362
rect 3551 10310 3553 10362
rect 3307 10308 3313 10310
rect 3369 10308 3393 10310
rect 3449 10308 3473 10310
rect 3529 10308 3553 10310
rect 3609 10308 3615 10310
rect 3307 10299 3615 10308
rect 3160 10254 3280 10282
rect 2835 9820 3143 9829
rect 2835 9818 2841 9820
rect 2897 9818 2921 9820
rect 2977 9818 3001 9820
rect 3057 9818 3081 9820
rect 3137 9818 3143 9820
rect 2897 9766 2899 9818
rect 3079 9766 3081 9818
rect 2835 9764 2841 9766
rect 2897 9764 2921 9766
rect 2977 9764 3001 9766
rect 3057 9764 3081 9766
rect 3137 9764 3143 9766
rect 2835 9755 3143 9764
rect 3252 9602 3280 10254
rect 3608 9988 3660 9994
rect 3608 9930 3660 9936
rect 3160 9586 3280 9602
rect 3160 9580 3292 9586
rect 3160 9574 3240 9580
rect 2688 9376 2740 9382
rect 2688 9318 2740 9324
rect 2364 9276 2672 9285
rect 2364 9274 2370 9276
rect 2426 9274 2450 9276
rect 2506 9274 2530 9276
rect 2586 9274 2610 9276
rect 2666 9274 2672 9276
rect 2426 9222 2428 9274
rect 2608 9222 2610 9274
rect 2364 9220 2370 9222
rect 2426 9220 2450 9222
rect 2506 9220 2530 9222
rect 2586 9220 2610 9222
rect 2666 9220 2672 9222
rect 2364 9211 2672 9220
rect 2148 8486 2268 8514
rect 1860 7948 1912 7954
rect 1860 7890 1912 7896
rect 1872 7750 1900 7890
rect 2148 7834 2176 8486
rect 2364 8188 2672 8197
rect 2364 8186 2370 8188
rect 2426 8186 2450 8188
rect 2506 8186 2530 8188
rect 2586 8186 2610 8188
rect 2666 8186 2672 8188
rect 2426 8134 2428 8186
rect 2608 8134 2610 8186
rect 2364 8132 2370 8134
rect 2426 8132 2450 8134
rect 2506 8132 2530 8134
rect 2586 8132 2610 8134
rect 2666 8132 2672 8134
rect 2364 8123 2672 8132
rect 2056 7806 2268 7834
rect 2056 7750 2084 7806
rect 1860 7744 1912 7750
rect 1860 7686 1912 7692
rect 2044 7744 2096 7750
rect 2044 7686 2096 7692
rect 2240 7698 2268 7806
rect 2240 7670 2360 7698
rect 1892 7644 2200 7653
rect 1892 7642 1898 7644
rect 1954 7642 1978 7644
rect 2034 7642 2058 7644
rect 2114 7642 2138 7644
rect 2194 7642 2200 7644
rect 1954 7590 1956 7642
rect 2136 7590 2138 7642
rect 1892 7588 1898 7590
rect 1954 7588 1978 7590
rect 2034 7588 2058 7590
rect 2114 7588 2138 7590
rect 2194 7588 2200 7590
rect 1892 7579 2200 7588
rect 1768 7540 1820 7546
rect 1768 7482 1820 7488
rect 1584 7472 1636 7478
rect 1584 7414 1636 7420
rect 1421 7100 1729 7109
rect 1421 7098 1427 7100
rect 1483 7098 1507 7100
rect 1563 7098 1587 7100
rect 1643 7098 1667 7100
rect 1723 7098 1729 7100
rect 1483 7046 1485 7098
rect 1665 7046 1667 7098
rect 1421 7044 1427 7046
rect 1483 7044 1507 7046
rect 1563 7044 1587 7046
rect 1643 7044 1667 7046
rect 1723 7044 1729 7046
rect 1421 7035 1729 7044
rect 1780 6118 1808 7482
rect 2332 7478 2360 7670
rect 2228 7472 2280 7478
rect 2228 7414 2280 7420
rect 2320 7472 2372 7478
rect 2320 7414 2372 7420
rect 1892 6556 2200 6565
rect 1892 6554 1898 6556
rect 1954 6554 1978 6556
rect 2034 6554 2058 6556
rect 2114 6554 2138 6556
rect 2194 6554 2200 6556
rect 1954 6502 1956 6554
rect 2136 6502 2138 6554
rect 1892 6500 1898 6502
rect 1954 6500 1978 6502
rect 2034 6500 2058 6502
rect 2114 6500 2138 6502
rect 2194 6500 2200 6502
rect 1892 6491 2200 6500
rect 2240 6254 2268 7414
rect 2364 7100 2672 7109
rect 2364 7098 2370 7100
rect 2426 7098 2450 7100
rect 2506 7098 2530 7100
rect 2586 7098 2610 7100
rect 2666 7098 2672 7100
rect 2426 7046 2428 7098
rect 2608 7046 2610 7098
rect 2364 7044 2370 7046
rect 2426 7044 2450 7046
rect 2506 7044 2530 7046
rect 2586 7044 2610 7046
rect 2666 7044 2672 7046
rect 2364 7035 2672 7044
rect 2596 6724 2648 6730
rect 2596 6666 2648 6672
rect 2228 6248 2280 6254
rect 2228 6190 2280 6196
rect 2608 6202 2636 6666
rect 2700 6390 2728 9318
rect 3160 9194 3188 9574
rect 3240 9522 3292 9528
rect 3620 9518 3648 9930
rect 3608 9512 3660 9518
rect 3608 9454 3660 9460
rect 3307 9276 3615 9285
rect 3307 9274 3313 9276
rect 3369 9274 3393 9276
rect 3449 9274 3473 9276
rect 3529 9274 3553 9276
rect 3609 9274 3615 9276
rect 3369 9222 3371 9274
rect 3551 9222 3553 9274
rect 3307 9220 3313 9222
rect 3369 9220 3393 9222
rect 3449 9220 3473 9222
rect 3529 9220 3553 9222
rect 3609 9220 3615 9222
rect 3307 9211 3615 9220
rect 3160 9166 3280 9194
rect 2835 8732 3143 8741
rect 2835 8730 2841 8732
rect 2897 8730 2921 8732
rect 2977 8730 3001 8732
rect 3057 8730 3081 8732
rect 3137 8730 3143 8732
rect 2897 8678 2899 8730
rect 3079 8678 3081 8730
rect 2835 8676 2841 8678
rect 2897 8676 2921 8678
rect 2977 8676 3001 8678
rect 3057 8676 3081 8678
rect 3137 8676 3143 8678
rect 2835 8667 3143 8676
rect 3252 8514 3280 9166
rect 3516 9172 3568 9178
rect 3516 9114 3568 9120
rect 3608 9172 3660 9178
rect 3608 9114 3660 9120
rect 3160 8486 3280 8514
rect 3160 8106 3188 8486
rect 3528 8430 3556 9114
rect 3620 8634 3648 9114
rect 3712 9042 3740 15535
rect 3778 15260 4086 15269
rect 3778 15258 3784 15260
rect 3840 15258 3864 15260
rect 3920 15258 3944 15260
rect 4000 15258 4024 15260
rect 4080 15258 4086 15260
rect 3840 15206 3842 15258
rect 4022 15206 4024 15258
rect 3778 15204 3784 15206
rect 3840 15204 3864 15206
rect 3920 15204 3944 15206
rect 4000 15204 4024 15206
rect 4080 15204 4086 15206
rect 3778 15195 4086 15204
rect 4250 14716 4558 14725
rect 4250 14714 4256 14716
rect 4312 14714 4336 14716
rect 4392 14714 4416 14716
rect 4472 14714 4496 14716
rect 4552 14714 4558 14716
rect 4312 14662 4314 14714
rect 4494 14662 4496 14714
rect 4250 14660 4256 14662
rect 4312 14660 4336 14662
rect 4392 14660 4416 14662
rect 4472 14660 4496 14662
rect 4552 14660 4558 14662
rect 4250 14651 4558 14660
rect 3778 14172 4086 14181
rect 3778 14170 3784 14172
rect 3840 14170 3864 14172
rect 3920 14170 3944 14172
rect 4000 14170 4024 14172
rect 4080 14170 4086 14172
rect 3840 14118 3842 14170
rect 4022 14118 4024 14170
rect 3778 14116 3784 14118
rect 3840 14116 3864 14118
rect 3920 14116 3944 14118
rect 4000 14116 4024 14118
rect 4080 14116 4086 14118
rect 3778 14107 4086 14116
rect 4250 13628 4558 13637
rect 4250 13626 4256 13628
rect 4312 13626 4336 13628
rect 4392 13626 4416 13628
rect 4472 13626 4496 13628
rect 4552 13626 4558 13628
rect 4312 13574 4314 13626
rect 4494 13574 4496 13626
rect 4250 13572 4256 13574
rect 4312 13572 4336 13574
rect 4392 13572 4416 13574
rect 4472 13572 4496 13574
rect 4552 13572 4558 13574
rect 4250 13563 4558 13572
rect 3778 13084 4086 13093
rect 3778 13082 3784 13084
rect 3840 13082 3864 13084
rect 3920 13082 3944 13084
rect 4000 13082 4024 13084
rect 4080 13082 4086 13084
rect 3840 13030 3842 13082
rect 4022 13030 4024 13082
rect 3778 13028 3784 13030
rect 3840 13028 3864 13030
rect 3920 13028 3944 13030
rect 4000 13028 4024 13030
rect 4080 13028 4086 13030
rect 3778 13019 4086 13028
rect 4250 12540 4558 12549
rect 4250 12538 4256 12540
rect 4312 12538 4336 12540
rect 4392 12538 4416 12540
rect 4472 12538 4496 12540
rect 4552 12538 4558 12540
rect 4312 12486 4314 12538
rect 4494 12486 4496 12538
rect 4250 12484 4256 12486
rect 4312 12484 4336 12486
rect 4392 12484 4416 12486
rect 4472 12484 4496 12486
rect 4552 12484 4558 12486
rect 4250 12475 4558 12484
rect 3778 11996 4086 12005
rect 3778 11994 3784 11996
rect 3840 11994 3864 11996
rect 3920 11994 3944 11996
rect 4000 11994 4024 11996
rect 4080 11994 4086 11996
rect 3840 11942 3842 11994
rect 4022 11942 4024 11994
rect 3778 11940 3784 11942
rect 3840 11940 3864 11942
rect 3920 11940 3944 11942
rect 4000 11940 4024 11942
rect 4080 11940 4086 11942
rect 3778 11931 4086 11940
rect 3884 11688 3936 11694
rect 3884 11630 3936 11636
rect 4160 11688 4212 11694
rect 4160 11630 4212 11636
rect 3896 11558 3924 11630
rect 3884 11552 3936 11558
rect 3884 11494 3936 11500
rect 3778 10908 4086 10917
rect 3778 10906 3784 10908
rect 3840 10906 3864 10908
rect 3920 10906 3944 10908
rect 4000 10906 4024 10908
rect 4080 10906 4086 10908
rect 3840 10854 3842 10906
rect 4022 10854 4024 10906
rect 3778 10852 3784 10854
rect 3840 10852 3864 10854
rect 3920 10852 3944 10854
rect 4000 10852 4024 10854
rect 4080 10852 4086 10854
rect 3778 10843 4086 10852
rect 4172 10606 4200 11630
rect 4250 11452 4558 11461
rect 4250 11450 4256 11452
rect 4312 11450 4336 11452
rect 4392 11450 4416 11452
rect 4472 11450 4496 11452
rect 4552 11450 4558 11452
rect 4312 11398 4314 11450
rect 4494 11398 4496 11450
rect 4250 11396 4256 11398
rect 4312 11396 4336 11398
rect 4392 11396 4416 11398
rect 4472 11396 4496 11398
rect 4552 11396 4558 11398
rect 4250 11387 4558 11396
rect 3884 10600 3936 10606
rect 3884 10542 3936 10548
rect 4160 10600 4212 10606
rect 4160 10542 4212 10548
rect 3896 9926 3924 10542
rect 3884 9920 3936 9926
rect 3884 9862 3936 9868
rect 3778 9820 4086 9829
rect 3778 9818 3784 9820
rect 3840 9818 3864 9820
rect 3920 9818 3944 9820
rect 4000 9818 4024 9820
rect 4080 9818 4086 9820
rect 3840 9766 3842 9818
rect 4022 9766 4024 9818
rect 3778 9764 3784 9766
rect 3840 9764 3864 9766
rect 3920 9764 3944 9766
rect 4000 9764 4024 9766
rect 4080 9764 4086 9766
rect 3778 9755 4086 9764
rect 3884 9716 3936 9722
rect 3884 9658 3936 9664
rect 3792 9376 3844 9382
rect 3792 9318 3844 9324
rect 3700 9036 3752 9042
rect 3700 8978 3752 8984
rect 3804 8922 3832 9318
rect 3896 9178 3924 9658
rect 4172 9518 4200 10542
rect 4250 10364 4558 10373
rect 4250 10362 4256 10364
rect 4312 10362 4336 10364
rect 4392 10362 4416 10364
rect 4472 10362 4496 10364
rect 4552 10362 4558 10364
rect 4312 10310 4314 10362
rect 4494 10310 4496 10362
rect 4250 10308 4256 10310
rect 4312 10308 4336 10310
rect 4392 10308 4416 10310
rect 4472 10308 4496 10310
rect 4552 10308 4558 10310
rect 4250 10299 4558 10308
rect 4632 10010 4660 18663
rect 4721 18524 5029 18533
rect 4721 18522 4727 18524
rect 4783 18522 4807 18524
rect 4863 18522 4887 18524
rect 4943 18522 4967 18524
rect 5023 18522 5029 18524
rect 4783 18470 4785 18522
rect 4965 18470 4967 18522
rect 4721 18468 4727 18470
rect 4783 18468 4807 18470
rect 4863 18468 4887 18470
rect 4943 18468 4967 18470
rect 5023 18468 5029 18470
rect 4721 18459 5029 18468
rect 4721 17436 5029 17445
rect 4721 17434 4727 17436
rect 4783 17434 4807 17436
rect 4863 17434 4887 17436
rect 4943 17434 4967 17436
rect 5023 17434 5029 17436
rect 4783 17382 4785 17434
rect 4965 17382 4967 17434
rect 4721 17380 4727 17382
rect 4783 17380 4807 17382
rect 4863 17380 4887 17382
rect 4943 17380 4967 17382
rect 5023 17380 5029 17382
rect 4721 17371 5029 17380
rect 5078 17232 5134 17241
rect 5078 17167 5134 17176
rect 4721 16348 5029 16357
rect 4721 16346 4727 16348
rect 4783 16346 4807 16348
rect 4863 16346 4887 16348
rect 4943 16346 4967 16348
rect 5023 16346 5029 16348
rect 4783 16294 4785 16346
rect 4965 16294 4967 16346
rect 4721 16292 4727 16294
rect 4783 16292 4807 16294
rect 4863 16292 4887 16294
rect 4943 16292 4967 16294
rect 5023 16292 5029 16294
rect 4721 16283 5029 16292
rect 4721 15260 5029 15269
rect 4721 15258 4727 15260
rect 4783 15258 4807 15260
rect 4863 15258 4887 15260
rect 4943 15258 4967 15260
rect 5023 15258 5029 15260
rect 4783 15206 4785 15258
rect 4965 15206 4967 15258
rect 4721 15204 4727 15206
rect 4783 15204 4807 15206
rect 4863 15204 4887 15206
rect 4943 15204 4967 15206
rect 5023 15204 5029 15206
rect 4721 15195 5029 15204
rect 4721 14172 5029 14181
rect 4721 14170 4727 14172
rect 4783 14170 4807 14172
rect 4863 14170 4887 14172
rect 4943 14170 4967 14172
rect 5023 14170 5029 14172
rect 4783 14118 4785 14170
rect 4965 14118 4967 14170
rect 4721 14116 4727 14118
rect 4783 14116 4807 14118
rect 4863 14116 4887 14118
rect 4943 14116 4967 14118
rect 5023 14116 5029 14118
rect 4721 14107 5029 14116
rect 4721 13084 5029 13093
rect 4721 13082 4727 13084
rect 4783 13082 4807 13084
rect 4863 13082 4887 13084
rect 4943 13082 4967 13084
rect 5023 13082 5029 13084
rect 4783 13030 4785 13082
rect 4965 13030 4967 13082
rect 4721 13028 4727 13030
rect 4783 13028 4807 13030
rect 4863 13028 4887 13030
rect 4943 13028 4967 13030
rect 5023 13028 5029 13030
rect 4721 13019 5029 13028
rect 4721 11996 5029 12005
rect 4721 11994 4727 11996
rect 4783 11994 4807 11996
rect 4863 11994 4887 11996
rect 4943 11994 4967 11996
rect 5023 11994 5029 11996
rect 4783 11942 4785 11994
rect 4965 11942 4967 11994
rect 4721 11940 4727 11942
rect 4783 11940 4807 11942
rect 4863 11940 4887 11942
rect 4943 11940 4967 11942
rect 5023 11940 5029 11942
rect 4721 11931 5029 11940
rect 5092 11762 5120 17167
rect 5080 11756 5132 11762
rect 5080 11698 5132 11704
rect 5080 11552 5132 11558
rect 5080 11494 5132 11500
rect 4721 10908 5029 10917
rect 4721 10906 4727 10908
rect 4783 10906 4807 10908
rect 4863 10906 4887 10908
rect 4943 10906 4967 10908
rect 5023 10906 5029 10908
rect 4783 10854 4785 10906
rect 4965 10854 4967 10906
rect 4721 10852 4727 10854
rect 4783 10852 4807 10854
rect 4863 10852 4887 10854
rect 4943 10852 4967 10854
rect 5023 10852 5029 10854
rect 4721 10843 5029 10852
rect 4540 9982 4660 10010
rect 4160 9512 4212 9518
rect 4160 9454 4212 9460
rect 3884 9172 3936 9178
rect 3884 9114 3936 9120
rect 3712 8894 3832 8922
rect 3608 8628 3660 8634
rect 3608 8570 3660 8576
rect 3712 8498 3740 8894
rect 3778 8732 4086 8741
rect 3778 8730 3784 8732
rect 3840 8730 3864 8732
rect 3920 8730 3944 8732
rect 4000 8730 4024 8732
rect 4080 8730 4086 8732
rect 3840 8678 3842 8730
rect 4022 8678 4024 8730
rect 3778 8676 3784 8678
rect 3840 8676 3864 8678
rect 3920 8676 3944 8678
rect 4000 8676 4024 8678
rect 4080 8676 4086 8678
rect 3778 8667 4086 8676
rect 3700 8492 3752 8498
rect 3700 8434 3752 8440
rect 4172 8430 4200 9454
rect 4540 9382 4568 9982
rect 4620 9920 4672 9926
rect 4620 9862 4672 9868
rect 4528 9376 4580 9382
rect 4528 9318 4580 9324
rect 4250 9276 4558 9285
rect 4250 9274 4256 9276
rect 4312 9274 4336 9276
rect 4392 9274 4416 9276
rect 4472 9274 4496 9276
rect 4552 9274 4558 9276
rect 4312 9222 4314 9274
rect 4494 9222 4496 9274
rect 4250 9220 4256 9222
rect 4312 9220 4336 9222
rect 4392 9220 4416 9222
rect 4472 9220 4496 9222
rect 4552 9220 4558 9222
rect 4250 9211 4558 9220
rect 3516 8424 3568 8430
rect 3516 8366 3568 8372
rect 4160 8424 4212 8430
rect 4160 8366 4212 8372
rect 3307 8188 3615 8197
rect 3307 8186 3313 8188
rect 3369 8186 3393 8188
rect 3449 8186 3473 8188
rect 3529 8186 3553 8188
rect 3609 8186 3615 8188
rect 3369 8134 3371 8186
rect 3551 8134 3553 8186
rect 3307 8132 3313 8134
rect 3369 8132 3393 8134
rect 3449 8132 3473 8134
rect 3529 8132 3553 8134
rect 3609 8132 3615 8134
rect 3307 8123 3615 8132
rect 3160 8078 3280 8106
rect 2835 7644 3143 7653
rect 2835 7642 2841 7644
rect 2897 7642 2921 7644
rect 2977 7642 3001 7644
rect 3057 7642 3081 7644
rect 3137 7642 3143 7644
rect 2897 7590 2899 7642
rect 3079 7590 3081 7642
rect 2835 7588 2841 7590
rect 2897 7588 2921 7590
rect 2977 7588 3001 7590
rect 3057 7588 3081 7590
rect 3137 7588 3143 7590
rect 2835 7579 3143 7588
rect 2780 7472 2832 7478
rect 3252 7426 3280 8078
rect 3700 7744 3752 7750
rect 3700 7686 3752 7692
rect 2780 7414 2832 7420
rect 2792 6730 2820 7414
rect 3160 7398 3280 7426
rect 3160 6798 3188 7398
rect 3712 7342 3740 7686
rect 3778 7644 4086 7653
rect 3778 7642 3784 7644
rect 3840 7642 3864 7644
rect 3920 7642 3944 7644
rect 4000 7642 4024 7644
rect 4080 7642 4086 7644
rect 3840 7590 3842 7642
rect 4022 7590 4024 7642
rect 3778 7588 3784 7590
rect 3840 7588 3864 7590
rect 3920 7588 3944 7590
rect 4000 7588 4024 7590
rect 4080 7588 4086 7590
rect 3778 7579 4086 7588
rect 4172 7342 4200 8366
rect 4250 8188 4558 8197
rect 4250 8186 4256 8188
rect 4312 8186 4336 8188
rect 4392 8186 4416 8188
rect 4472 8186 4496 8188
rect 4552 8186 4558 8188
rect 4312 8134 4314 8186
rect 4494 8134 4496 8186
rect 4250 8132 4256 8134
rect 4312 8132 4336 8134
rect 4392 8132 4416 8134
rect 4472 8132 4496 8134
rect 4552 8132 4558 8134
rect 4250 8123 4558 8132
rect 3700 7336 3752 7342
rect 3700 7278 3752 7284
rect 4160 7336 4212 7342
rect 4160 7278 4212 7284
rect 3307 7100 3615 7109
rect 3307 7098 3313 7100
rect 3369 7098 3393 7100
rect 3449 7098 3473 7100
rect 3529 7098 3553 7100
rect 3609 7098 3615 7100
rect 3369 7046 3371 7098
rect 3551 7046 3553 7098
rect 3307 7044 3313 7046
rect 3369 7044 3393 7046
rect 3449 7044 3473 7046
rect 3529 7044 3553 7046
rect 3609 7044 3615 7046
rect 3307 7035 3615 7044
rect 3712 6882 3740 7278
rect 3528 6854 3740 6882
rect 3148 6792 3200 6798
rect 3148 6734 3200 6740
rect 2780 6724 2832 6730
rect 2780 6666 2832 6672
rect 2835 6556 3143 6565
rect 2835 6554 2841 6556
rect 2897 6554 2921 6556
rect 2977 6554 3001 6556
rect 3057 6554 3081 6556
rect 3137 6554 3143 6556
rect 2897 6502 2899 6554
rect 3079 6502 3081 6554
rect 2835 6500 2841 6502
rect 2897 6500 2921 6502
rect 2977 6500 3001 6502
rect 3057 6500 3081 6502
rect 3137 6500 3143 6502
rect 2835 6491 3143 6500
rect 2688 6384 2740 6390
rect 3528 6361 3556 6854
rect 3606 6760 3662 6769
rect 3606 6695 3662 6704
rect 2688 6326 2740 6332
rect 3514 6352 3570 6361
rect 3514 6287 3570 6296
rect 3620 6202 3648 6695
rect 3700 6656 3752 6662
rect 3700 6598 3752 6604
rect 3712 6322 3740 6598
rect 3778 6556 4086 6565
rect 3778 6554 3784 6556
rect 3840 6554 3864 6556
rect 3920 6554 3944 6556
rect 4000 6554 4024 6556
rect 4080 6554 4086 6556
rect 3840 6502 3842 6554
rect 4022 6502 4024 6554
rect 3778 6500 3784 6502
rect 3840 6500 3864 6502
rect 3920 6500 3944 6502
rect 4000 6500 4024 6502
rect 4080 6500 4086 6502
rect 3778 6491 4086 6500
rect 3790 6352 3846 6361
rect 3700 6316 3752 6322
rect 3790 6287 3846 6296
rect 3700 6258 3752 6264
rect 2608 6174 2728 6202
rect 3620 6174 3740 6202
rect 1768 6112 1820 6118
rect 1768 6054 1820 6060
rect 2228 6112 2280 6118
rect 2228 6054 2280 6060
rect 1421 6012 1729 6021
rect 1421 6010 1427 6012
rect 1483 6010 1507 6012
rect 1563 6010 1587 6012
rect 1643 6010 1667 6012
rect 1723 6010 1729 6012
rect 1483 5958 1485 6010
rect 1665 5958 1667 6010
rect 1421 5956 1427 5958
rect 1483 5956 1507 5958
rect 1563 5956 1587 5958
rect 1643 5956 1667 5958
rect 1723 5956 1729 5958
rect 1421 5947 1729 5956
rect 1768 5772 1820 5778
rect 1768 5714 1820 5720
rect 1308 5636 1360 5642
rect 1308 5578 1360 5584
rect 1780 5250 1808 5714
rect 1892 5468 2200 5477
rect 1892 5466 1898 5468
rect 1954 5466 1978 5468
rect 2034 5466 2058 5468
rect 2114 5466 2138 5468
rect 2194 5466 2200 5468
rect 1954 5414 1956 5466
rect 2136 5414 2138 5466
rect 1892 5412 1898 5414
rect 1954 5412 1978 5414
rect 2034 5412 2058 5414
rect 2114 5412 2138 5414
rect 2194 5412 2200 5414
rect 1892 5403 2200 5412
rect 1780 5222 1900 5250
rect 2240 5234 2268 6054
rect 2364 6012 2672 6021
rect 2364 6010 2370 6012
rect 2426 6010 2450 6012
rect 2506 6010 2530 6012
rect 2586 6010 2610 6012
rect 2666 6010 2672 6012
rect 2426 5958 2428 6010
rect 2608 5958 2610 6010
rect 2364 5956 2370 5958
rect 2426 5956 2450 5958
rect 2506 5956 2530 5958
rect 2586 5956 2610 5958
rect 2666 5956 2672 5958
rect 2364 5947 2672 5956
rect 1872 5166 1900 5222
rect 2228 5228 2280 5234
rect 2228 5170 2280 5176
rect 1860 5160 1912 5166
rect 2700 5114 2728 6174
rect 3307 6012 3615 6021
rect 3307 6010 3313 6012
rect 3369 6010 3393 6012
rect 3449 6010 3473 6012
rect 3529 6010 3553 6012
rect 3609 6010 3615 6012
rect 3369 5958 3371 6010
rect 3551 5958 3553 6010
rect 3307 5956 3313 5958
rect 3369 5956 3393 5958
rect 3449 5956 3473 5958
rect 3529 5956 3553 5958
rect 3609 5956 3615 5958
rect 3307 5947 3615 5956
rect 3712 5914 3740 6174
rect 3700 5908 3752 5914
rect 3700 5850 3752 5856
rect 3240 5840 3292 5846
rect 3240 5782 3292 5788
rect 2835 5468 3143 5477
rect 2835 5466 2841 5468
rect 2897 5466 2921 5468
rect 2977 5466 3001 5468
rect 3057 5466 3081 5468
rect 3137 5466 3143 5468
rect 2897 5414 2899 5466
rect 3079 5414 3081 5466
rect 2835 5412 2841 5414
rect 2897 5412 2921 5414
rect 2977 5412 3001 5414
rect 3057 5412 3081 5414
rect 3137 5412 3143 5414
rect 2835 5403 3143 5412
rect 3252 5234 3280 5782
rect 3804 5534 3832 6287
rect 4172 6254 4200 7278
rect 4250 7100 4558 7109
rect 4250 7098 4256 7100
rect 4312 7098 4336 7100
rect 4392 7098 4416 7100
rect 4472 7098 4496 7100
rect 4552 7098 4558 7100
rect 4312 7046 4314 7098
rect 4494 7046 4496 7098
rect 4250 7044 4256 7046
rect 4312 7044 4336 7046
rect 4392 7044 4416 7046
rect 4472 7044 4496 7046
rect 4552 7044 4558 7046
rect 4250 7035 4558 7044
rect 4632 6338 4660 9862
rect 4721 9820 5029 9829
rect 4721 9818 4727 9820
rect 4783 9818 4807 9820
rect 4863 9818 4887 9820
rect 4943 9818 4967 9820
rect 5023 9818 5029 9820
rect 4783 9766 4785 9818
rect 4965 9766 4967 9818
rect 4721 9764 4727 9766
rect 4783 9764 4807 9766
rect 4863 9764 4887 9766
rect 4943 9764 4967 9766
rect 5023 9764 5029 9766
rect 4721 9755 5029 9764
rect 5092 8838 5120 11494
rect 5184 10674 5212 21383
rect 5172 10668 5224 10674
rect 5172 10610 5224 10616
rect 5276 9994 5304 23174
rect 5538 19952 5594 19961
rect 5538 19887 5594 19896
rect 5354 14512 5410 14521
rect 5354 14447 5410 14456
rect 5264 9988 5316 9994
rect 5264 9930 5316 9936
rect 5170 9480 5226 9489
rect 5170 9415 5226 9424
rect 5080 8832 5132 8838
rect 5080 8774 5132 8780
rect 4721 8732 5029 8741
rect 4721 8730 4727 8732
rect 4783 8730 4807 8732
rect 4863 8730 4887 8732
rect 4943 8730 4967 8732
rect 5023 8730 5029 8732
rect 4783 8678 4785 8730
rect 4965 8678 4967 8730
rect 4721 8676 4727 8678
rect 4783 8676 4807 8678
rect 4863 8676 4887 8678
rect 4943 8676 4967 8678
rect 5023 8676 5029 8678
rect 4721 8667 5029 8676
rect 5078 8256 5134 8265
rect 5078 8191 5134 8200
rect 4721 7644 5029 7653
rect 4721 7642 4727 7644
rect 4783 7642 4807 7644
rect 4863 7642 4887 7644
rect 4943 7642 4967 7644
rect 5023 7642 5029 7644
rect 4783 7590 4785 7642
rect 4965 7590 4967 7642
rect 4721 7588 4727 7590
rect 4783 7588 4807 7590
rect 4863 7588 4887 7590
rect 4943 7588 4967 7590
rect 5023 7588 5029 7590
rect 4721 7579 5029 7588
rect 4721 6556 5029 6565
rect 4721 6554 4727 6556
rect 4783 6554 4807 6556
rect 4863 6554 4887 6556
rect 4943 6554 4967 6556
rect 5023 6554 5029 6556
rect 4783 6502 4785 6554
rect 4965 6502 4967 6554
rect 4721 6500 4727 6502
rect 4783 6500 4807 6502
rect 4863 6500 4887 6502
rect 4943 6500 4967 6502
rect 5023 6500 5029 6502
rect 4721 6491 5029 6500
rect 4632 6310 4752 6338
rect 4160 6248 4212 6254
rect 4160 6190 4212 6196
rect 4620 6248 4672 6254
rect 4620 6190 4672 6196
rect 3712 5506 3832 5534
rect 3240 5228 3292 5234
rect 3240 5170 3292 5176
rect 1860 5102 1912 5108
rect 1421 4924 1729 4933
rect 1421 4922 1427 4924
rect 1483 4922 1507 4924
rect 1563 4922 1587 4924
rect 1643 4922 1667 4924
rect 1723 4922 1729 4924
rect 1483 4870 1485 4922
rect 1665 4870 1667 4922
rect 1421 4868 1427 4870
rect 1483 4868 1507 4870
rect 1563 4868 1587 4870
rect 1643 4868 1667 4870
rect 1723 4868 1729 4870
rect 1421 4859 1729 4868
rect 1872 4622 1900 5102
rect 2240 5086 2728 5114
rect 3148 5160 3200 5166
rect 3148 5102 3200 5108
rect 1860 4616 1912 4622
rect 1860 4558 1912 4564
rect 1892 4380 2200 4389
rect 1892 4378 1898 4380
rect 1954 4378 1978 4380
rect 2034 4378 2058 4380
rect 2114 4378 2138 4380
rect 2194 4378 2200 4380
rect 1954 4326 1956 4378
rect 2136 4326 2138 4378
rect 1892 4324 1898 4326
rect 1954 4324 1978 4326
rect 2034 4324 2058 4326
rect 2114 4324 2138 4326
rect 2194 4324 2200 4326
rect 1892 4315 2200 4324
rect 1421 3836 1729 3845
rect 1421 3834 1427 3836
rect 1483 3834 1507 3836
rect 1563 3834 1587 3836
rect 1643 3834 1667 3836
rect 1723 3834 1729 3836
rect 1483 3782 1485 3834
rect 1665 3782 1667 3834
rect 1421 3780 1427 3782
rect 1483 3780 1507 3782
rect 1563 3780 1587 3782
rect 1643 3780 1667 3782
rect 1723 3780 1729 3782
rect 1421 3771 1729 3780
rect 1892 3292 2200 3301
rect 1892 3290 1898 3292
rect 1954 3290 1978 3292
rect 2034 3290 2058 3292
rect 2114 3290 2138 3292
rect 2194 3290 2200 3292
rect 1954 3238 1956 3290
rect 2136 3238 2138 3290
rect 1892 3236 1898 3238
rect 1954 3236 1978 3238
rect 2034 3236 2058 3238
rect 2114 3236 2138 3238
rect 2194 3236 2200 3238
rect 1892 3227 2200 3236
rect 1421 2748 1729 2757
rect 1421 2746 1427 2748
rect 1483 2746 1507 2748
rect 1563 2746 1587 2748
rect 1643 2746 1667 2748
rect 1723 2746 1729 2748
rect 1483 2694 1485 2746
rect 1665 2694 1667 2746
rect 1421 2692 1427 2694
rect 1483 2692 1507 2694
rect 1563 2692 1587 2694
rect 1643 2692 1667 2694
rect 1723 2692 1729 2694
rect 1421 2683 1729 2692
rect 1892 2204 2200 2213
rect 1892 2202 1898 2204
rect 1954 2202 1978 2204
rect 2034 2202 2058 2204
rect 2114 2202 2138 2204
rect 2194 2202 2200 2204
rect 1954 2150 1956 2202
rect 2136 2150 2138 2202
rect 1892 2148 1898 2150
rect 1954 2148 1978 2150
rect 2034 2148 2058 2150
rect 2114 2148 2138 2150
rect 2194 2148 2200 2150
rect 1892 2139 2200 2148
rect 2240 1902 2268 5086
rect 2688 5024 2740 5030
rect 2688 4966 2740 4972
rect 2364 4924 2672 4933
rect 2364 4922 2370 4924
rect 2426 4922 2450 4924
rect 2506 4922 2530 4924
rect 2586 4922 2610 4924
rect 2666 4922 2672 4924
rect 2426 4870 2428 4922
rect 2608 4870 2610 4922
rect 2364 4868 2370 4870
rect 2426 4868 2450 4870
rect 2506 4868 2530 4870
rect 2586 4868 2610 4870
rect 2666 4868 2672 4870
rect 2364 4859 2672 4868
rect 2412 4616 2464 4622
rect 2412 4558 2464 4564
rect 2424 4078 2452 4558
rect 2412 4072 2464 4078
rect 2412 4014 2464 4020
rect 2364 3836 2672 3845
rect 2364 3834 2370 3836
rect 2426 3834 2450 3836
rect 2506 3834 2530 3836
rect 2586 3834 2610 3836
rect 2666 3834 2672 3836
rect 2426 3782 2428 3834
rect 2608 3782 2610 3834
rect 2364 3780 2370 3782
rect 2426 3780 2450 3782
rect 2506 3780 2530 3782
rect 2586 3780 2610 3782
rect 2666 3780 2672 3782
rect 2364 3771 2672 3780
rect 2364 2748 2672 2757
rect 2364 2746 2370 2748
rect 2426 2746 2450 2748
rect 2506 2746 2530 2748
rect 2586 2746 2610 2748
rect 2666 2746 2672 2748
rect 2426 2694 2428 2746
rect 2608 2694 2610 2746
rect 2364 2692 2370 2694
rect 2426 2692 2450 2694
rect 2506 2692 2530 2694
rect 2586 2692 2610 2694
rect 2666 2692 2672 2694
rect 2364 2683 2672 2692
rect 2700 2417 2728 4966
rect 3160 4842 3188 5102
rect 3307 4924 3615 4933
rect 3307 4922 3313 4924
rect 3369 4922 3393 4924
rect 3449 4922 3473 4924
rect 3529 4922 3553 4924
rect 3609 4922 3615 4924
rect 3369 4870 3371 4922
rect 3551 4870 3553 4922
rect 3307 4868 3313 4870
rect 3369 4868 3393 4870
rect 3449 4868 3473 4870
rect 3529 4868 3553 4870
rect 3609 4868 3615 4870
rect 3307 4859 3615 4868
rect 3160 4814 3280 4842
rect 2835 4380 3143 4389
rect 2835 4378 2841 4380
rect 2897 4378 2921 4380
rect 2977 4378 3001 4380
rect 3057 4378 3081 4380
rect 3137 4378 3143 4380
rect 2897 4326 2899 4378
rect 3079 4326 3081 4378
rect 2835 4324 2841 4326
rect 2897 4324 2921 4326
rect 2977 4324 3001 4326
rect 3057 4324 3081 4326
rect 3137 4324 3143 4326
rect 2835 4315 3143 4324
rect 3252 4162 3280 4814
rect 3160 4134 3280 4162
rect 3160 4078 3188 4134
rect 3148 4072 3200 4078
rect 3148 4014 3200 4020
rect 3160 3754 3188 4014
rect 3307 3836 3615 3845
rect 3307 3834 3313 3836
rect 3369 3834 3393 3836
rect 3449 3834 3473 3836
rect 3529 3834 3553 3836
rect 3609 3834 3615 3836
rect 3369 3782 3371 3834
rect 3551 3782 3553 3834
rect 3307 3780 3313 3782
rect 3369 3780 3393 3782
rect 3449 3780 3473 3782
rect 3529 3780 3553 3782
rect 3609 3780 3615 3782
rect 3307 3771 3615 3780
rect 3160 3726 3280 3754
rect 2835 3292 3143 3301
rect 2835 3290 2841 3292
rect 2897 3290 2921 3292
rect 2977 3290 3001 3292
rect 3057 3290 3081 3292
rect 3137 3290 3143 3292
rect 2897 3238 2899 3290
rect 3079 3238 3081 3290
rect 2835 3236 2841 3238
rect 2897 3236 2921 3238
rect 2977 3236 3001 3238
rect 3057 3236 3081 3238
rect 3137 3236 3143 3238
rect 2835 3227 3143 3236
rect 3252 3074 3280 3726
rect 3160 3046 3280 3074
rect 3712 3058 3740 5506
rect 3778 5468 4086 5477
rect 3778 5466 3784 5468
rect 3840 5466 3864 5468
rect 3920 5466 3944 5468
rect 4000 5466 4024 5468
rect 4080 5466 4086 5468
rect 3840 5414 3842 5466
rect 4022 5414 4024 5466
rect 3778 5412 3784 5414
rect 3840 5412 3864 5414
rect 3920 5412 3944 5414
rect 4000 5412 4024 5414
rect 4080 5412 4086 5414
rect 3778 5403 4086 5412
rect 4172 4826 4200 6190
rect 4250 6012 4558 6021
rect 4250 6010 4256 6012
rect 4312 6010 4336 6012
rect 4392 6010 4416 6012
rect 4472 6010 4496 6012
rect 4552 6010 4558 6012
rect 4312 5958 4314 6010
rect 4494 5958 4496 6010
rect 4250 5956 4256 5958
rect 4312 5956 4336 5958
rect 4392 5956 4416 5958
rect 4472 5956 4496 5958
rect 4552 5956 4558 5958
rect 4250 5947 4558 5956
rect 4250 4924 4558 4933
rect 4250 4922 4256 4924
rect 4312 4922 4336 4924
rect 4392 4922 4416 4924
rect 4472 4922 4496 4924
rect 4552 4922 4558 4924
rect 4312 4870 4314 4922
rect 4494 4870 4496 4922
rect 4250 4868 4256 4870
rect 4312 4868 4336 4870
rect 4392 4868 4416 4870
rect 4472 4868 4496 4870
rect 4552 4868 4558 4870
rect 4250 4859 4558 4868
rect 4160 4820 4212 4826
rect 4160 4762 4212 4768
rect 4160 4616 4212 4622
rect 4160 4558 4212 4564
rect 3778 4380 4086 4389
rect 3778 4378 3784 4380
rect 3840 4378 3864 4380
rect 3920 4378 3944 4380
rect 4000 4378 4024 4380
rect 4080 4378 4086 4380
rect 3840 4326 3842 4378
rect 4022 4326 4024 4378
rect 3778 4324 3784 4326
rect 3840 4324 3864 4326
rect 3920 4324 3944 4326
rect 4000 4324 4024 4326
rect 4080 4324 4086 4326
rect 3778 4315 4086 4324
rect 3778 3292 4086 3301
rect 3778 3290 3784 3292
rect 3840 3290 3864 3292
rect 3920 3290 3944 3292
rect 4000 3290 4024 3292
rect 4080 3290 4086 3292
rect 3840 3238 3842 3290
rect 4022 3238 4024 3290
rect 3778 3236 3784 3238
rect 3840 3236 3864 3238
rect 3920 3236 3944 3238
rect 4000 3236 4024 3238
rect 4080 3236 4086 3238
rect 3778 3227 4086 3236
rect 3700 3052 3752 3058
rect 3160 2990 3188 3046
rect 3700 2994 3752 3000
rect 3148 2984 3200 2990
rect 3148 2926 3200 2932
rect 3160 2666 3188 2926
rect 3307 2748 3615 2757
rect 3307 2746 3313 2748
rect 3369 2746 3393 2748
rect 3449 2746 3473 2748
rect 3529 2746 3553 2748
rect 3609 2746 3615 2748
rect 3369 2694 3371 2746
rect 3551 2694 3553 2746
rect 3307 2692 3313 2694
rect 3369 2692 3393 2694
rect 3449 2692 3473 2694
rect 3529 2692 3553 2694
rect 3609 2692 3615 2694
rect 3307 2683 3615 2692
rect 3160 2638 3280 2666
rect 2686 2408 2742 2417
rect 2686 2343 2742 2352
rect 2835 2204 3143 2213
rect 2835 2202 2841 2204
rect 2897 2202 2921 2204
rect 2977 2202 3001 2204
rect 3057 2202 3081 2204
rect 3137 2202 3143 2204
rect 2897 2150 2899 2202
rect 3079 2150 3081 2202
rect 2835 2148 2841 2150
rect 2897 2148 2921 2150
rect 2977 2148 3001 2150
rect 3057 2148 3081 2150
rect 3137 2148 3143 2150
rect 2835 2139 3143 2148
rect 3252 1986 3280 2638
rect 3778 2204 4086 2213
rect 3778 2202 3784 2204
rect 3840 2202 3864 2204
rect 3920 2202 3944 2204
rect 4000 2202 4024 2204
rect 4080 2202 4086 2204
rect 3840 2150 3842 2202
rect 4022 2150 4024 2202
rect 3778 2148 3784 2150
rect 3840 2148 3864 2150
rect 3920 2148 3944 2150
rect 4000 2148 4024 2150
rect 4080 2148 4086 2150
rect 3778 2139 4086 2148
rect 4172 2038 4200 4558
rect 4250 3836 4558 3845
rect 4250 3834 4256 3836
rect 4312 3834 4336 3836
rect 4392 3834 4416 3836
rect 4472 3834 4496 3836
rect 4552 3834 4558 3836
rect 4312 3782 4314 3834
rect 4494 3782 4496 3834
rect 4250 3780 4256 3782
rect 4312 3780 4336 3782
rect 4392 3780 4416 3782
rect 4472 3780 4496 3782
rect 4552 3780 4558 3782
rect 4250 3771 4558 3780
rect 4250 2748 4558 2757
rect 4250 2746 4256 2748
rect 4312 2746 4336 2748
rect 4392 2746 4416 2748
rect 4472 2746 4496 2748
rect 4552 2746 4558 2748
rect 4312 2694 4314 2746
rect 4494 2694 4496 2746
rect 4250 2692 4256 2694
rect 4312 2692 4336 2694
rect 4392 2692 4416 2694
rect 4472 2692 4496 2694
rect 4552 2692 4558 2694
rect 4250 2683 4558 2692
rect 3160 1958 3280 1986
rect 4160 2032 4212 2038
rect 4160 1974 4212 1980
rect 1768 1896 1820 1902
rect 1768 1838 1820 1844
rect 2228 1896 2280 1902
rect 2228 1838 2280 1844
rect 1421 1660 1729 1669
rect 1421 1658 1427 1660
rect 1483 1658 1507 1660
rect 1563 1658 1587 1660
rect 1643 1658 1667 1660
rect 1723 1658 1729 1660
rect 1483 1606 1485 1658
rect 1665 1606 1667 1658
rect 1421 1604 1427 1606
rect 1483 1604 1507 1606
rect 1563 1604 1587 1606
rect 1643 1604 1667 1606
rect 1723 1604 1729 1606
rect 1421 1595 1729 1604
rect 1780 898 1808 1838
rect 2364 1660 2672 1669
rect 2364 1658 2370 1660
rect 2426 1658 2450 1660
rect 2506 1658 2530 1660
rect 2586 1658 2610 1660
rect 2666 1658 2672 1660
rect 2426 1606 2428 1658
rect 2608 1606 2610 1658
rect 2364 1604 2370 1606
rect 2426 1604 2450 1606
rect 2506 1604 2530 1606
rect 2586 1604 2610 1606
rect 2666 1604 2672 1606
rect 2364 1595 2672 1604
rect 3160 1358 3188 1958
rect 4160 1896 4212 1902
rect 4160 1838 4212 1844
rect 3307 1660 3615 1669
rect 3307 1658 3313 1660
rect 3369 1658 3393 1660
rect 3449 1658 3473 1660
rect 3529 1658 3553 1660
rect 3609 1658 3615 1660
rect 3369 1606 3371 1658
rect 3551 1606 3553 1658
rect 3307 1604 3313 1606
rect 3369 1604 3393 1606
rect 3449 1604 3473 1606
rect 3529 1604 3553 1606
rect 3609 1604 3615 1606
rect 3307 1595 3615 1604
rect 2596 1352 2648 1358
rect 2596 1294 2648 1300
rect 3148 1352 3200 1358
rect 3148 1294 3200 1300
rect 1892 1116 2200 1125
rect 1892 1114 1898 1116
rect 1954 1114 1978 1116
rect 2034 1114 2058 1116
rect 2114 1114 2138 1116
rect 2194 1114 2200 1116
rect 1954 1062 1956 1114
rect 2136 1062 2138 1114
rect 1892 1060 1898 1062
rect 1954 1060 1978 1062
rect 2034 1060 2058 1062
rect 2114 1060 2138 1062
rect 2194 1060 2200 1062
rect 1892 1051 2200 1060
rect 1780 870 1900 898
rect 1872 800 1900 870
rect 2608 800 2636 1294
rect 3332 1284 3384 1290
rect 3332 1226 3384 1232
rect 2835 1116 3143 1125
rect 2835 1114 2841 1116
rect 2897 1114 2921 1116
rect 2977 1114 3001 1116
rect 3057 1114 3081 1116
rect 3137 1114 3143 1116
rect 2897 1062 2899 1114
rect 3079 1062 3081 1114
rect 2835 1060 2841 1062
rect 2897 1060 2921 1062
rect 2977 1060 3001 1062
rect 3057 1060 3081 1062
rect 3137 1060 3143 1062
rect 2835 1051 3143 1060
rect 3344 800 3372 1226
rect 3778 1116 4086 1125
rect 3778 1114 3784 1116
rect 3840 1114 3864 1116
rect 3920 1114 3944 1116
rect 4000 1114 4024 1116
rect 4080 1114 4086 1116
rect 3840 1062 3842 1114
rect 4022 1062 4024 1114
rect 3778 1060 3784 1062
rect 3840 1060 3864 1062
rect 3920 1060 3944 1062
rect 4000 1060 4024 1062
rect 4080 1060 4086 1062
rect 3778 1051 4086 1060
rect 4172 898 4200 1838
rect 4250 1660 4558 1669
rect 4250 1658 4256 1660
rect 4312 1658 4336 1660
rect 4392 1658 4416 1660
rect 4472 1658 4496 1660
rect 4552 1658 4558 1660
rect 4312 1606 4314 1658
rect 4494 1606 4496 1658
rect 4250 1604 4256 1606
rect 4312 1604 4336 1606
rect 4392 1604 4416 1606
rect 4472 1604 4496 1606
rect 4552 1604 4558 1606
rect 4250 1595 4558 1604
rect 4080 870 4200 898
rect 4632 898 4660 6190
rect 4724 5846 4752 6310
rect 4712 5840 4764 5846
rect 4712 5782 4764 5788
rect 5092 5534 5120 8191
rect 5184 7002 5212 9415
rect 5264 8832 5316 8838
rect 5264 8774 5316 8780
rect 5172 6996 5224 7002
rect 5172 6938 5224 6944
rect 5092 5506 5212 5534
rect 4721 5468 5029 5477
rect 4721 5466 4727 5468
rect 4783 5466 4807 5468
rect 4863 5466 4887 5468
rect 4943 5466 4967 5468
rect 5023 5466 5029 5468
rect 4783 5414 4785 5466
rect 4965 5414 4967 5466
rect 4721 5412 4727 5414
rect 4783 5412 4807 5414
rect 4863 5412 4887 5414
rect 4943 5412 4967 5414
rect 5023 5412 5029 5414
rect 4721 5403 5029 5412
rect 5184 5370 5212 5506
rect 5172 5364 5224 5370
rect 5172 5306 5224 5312
rect 5078 5264 5134 5273
rect 5078 5199 5134 5208
rect 4721 4380 5029 4389
rect 4721 4378 4727 4380
rect 4783 4378 4807 4380
rect 4863 4378 4887 4380
rect 4943 4378 4967 4380
rect 5023 4378 5029 4380
rect 4783 4326 4785 4378
rect 4965 4326 4967 4378
rect 4721 4324 4727 4326
rect 4783 4324 4807 4326
rect 4863 4324 4887 4326
rect 4943 4324 4967 4326
rect 5023 4324 5029 4326
rect 4721 4315 5029 4324
rect 5092 4282 5120 5199
rect 5276 4690 5304 8774
rect 5368 7410 5396 14447
rect 5446 12472 5502 12481
rect 5446 12407 5502 12416
rect 5460 7954 5488 12407
rect 5552 10130 5580 19887
rect 5540 10124 5592 10130
rect 5540 10066 5592 10072
rect 5540 8492 5592 8498
rect 5540 8434 5592 8440
rect 5448 7948 5500 7954
rect 5448 7890 5500 7896
rect 5356 7404 5408 7410
rect 5356 7346 5408 7352
rect 5552 5534 5580 8434
rect 5460 5506 5580 5534
rect 5264 4684 5316 4690
rect 5264 4626 5316 4632
rect 5172 4480 5224 4486
rect 5172 4422 5224 4428
rect 5080 4276 5132 4282
rect 5080 4218 5132 4224
rect 5078 3768 5134 3777
rect 5184 3754 5212 4422
rect 5460 4146 5488 5506
rect 5448 4140 5500 4146
rect 5448 4082 5500 4088
rect 5134 3726 5212 3754
rect 5078 3703 5134 3712
rect 4721 3292 5029 3301
rect 4721 3290 4727 3292
rect 4783 3290 4807 3292
rect 4863 3290 4887 3292
rect 4943 3290 4967 3292
rect 5023 3290 5029 3292
rect 4783 3238 4785 3290
rect 4965 3238 4967 3290
rect 4721 3236 4727 3238
rect 4783 3236 4807 3238
rect 4863 3236 4887 3238
rect 4943 3236 4967 3238
rect 5023 3236 5029 3238
rect 4721 3227 5029 3236
rect 5080 2848 5132 2854
rect 5080 2790 5132 2796
rect 4721 2204 5029 2213
rect 4721 2202 4727 2204
rect 4783 2202 4807 2204
rect 4863 2202 4887 2204
rect 4943 2202 4967 2204
rect 5023 2202 5029 2204
rect 4783 2150 4785 2202
rect 4965 2150 4967 2202
rect 4721 2148 4727 2150
rect 4783 2148 4807 2150
rect 4863 2148 4887 2150
rect 4943 2148 4967 2150
rect 5023 2148 5029 2150
rect 4721 2139 5029 2148
rect 4721 1116 5029 1125
rect 4721 1114 4727 1116
rect 4783 1114 4807 1116
rect 4863 1114 4887 1116
rect 4943 1114 4967 1116
rect 5023 1114 5029 1116
rect 4783 1062 4785 1114
rect 4965 1062 4967 1114
rect 4721 1060 4727 1062
rect 4783 1060 4807 1062
rect 4863 1060 4887 1062
rect 4943 1060 4967 1062
rect 5023 1060 5029 1062
rect 4721 1051 5029 1060
rect 4632 870 4844 898
rect 4080 800 4108 870
rect 4816 800 4844 870
rect 386 0 442 800
rect 1122 0 1178 800
rect 1858 0 1914 800
rect 2594 0 2650 800
rect 3330 0 3386 800
rect 4066 0 4122 800
rect 4802 0 4858 800
rect 5092 785 5120 2790
rect 5540 2032 5592 2038
rect 5540 1974 5592 1980
rect 5552 800 5580 1974
rect 5078 776 5134 785
rect 5078 711 5134 720
rect 5538 0 5594 800
<< via2 >>
rect 5078 23160 5134 23216
rect 1898 22874 1954 22876
rect 1978 22874 2034 22876
rect 2058 22874 2114 22876
rect 2138 22874 2194 22876
rect 1898 22822 1944 22874
rect 1944 22822 1954 22874
rect 1978 22822 2008 22874
rect 2008 22822 2020 22874
rect 2020 22822 2034 22874
rect 2058 22822 2072 22874
rect 2072 22822 2084 22874
rect 2084 22822 2114 22874
rect 2138 22822 2148 22874
rect 2148 22822 2194 22874
rect 1898 22820 1954 22822
rect 1978 22820 2034 22822
rect 2058 22820 2114 22822
rect 2138 22820 2194 22822
rect 2841 22874 2897 22876
rect 2921 22874 2977 22876
rect 3001 22874 3057 22876
rect 3081 22874 3137 22876
rect 2841 22822 2887 22874
rect 2887 22822 2897 22874
rect 2921 22822 2951 22874
rect 2951 22822 2963 22874
rect 2963 22822 2977 22874
rect 3001 22822 3015 22874
rect 3015 22822 3027 22874
rect 3027 22822 3057 22874
rect 3081 22822 3091 22874
rect 3091 22822 3137 22874
rect 2841 22820 2897 22822
rect 2921 22820 2977 22822
rect 3001 22820 3057 22822
rect 3081 22820 3137 22822
rect 3784 22874 3840 22876
rect 3864 22874 3920 22876
rect 3944 22874 4000 22876
rect 4024 22874 4080 22876
rect 3784 22822 3830 22874
rect 3830 22822 3840 22874
rect 3864 22822 3894 22874
rect 3894 22822 3906 22874
rect 3906 22822 3920 22874
rect 3944 22822 3958 22874
rect 3958 22822 3970 22874
rect 3970 22822 4000 22874
rect 4024 22822 4034 22874
rect 4034 22822 4080 22874
rect 3784 22820 3840 22822
rect 3864 22820 3920 22822
rect 3944 22820 4000 22822
rect 4024 22820 4080 22822
rect 4727 22874 4783 22876
rect 4807 22874 4863 22876
rect 4887 22874 4943 22876
rect 4967 22874 5023 22876
rect 4727 22822 4773 22874
rect 4773 22822 4783 22874
rect 4807 22822 4837 22874
rect 4837 22822 4849 22874
rect 4849 22822 4863 22874
rect 4887 22822 4901 22874
rect 4901 22822 4913 22874
rect 4913 22822 4943 22874
rect 4967 22822 4977 22874
rect 4977 22822 5023 22874
rect 4727 22820 4783 22822
rect 4807 22820 4863 22822
rect 4887 22820 4943 22822
rect 4967 22820 5023 22822
rect 1427 22330 1483 22332
rect 1507 22330 1563 22332
rect 1587 22330 1643 22332
rect 1667 22330 1723 22332
rect 1427 22278 1473 22330
rect 1473 22278 1483 22330
rect 1507 22278 1537 22330
rect 1537 22278 1549 22330
rect 1549 22278 1563 22330
rect 1587 22278 1601 22330
rect 1601 22278 1613 22330
rect 1613 22278 1643 22330
rect 1667 22278 1677 22330
rect 1677 22278 1723 22330
rect 1427 22276 1483 22278
rect 1507 22276 1563 22278
rect 1587 22276 1643 22278
rect 1667 22276 1723 22278
rect 2370 22330 2426 22332
rect 2450 22330 2506 22332
rect 2530 22330 2586 22332
rect 2610 22330 2666 22332
rect 2370 22278 2416 22330
rect 2416 22278 2426 22330
rect 2450 22278 2480 22330
rect 2480 22278 2492 22330
rect 2492 22278 2506 22330
rect 2530 22278 2544 22330
rect 2544 22278 2556 22330
rect 2556 22278 2586 22330
rect 2610 22278 2620 22330
rect 2620 22278 2666 22330
rect 2370 22276 2426 22278
rect 2450 22276 2506 22278
rect 2530 22276 2586 22278
rect 2610 22276 2666 22278
rect 3313 22330 3369 22332
rect 3393 22330 3449 22332
rect 3473 22330 3529 22332
rect 3553 22330 3609 22332
rect 3313 22278 3359 22330
rect 3359 22278 3369 22330
rect 3393 22278 3423 22330
rect 3423 22278 3435 22330
rect 3435 22278 3449 22330
rect 3473 22278 3487 22330
rect 3487 22278 3499 22330
rect 3499 22278 3529 22330
rect 3553 22278 3563 22330
rect 3563 22278 3609 22330
rect 3313 22276 3369 22278
rect 3393 22276 3449 22278
rect 3473 22276 3529 22278
rect 3553 22276 3609 22278
rect 4256 22330 4312 22332
rect 4336 22330 4392 22332
rect 4416 22330 4472 22332
rect 4496 22330 4552 22332
rect 4256 22278 4302 22330
rect 4302 22278 4312 22330
rect 4336 22278 4366 22330
rect 4366 22278 4378 22330
rect 4378 22278 4392 22330
rect 4416 22278 4430 22330
rect 4430 22278 4442 22330
rect 4442 22278 4472 22330
rect 4496 22278 4506 22330
rect 4506 22278 4552 22330
rect 4256 22276 4312 22278
rect 4336 22276 4392 22278
rect 4416 22276 4472 22278
rect 4496 22276 4552 22278
rect 1898 21786 1954 21788
rect 1978 21786 2034 21788
rect 2058 21786 2114 21788
rect 2138 21786 2194 21788
rect 1898 21734 1944 21786
rect 1944 21734 1954 21786
rect 1978 21734 2008 21786
rect 2008 21734 2020 21786
rect 2020 21734 2034 21786
rect 2058 21734 2072 21786
rect 2072 21734 2084 21786
rect 2084 21734 2114 21786
rect 2138 21734 2148 21786
rect 2148 21734 2194 21786
rect 1898 21732 1954 21734
rect 1978 21732 2034 21734
rect 2058 21732 2114 21734
rect 2138 21732 2194 21734
rect 2841 21786 2897 21788
rect 2921 21786 2977 21788
rect 3001 21786 3057 21788
rect 3081 21786 3137 21788
rect 2841 21734 2887 21786
rect 2887 21734 2897 21786
rect 2921 21734 2951 21786
rect 2951 21734 2963 21786
rect 2963 21734 2977 21786
rect 3001 21734 3015 21786
rect 3015 21734 3027 21786
rect 3027 21734 3057 21786
rect 3081 21734 3091 21786
rect 3091 21734 3137 21786
rect 2841 21732 2897 21734
rect 2921 21732 2977 21734
rect 3001 21732 3057 21734
rect 3081 21732 3137 21734
rect 3784 21786 3840 21788
rect 3864 21786 3920 21788
rect 3944 21786 4000 21788
rect 4024 21786 4080 21788
rect 3784 21734 3830 21786
rect 3830 21734 3840 21786
rect 3864 21734 3894 21786
rect 3894 21734 3906 21786
rect 3906 21734 3920 21786
rect 3944 21734 3958 21786
rect 3958 21734 3970 21786
rect 3970 21734 4000 21786
rect 4024 21734 4034 21786
rect 4034 21734 4080 21786
rect 3784 21732 3840 21734
rect 3864 21732 3920 21734
rect 3944 21732 4000 21734
rect 4024 21732 4080 21734
rect 4727 21786 4783 21788
rect 4807 21786 4863 21788
rect 4887 21786 4943 21788
rect 4967 21786 5023 21788
rect 4727 21734 4773 21786
rect 4773 21734 4783 21786
rect 4807 21734 4837 21786
rect 4837 21734 4849 21786
rect 4849 21734 4863 21786
rect 4887 21734 4901 21786
rect 4901 21734 4913 21786
rect 4913 21734 4943 21786
rect 4967 21734 4977 21786
rect 4977 21734 5023 21786
rect 4727 21732 4783 21734
rect 4807 21732 4863 21734
rect 4887 21732 4943 21734
rect 4967 21732 5023 21734
rect 5170 21392 5226 21448
rect 1427 21242 1483 21244
rect 1507 21242 1563 21244
rect 1587 21242 1643 21244
rect 1667 21242 1723 21244
rect 1427 21190 1473 21242
rect 1473 21190 1483 21242
rect 1507 21190 1537 21242
rect 1537 21190 1549 21242
rect 1549 21190 1563 21242
rect 1587 21190 1601 21242
rect 1601 21190 1613 21242
rect 1613 21190 1643 21242
rect 1667 21190 1677 21242
rect 1677 21190 1723 21242
rect 1427 21188 1483 21190
rect 1507 21188 1563 21190
rect 1587 21188 1643 21190
rect 1667 21188 1723 21190
rect 2370 21242 2426 21244
rect 2450 21242 2506 21244
rect 2530 21242 2586 21244
rect 2610 21242 2666 21244
rect 2370 21190 2416 21242
rect 2416 21190 2426 21242
rect 2450 21190 2480 21242
rect 2480 21190 2492 21242
rect 2492 21190 2506 21242
rect 2530 21190 2544 21242
rect 2544 21190 2556 21242
rect 2556 21190 2586 21242
rect 2610 21190 2620 21242
rect 2620 21190 2666 21242
rect 2370 21188 2426 21190
rect 2450 21188 2506 21190
rect 2530 21188 2586 21190
rect 2610 21188 2666 21190
rect 3313 21242 3369 21244
rect 3393 21242 3449 21244
rect 3473 21242 3529 21244
rect 3553 21242 3609 21244
rect 3313 21190 3359 21242
rect 3359 21190 3369 21242
rect 3393 21190 3423 21242
rect 3423 21190 3435 21242
rect 3435 21190 3449 21242
rect 3473 21190 3487 21242
rect 3487 21190 3499 21242
rect 3499 21190 3529 21242
rect 3553 21190 3563 21242
rect 3563 21190 3609 21242
rect 3313 21188 3369 21190
rect 3393 21188 3449 21190
rect 3473 21188 3529 21190
rect 3553 21188 3609 21190
rect 4256 21242 4312 21244
rect 4336 21242 4392 21244
rect 4416 21242 4472 21244
rect 4496 21242 4552 21244
rect 4256 21190 4302 21242
rect 4302 21190 4312 21242
rect 4336 21190 4366 21242
rect 4366 21190 4378 21242
rect 4378 21190 4392 21242
rect 4416 21190 4430 21242
rect 4430 21190 4442 21242
rect 4442 21190 4472 21242
rect 4496 21190 4506 21242
rect 4506 21190 4552 21242
rect 4256 21188 4312 21190
rect 4336 21188 4392 21190
rect 4416 21188 4472 21190
rect 4496 21188 4552 21190
rect 1898 20698 1954 20700
rect 1978 20698 2034 20700
rect 2058 20698 2114 20700
rect 2138 20698 2194 20700
rect 1898 20646 1944 20698
rect 1944 20646 1954 20698
rect 1978 20646 2008 20698
rect 2008 20646 2020 20698
rect 2020 20646 2034 20698
rect 2058 20646 2072 20698
rect 2072 20646 2084 20698
rect 2084 20646 2114 20698
rect 2138 20646 2148 20698
rect 2148 20646 2194 20698
rect 1898 20644 1954 20646
rect 1978 20644 2034 20646
rect 2058 20644 2114 20646
rect 2138 20644 2194 20646
rect 2841 20698 2897 20700
rect 2921 20698 2977 20700
rect 3001 20698 3057 20700
rect 3081 20698 3137 20700
rect 2841 20646 2887 20698
rect 2887 20646 2897 20698
rect 2921 20646 2951 20698
rect 2951 20646 2963 20698
rect 2963 20646 2977 20698
rect 3001 20646 3015 20698
rect 3015 20646 3027 20698
rect 3027 20646 3057 20698
rect 3081 20646 3091 20698
rect 3091 20646 3137 20698
rect 2841 20644 2897 20646
rect 2921 20644 2977 20646
rect 3001 20644 3057 20646
rect 3081 20644 3137 20646
rect 3784 20698 3840 20700
rect 3864 20698 3920 20700
rect 3944 20698 4000 20700
rect 4024 20698 4080 20700
rect 3784 20646 3830 20698
rect 3830 20646 3840 20698
rect 3864 20646 3894 20698
rect 3894 20646 3906 20698
rect 3906 20646 3920 20698
rect 3944 20646 3958 20698
rect 3958 20646 3970 20698
rect 3970 20646 4000 20698
rect 4024 20646 4034 20698
rect 4034 20646 4080 20698
rect 3784 20644 3840 20646
rect 3864 20644 3920 20646
rect 3944 20644 4000 20646
rect 4024 20644 4080 20646
rect 4727 20698 4783 20700
rect 4807 20698 4863 20700
rect 4887 20698 4943 20700
rect 4967 20698 5023 20700
rect 4727 20646 4773 20698
rect 4773 20646 4783 20698
rect 4807 20646 4837 20698
rect 4837 20646 4849 20698
rect 4849 20646 4863 20698
rect 4887 20646 4901 20698
rect 4901 20646 4913 20698
rect 4913 20646 4943 20698
rect 4967 20646 4977 20698
rect 4977 20646 5023 20698
rect 4727 20644 4783 20646
rect 4807 20644 4863 20646
rect 4887 20644 4943 20646
rect 4967 20644 5023 20646
rect 1427 20154 1483 20156
rect 1507 20154 1563 20156
rect 1587 20154 1643 20156
rect 1667 20154 1723 20156
rect 1427 20102 1473 20154
rect 1473 20102 1483 20154
rect 1507 20102 1537 20154
rect 1537 20102 1549 20154
rect 1549 20102 1563 20154
rect 1587 20102 1601 20154
rect 1601 20102 1613 20154
rect 1613 20102 1643 20154
rect 1667 20102 1677 20154
rect 1677 20102 1723 20154
rect 1427 20100 1483 20102
rect 1507 20100 1563 20102
rect 1587 20100 1643 20102
rect 1667 20100 1723 20102
rect 2370 20154 2426 20156
rect 2450 20154 2506 20156
rect 2530 20154 2586 20156
rect 2610 20154 2666 20156
rect 2370 20102 2416 20154
rect 2416 20102 2426 20154
rect 2450 20102 2480 20154
rect 2480 20102 2492 20154
rect 2492 20102 2506 20154
rect 2530 20102 2544 20154
rect 2544 20102 2556 20154
rect 2556 20102 2586 20154
rect 2610 20102 2620 20154
rect 2620 20102 2666 20154
rect 2370 20100 2426 20102
rect 2450 20100 2506 20102
rect 2530 20100 2586 20102
rect 2610 20100 2666 20102
rect 3313 20154 3369 20156
rect 3393 20154 3449 20156
rect 3473 20154 3529 20156
rect 3553 20154 3609 20156
rect 3313 20102 3359 20154
rect 3359 20102 3369 20154
rect 3393 20102 3423 20154
rect 3423 20102 3435 20154
rect 3435 20102 3449 20154
rect 3473 20102 3487 20154
rect 3487 20102 3499 20154
rect 3499 20102 3529 20154
rect 3553 20102 3563 20154
rect 3563 20102 3609 20154
rect 3313 20100 3369 20102
rect 3393 20100 3449 20102
rect 3473 20100 3529 20102
rect 3553 20100 3609 20102
rect 4256 20154 4312 20156
rect 4336 20154 4392 20156
rect 4416 20154 4472 20156
rect 4496 20154 4552 20156
rect 4256 20102 4302 20154
rect 4302 20102 4312 20154
rect 4336 20102 4366 20154
rect 4366 20102 4378 20154
rect 4378 20102 4392 20154
rect 4416 20102 4430 20154
rect 4430 20102 4442 20154
rect 4442 20102 4472 20154
rect 4496 20102 4506 20154
rect 4506 20102 4552 20154
rect 4256 20100 4312 20102
rect 4336 20100 4392 20102
rect 4416 20100 4472 20102
rect 4496 20100 4552 20102
rect 1898 19610 1954 19612
rect 1978 19610 2034 19612
rect 2058 19610 2114 19612
rect 2138 19610 2194 19612
rect 1898 19558 1944 19610
rect 1944 19558 1954 19610
rect 1978 19558 2008 19610
rect 2008 19558 2020 19610
rect 2020 19558 2034 19610
rect 2058 19558 2072 19610
rect 2072 19558 2084 19610
rect 2084 19558 2114 19610
rect 2138 19558 2148 19610
rect 2148 19558 2194 19610
rect 1898 19556 1954 19558
rect 1978 19556 2034 19558
rect 2058 19556 2114 19558
rect 2138 19556 2194 19558
rect 2841 19610 2897 19612
rect 2921 19610 2977 19612
rect 3001 19610 3057 19612
rect 3081 19610 3137 19612
rect 2841 19558 2887 19610
rect 2887 19558 2897 19610
rect 2921 19558 2951 19610
rect 2951 19558 2963 19610
rect 2963 19558 2977 19610
rect 3001 19558 3015 19610
rect 3015 19558 3027 19610
rect 3027 19558 3057 19610
rect 3081 19558 3091 19610
rect 3091 19558 3137 19610
rect 2841 19556 2897 19558
rect 2921 19556 2977 19558
rect 3001 19556 3057 19558
rect 3081 19556 3137 19558
rect 3784 19610 3840 19612
rect 3864 19610 3920 19612
rect 3944 19610 4000 19612
rect 4024 19610 4080 19612
rect 3784 19558 3830 19610
rect 3830 19558 3840 19610
rect 3864 19558 3894 19610
rect 3894 19558 3906 19610
rect 3906 19558 3920 19610
rect 3944 19558 3958 19610
rect 3958 19558 3970 19610
rect 3970 19558 4000 19610
rect 4024 19558 4034 19610
rect 4034 19558 4080 19610
rect 3784 19556 3840 19558
rect 3864 19556 3920 19558
rect 3944 19556 4000 19558
rect 4024 19556 4080 19558
rect 4727 19610 4783 19612
rect 4807 19610 4863 19612
rect 4887 19610 4943 19612
rect 4967 19610 5023 19612
rect 4727 19558 4773 19610
rect 4773 19558 4783 19610
rect 4807 19558 4837 19610
rect 4837 19558 4849 19610
rect 4849 19558 4863 19610
rect 4887 19558 4901 19610
rect 4901 19558 4913 19610
rect 4913 19558 4943 19610
rect 4967 19558 4977 19610
rect 4977 19558 5023 19610
rect 4727 19556 4783 19558
rect 4807 19556 4863 19558
rect 4887 19556 4943 19558
rect 4967 19556 5023 19558
rect 1427 19066 1483 19068
rect 1507 19066 1563 19068
rect 1587 19066 1643 19068
rect 1667 19066 1723 19068
rect 1427 19014 1473 19066
rect 1473 19014 1483 19066
rect 1507 19014 1537 19066
rect 1537 19014 1549 19066
rect 1549 19014 1563 19066
rect 1587 19014 1601 19066
rect 1601 19014 1613 19066
rect 1613 19014 1643 19066
rect 1667 19014 1677 19066
rect 1677 19014 1723 19066
rect 1427 19012 1483 19014
rect 1507 19012 1563 19014
rect 1587 19012 1643 19014
rect 1667 19012 1723 19014
rect 2370 19066 2426 19068
rect 2450 19066 2506 19068
rect 2530 19066 2586 19068
rect 2610 19066 2666 19068
rect 2370 19014 2416 19066
rect 2416 19014 2426 19066
rect 2450 19014 2480 19066
rect 2480 19014 2492 19066
rect 2492 19014 2506 19066
rect 2530 19014 2544 19066
rect 2544 19014 2556 19066
rect 2556 19014 2586 19066
rect 2610 19014 2620 19066
rect 2620 19014 2666 19066
rect 2370 19012 2426 19014
rect 2450 19012 2506 19014
rect 2530 19012 2586 19014
rect 2610 19012 2666 19014
rect 3313 19066 3369 19068
rect 3393 19066 3449 19068
rect 3473 19066 3529 19068
rect 3553 19066 3609 19068
rect 3313 19014 3359 19066
rect 3359 19014 3369 19066
rect 3393 19014 3423 19066
rect 3423 19014 3435 19066
rect 3435 19014 3449 19066
rect 3473 19014 3487 19066
rect 3487 19014 3499 19066
rect 3499 19014 3529 19066
rect 3553 19014 3563 19066
rect 3563 19014 3609 19066
rect 3313 19012 3369 19014
rect 3393 19012 3449 19014
rect 3473 19012 3529 19014
rect 3553 19012 3609 19014
rect 4256 19066 4312 19068
rect 4336 19066 4392 19068
rect 4416 19066 4472 19068
rect 4496 19066 4552 19068
rect 4256 19014 4302 19066
rect 4302 19014 4312 19066
rect 4336 19014 4366 19066
rect 4366 19014 4378 19066
rect 4378 19014 4392 19066
rect 4416 19014 4430 19066
rect 4430 19014 4442 19066
rect 4442 19014 4472 19066
rect 4496 19014 4506 19066
rect 4506 19014 4552 19066
rect 4256 19012 4312 19014
rect 4336 19012 4392 19014
rect 4416 19012 4472 19014
rect 4496 19012 4552 19014
rect 4618 18672 4674 18728
rect 1898 18522 1954 18524
rect 1978 18522 2034 18524
rect 2058 18522 2114 18524
rect 2138 18522 2194 18524
rect 1898 18470 1944 18522
rect 1944 18470 1954 18522
rect 1978 18470 2008 18522
rect 2008 18470 2020 18522
rect 2020 18470 2034 18522
rect 2058 18470 2072 18522
rect 2072 18470 2084 18522
rect 2084 18470 2114 18522
rect 2138 18470 2148 18522
rect 2148 18470 2194 18522
rect 1898 18468 1954 18470
rect 1978 18468 2034 18470
rect 2058 18468 2114 18470
rect 2138 18468 2194 18470
rect 2841 18522 2897 18524
rect 2921 18522 2977 18524
rect 3001 18522 3057 18524
rect 3081 18522 3137 18524
rect 2841 18470 2887 18522
rect 2887 18470 2897 18522
rect 2921 18470 2951 18522
rect 2951 18470 2963 18522
rect 2963 18470 2977 18522
rect 3001 18470 3015 18522
rect 3015 18470 3027 18522
rect 3027 18470 3057 18522
rect 3081 18470 3091 18522
rect 3091 18470 3137 18522
rect 2841 18468 2897 18470
rect 2921 18468 2977 18470
rect 3001 18468 3057 18470
rect 3081 18468 3137 18470
rect 3784 18522 3840 18524
rect 3864 18522 3920 18524
rect 3944 18522 4000 18524
rect 4024 18522 4080 18524
rect 3784 18470 3830 18522
rect 3830 18470 3840 18522
rect 3864 18470 3894 18522
rect 3894 18470 3906 18522
rect 3906 18470 3920 18522
rect 3944 18470 3958 18522
rect 3958 18470 3970 18522
rect 3970 18470 4000 18522
rect 4024 18470 4034 18522
rect 4034 18470 4080 18522
rect 3784 18468 3840 18470
rect 3864 18468 3920 18470
rect 3944 18468 4000 18470
rect 4024 18468 4080 18470
rect 1427 17978 1483 17980
rect 1507 17978 1563 17980
rect 1587 17978 1643 17980
rect 1667 17978 1723 17980
rect 1427 17926 1473 17978
rect 1473 17926 1483 17978
rect 1507 17926 1537 17978
rect 1537 17926 1549 17978
rect 1549 17926 1563 17978
rect 1587 17926 1601 17978
rect 1601 17926 1613 17978
rect 1613 17926 1643 17978
rect 1667 17926 1677 17978
rect 1677 17926 1723 17978
rect 1427 17924 1483 17926
rect 1507 17924 1563 17926
rect 1587 17924 1643 17926
rect 1667 17924 1723 17926
rect 2370 17978 2426 17980
rect 2450 17978 2506 17980
rect 2530 17978 2586 17980
rect 2610 17978 2666 17980
rect 2370 17926 2416 17978
rect 2416 17926 2426 17978
rect 2450 17926 2480 17978
rect 2480 17926 2492 17978
rect 2492 17926 2506 17978
rect 2530 17926 2544 17978
rect 2544 17926 2556 17978
rect 2556 17926 2586 17978
rect 2610 17926 2620 17978
rect 2620 17926 2666 17978
rect 2370 17924 2426 17926
rect 2450 17924 2506 17926
rect 2530 17924 2586 17926
rect 2610 17924 2666 17926
rect 3313 17978 3369 17980
rect 3393 17978 3449 17980
rect 3473 17978 3529 17980
rect 3553 17978 3609 17980
rect 3313 17926 3359 17978
rect 3359 17926 3369 17978
rect 3393 17926 3423 17978
rect 3423 17926 3435 17978
rect 3435 17926 3449 17978
rect 3473 17926 3487 17978
rect 3487 17926 3499 17978
rect 3499 17926 3529 17978
rect 3553 17926 3563 17978
rect 3563 17926 3609 17978
rect 3313 17924 3369 17926
rect 3393 17924 3449 17926
rect 3473 17924 3529 17926
rect 3553 17924 3609 17926
rect 4256 17978 4312 17980
rect 4336 17978 4392 17980
rect 4416 17978 4472 17980
rect 4496 17978 4552 17980
rect 4256 17926 4302 17978
rect 4302 17926 4312 17978
rect 4336 17926 4366 17978
rect 4366 17926 4378 17978
rect 4378 17926 4392 17978
rect 4416 17926 4430 17978
rect 4430 17926 4442 17978
rect 4442 17926 4472 17978
rect 4496 17926 4506 17978
rect 4506 17926 4552 17978
rect 4256 17924 4312 17926
rect 4336 17924 4392 17926
rect 4416 17924 4472 17926
rect 4496 17924 4552 17926
rect 1898 17434 1954 17436
rect 1978 17434 2034 17436
rect 2058 17434 2114 17436
rect 2138 17434 2194 17436
rect 1898 17382 1944 17434
rect 1944 17382 1954 17434
rect 1978 17382 2008 17434
rect 2008 17382 2020 17434
rect 2020 17382 2034 17434
rect 2058 17382 2072 17434
rect 2072 17382 2084 17434
rect 2084 17382 2114 17434
rect 2138 17382 2148 17434
rect 2148 17382 2194 17434
rect 1898 17380 1954 17382
rect 1978 17380 2034 17382
rect 2058 17380 2114 17382
rect 2138 17380 2194 17382
rect 2841 17434 2897 17436
rect 2921 17434 2977 17436
rect 3001 17434 3057 17436
rect 3081 17434 3137 17436
rect 2841 17382 2887 17434
rect 2887 17382 2897 17434
rect 2921 17382 2951 17434
rect 2951 17382 2963 17434
rect 2963 17382 2977 17434
rect 3001 17382 3015 17434
rect 3015 17382 3027 17434
rect 3027 17382 3057 17434
rect 3081 17382 3091 17434
rect 3091 17382 3137 17434
rect 2841 17380 2897 17382
rect 2921 17380 2977 17382
rect 3001 17380 3057 17382
rect 3081 17380 3137 17382
rect 3784 17434 3840 17436
rect 3864 17434 3920 17436
rect 3944 17434 4000 17436
rect 4024 17434 4080 17436
rect 3784 17382 3830 17434
rect 3830 17382 3840 17434
rect 3864 17382 3894 17434
rect 3894 17382 3906 17434
rect 3906 17382 3920 17434
rect 3944 17382 3958 17434
rect 3958 17382 3970 17434
rect 3970 17382 4000 17434
rect 4024 17382 4034 17434
rect 4034 17382 4080 17434
rect 3784 17380 3840 17382
rect 3864 17380 3920 17382
rect 3944 17380 4000 17382
rect 4024 17380 4080 17382
rect 1427 16890 1483 16892
rect 1507 16890 1563 16892
rect 1587 16890 1643 16892
rect 1667 16890 1723 16892
rect 1427 16838 1473 16890
rect 1473 16838 1483 16890
rect 1507 16838 1537 16890
rect 1537 16838 1549 16890
rect 1549 16838 1563 16890
rect 1587 16838 1601 16890
rect 1601 16838 1613 16890
rect 1613 16838 1643 16890
rect 1667 16838 1677 16890
rect 1677 16838 1723 16890
rect 1427 16836 1483 16838
rect 1507 16836 1563 16838
rect 1587 16836 1643 16838
rect 1667 16836 1723 16838
rect 2370 16890 2426 16892
rect 2450 16890 2506 16892
rect 2530 16890 2586 16892
rect 2610 16890 2666 16892
rect 2370 16838 2416 16890
rect 2416 16838 2426 16890
rect 2450 16838 2480 16890
rect 2480 16838 2492 16890
rect 2492 16838 2506 16890
rect 2530 16838 2544 16890
rect 2544 16838 2556 16890
rect 2556 16838 2586 16890
rect 2610 16838 2620 16890
rect 2620 16838 2666 16890
rect 2370 16836 2426 16838
rect 2450 16836 2506 16838
rect 2530 16836 2586 16838
rect 2610 16836 2666 16838
rect 3313 16890 3369 16892
rect 3393 16890 3449 16892
rect 3473 16890 3529 16892
rect 3553 16890 3609 16892
rect 3313 16838 3359 16890
rect 3359 16838 3369 16890
rect 3393 16838 3423 16890
rect 3423 16838 3435 16890
rect 3435 16838 3449 16890
rect 3473 16838 3487 16890
rect 3487 16838 3499 16890
rect 3499 16838 3529 16890
rect 3553 16838 3563 16890
rect 3563 16838 3609 16890
rect 3313 16836 3369 16838
rect 3393 16836 3449 16838
rect 3473 16836 3529 16838
rect 3553 16836 3609 16838
rect 4256 16890 4312 16892
rect 4336 16890 4392 16892
rect 4416 16890 4472 16892
rect 4496 16890 4552 16892
rect 4256 16838 4302 16890
rect 4302 16838 4312 16890
rect 4336 16838 4366 16890
rect 4366 16838 4378 16890
rect 4378 16838 4392 16890
rect 4416 16838 4430 16890
rect 4430 16838 4442 16890
rect 4442 16838 4472 16890
rect 4496 16838 4506 16890
rect 4506 16838 4552 16890
rect 4256 16836 4312 16838
rect 4336 16836 4392 16838
rect 4416 16836 4472 16838
rect 4496 16836 4552 16838
rect 1898 16346 1954 16348
rect 1978 16346 2034 16348
rect 2058 16346 2114 16348
rect 2138 16346 2194 16348
rect 1898 16294 1944 16346
rect 1944 16294 1954 16346
rect 1978 16294 2008 16346
rect 2008 16294 2020 16346
rect 2020 16294 2034 16346
rect 2058 16294 2072 16346
rect 2072 16294 2084 16346
rect 2084 16294 2114 16346
rect 2138 16294 2148 16346
rect 2148 16294 2194 16346
rect 1898 16292 1954 16294
rect 1978 16292 2034 16294
rect 2058 16292 2114 16294
rect 2138 16292 2194 16294
rect 2841 16346 2897 16348
rect 2921 16346 2977 16348
rect 3001 16346 3057 16348
rect 3081 16346 3137 16348
rect 2841 16294 2887 16346
rect 2887 16294 2897 16346
rect 2921 16294 2951 16346
rect 2951 16294 2963 16346
rect 2963 16294 2977 16346
rect 3001 16294 3015 16346
rect 3015 16294 3027 16346
rect 3027 16294 3057 16346
rect 3081 16294 3091 16346
rect 3091 16294 3137 16346
rect 2841 16292 2897 16294
rect 2921 16292 2977 16294
rect 3001 16292 3057 16294
rect 3081 16292 3137 16294
rect 3784 16346 3840 16348
rect 3864 16346 3920 16348
rect 3944 16346 4000 16348
rect 4024 16346 4080 16348
rect 3784 16294 3830 16346
rect 3830 16294 3840 16346
rect 3864 16294 3894 16346
rect 3894 16294 3906 16346
rect 3906 16294 3920 16346
rect 3944 16294 3958 16346
rect 3958 16294 3970 16346
rect 3970 16294 4000 16346
rect 4024 16294 4034 16346
rect 4034 16294 4080 16346
rect 3784 16292 3840 16294
rect 3864 16292 3920 16294
rect 3944 16292 4000 16294
rect 4024 16292 4080 16294
rect 1427 15802 1483 15804
rect 1507 15802 1563 15804
rect 1587 15802 1643 15804
rect 1667 15802 1723 15804
rect 1427 15750 1473 15802
rect 1473 15750 1483 15802
rect 1507 15750 1537 15802
rect 1537 15750 1549 15802
rect 1549 15750 1563 15802
rect 1587 15750 1601 15802
rect 1601 15750 1613 15802
rect 1613 15750 1643 15802
rect 1667 15750 1677 15802
rect 1677 15750 1723 15802
rect 1427 15748 1483 15750
rect 1507 15748 1563 15750
rect 1587 15748 1643 15750
rect 1667 15748 1723 15750
rect 2370 15802 2426 15804
rect 2450 15802 2506 15804
rect 2530 15802 2586 15804
rect 2610 15802 2666 15804
rect 2370 15750 2416 15802
rect 2416 15750 2426 15802
rect 2450 15750 2480 15802
rect 2480 15750 2492 15802
rect 2492 15750 2506 15802
rect 2530 15750 2544 15802
rect 2544 15750 2556 15802
rect 2556 15750 2586 15802
rect 2610 15750 2620 15802
rect 2620 15750 2666 15802
rect 2370 15748 2426 15750
rect 2450 15748 2506 15750
rect 2530 15748 2586 15750
rect 2610 15748 2666 15750
rect 3313 15802 3369 15804
rect 3393 15802 3449 15804
rect 3473 15802 3529 15804
rect 3553 15802 3609 15804
rect 3313 15750 3359 15802
rect 3359 15750 3369 15802
rect 3393 15750 3423 15802
rect 3423 15750 3435 15802
rect 3435 15750 3449 15802
rect 3473 15750 3487 15802
rect 3487 15750 3499 15802
rect 3499 15750 3529 15802
rect 3553 15750 3563 15802
rect 3563 15750 3609 15802
rect 3313 15748 3369 15750
rect 3393 15748 3449 15750
rect 3473 15748 3529 15750
rect 3553 15748 3609 15750
rect 4256 15802 4312 15804
rect 4336 15802 4392 15804
rect 4416 15802 4472 15804
rect 4496 15802 4552 15804
rect 4256 15750 4302 15802
rect 4302 15750 4312 15802
rect 4336 15750 4366 15802
rect 4366 15750 4378 15802
rect 4378 15750 4392 15802
rect 4416 15750 4430 15802
rect 4430 15750 4442 15802
rect 4442 15750 4472 15802
rect 4496 15750 4506 15802
rect 4506 15750 4552 15802
rect 4256 15748 4312 15750
rect 4336 15748 4392 15750
rect 4416 15748 4472 15750
rect 4496 15748 4552 15750
rect 3698 15544 3754 15600
rect 1898 15258 1954 15260
rect 1978 15258 2034 15260
rect 2058 15258 2114 15260
rect 2138 15258 2194 15260
rect 1898 15206 1944 15258
rect 1944 15206 1954 15258
rect 1978 15206 2008 15258
rect 2008 15206 2020 15258
rect 2020 15206 2034 15258
rect 2058 15206 2072 15258
rect 2072 15206 2084 15258
rect 2084 15206 2114 15258
rect 2138 15206 2148 15258
rect 2148 15206 2194 15258
rect 1898 15204 1954 15206
rect 1978 15204 2034 15206
rect 2058 15204 2114 15206
rect 2138 15204 2194 15206
rect 2841 15258 2897 15260
rect 2921 15258 2977 15260
rect 3001 15258 3057 15260
rect 3081 15258 3137 15260
rect 2841 15206 2887 15258
rect 2887 15206 2897 15258
rect 2921 15206 2951 15258
rect 2951 15206 2963 15258
rect 2963 15206 2977 15258
rect 3001 15206 3015 15258
rect 3015 15206 3027 15258
rect 3027 15206 3057 15258
rect 3081 15206 3091 15258
rect 3091 15206 3137 15258
rect 2841 15204 2897 15206
rect 2921 15204 2977 15206
rect 3001 15204 3057 15206
rect 3081 15204 3137 15206
rect 1427 14714 1483 14716
rect 1507 14714 1563 14716
rect 1587 14714 1643 14716
rect 1667 14714 1723 14716
rect 1427 14662 1473 14714
rect 1473 14662 1483 14714
rect 1507 14662 1537 14714
rect 1537 14662 1549 14714
rect 1549 14662 1563 14714
rect 1587 14662 1601 14714
rect 1601 14662 1613 14714
rect 1613 14662 1643 14714
rect 1667 14662 1677 14714
rect 1677 14662 1723 14714
rect 1427 14660 1483 14662
rect 1507 14660 1563 14662
rect 1587 14660 1643 14662
rect 1667 14660 1723 14662
rect 2370 14714 2426 14716
rect 2450 14714 2506 14716
rect 2530 14714 2586 14716
rect 2610 14714 2666 14716
rect 2370 14662 2416 14714
rect 2416 14662 2426 14714
rect 2450 14662 2480 14714
rect 2480 14662 2492 14714
rect 2492 14662 2506 14714
rect 2530 14662 2544 14714
rect 2544 14662 2556 14714
rect 2556 14662 2586 14714
rect 2610 14662 2620 14714
rect 2620 14662 2666 14714
rect 2370 14660 2426 14662
rect 2450 14660 2506 14662
rect 2530 14660 2586 14662
rect 2610 14660 2666 14662
rect 3313 14714 3369 14716
rect 3393 14714 3449 14716
rect 3473 14714 3529 14716
rect 3553 14714 3609 14716
rect 3313 14662 3359 14714
rect 3359 14662 3369 14714
rect 3393 14662 3423 14714
rect 3423 14662 3435 14714
rect 3435 14662 3449 14714
rect 3473 14662 3487 14714
rect 3487 14662 3499 14714
rect 3499 14662 3529 14714
rect 3553 14662 3563 14714
rect 3563 14662 3609 14714
rect 3313 14660 3369 14662
rect 3393 14660 3449 14662
rect 3473 14660 3529 14662
rect 3553 14660 3609 14662
rect 1898 14170 1954 14172
rect 1978 14170 2034 14172
rect 2058 14170 2114 14172
rect 2138 14170 2194 14172
rect 1898 14118 1944 14170
rect 1944 14118 1954 14170
rect 1978 14118 2008 14170
rect 2008 14118 2020 14170
rect 2020 14118 2034 14170
rect 2058 14118 2072 14170
rect 2072 14118 2084 14170
rect 2084 14118 2114 14170
rect 2138 14118 2148 14170
rect 2148 14118 2194 14170
rect 1898 14116 1954 14118
rect 1978 14116 2034 14118
rect 2058 14116 2114 14118
rect 2138 14116 2194 14118
rect 2841 14170 2897 14172
rect 2921 14170 2977 14172
rect 3001 14170 3057 14172
rect 3081 14170 3137 14172
rect 2841 14118 2887 14170
rect 2887 14118 2897 14170
rect 2921 14118 2951 14170
rect 2951 14118 2963 14170
rect 2963 14118 2977 14170
rect 3001 14118 3015 14170
rect 3015 14118 3027 14170
rect 3027 14118 3057 14170
rect 3081 14118 3091 14170
rect 3091 14118 3137 14170
rect 2841 14116 2897 14118
rect 2921 14116 2977 14118
rect 3001 14116 3057 14118
rect 3081 14116 3137 14118
rect 1427 13626 1483 13628
rect 1507 13626 1563 13628
rect 1587 13626 1643 13628
rect 1667 13626 1723 13628
rect 1427 13574 1473 13626
rect 1473 13574 1483 13626
rect 1507 13574 1537 13626
rect 1537 13574 1549 13626
rect 1549 13574 1563 13626
rect 1587 13574 1601 13626
rect 1601 13574 1613 13626
rect 1613 13574 1643 13626
rect 1667 13574 1677 13626
rect 1677 13574 1723 13626
rect 1427 13572 1483 13574
rect 1507 13572 1563 13574
rect 1587 13572 1643 13574
rect 1667 13572 1723 13574
rect 2370 13626 2426 13628
rect 2450 13626 2506 13628
rect 2530 13626 2586 13628
rect 2610 13626 2666 13628
rect 2370 13574 2416 13626
rect 2416 13574 2426 13626
rect 2450 13574 2480 13626
rect 2480 13574 2492 13626
rect 2492 13574 2506 13626
rect 2530 13574 2544 13626
rect 2544 13574 2556 13626
rect 2556 13574 2586 13626
rect 2610 13574 2620 13626
rect 2620 13574 2666 13626
rect 2370 13572 2426 13574
rect 2450 13572 2506 13574
rect 2530 13572 2586 13574
rect 2610 13572 2666 13574
rect 3313 13626 3369 13628
rect 3393 13626 3449 13628
rect 3473 13626 3529 13628
rect 3553 13626 3609 13628
rect 3313 13574 3359 13626
rect 3359 13574 3369 13626
rect 3393 13574 3423 13626
rect 3423 13574 3435 13626
rect 3435 13574 3449 13626
rect 3473 13574 3487 13626
rect 3487 13574 3499 13626
rect 3499 13574 3529 13626
rect 3553 13574 3563 13626
rect 3563 13574 3609 13626
rect 3313 13572 3369 13574
rect 3393 13572 3449 13574
rect 3473 13572 3529 13574
rect 3553 13572 3609 13574
rect 1898 13082 1954 13084
rect 1978 13082 2034 13084
rect 2058 13082 2114 13084
rect 2138 13082 2194 13084
rect 1898 13030 1944 13082
rect 1944 13030 1954 13082
rect 1978 13030 2008 13082
rect 2008 13030 2020 13082
rect 2020 13030 2034 13082
rect 2058 13030 2072 13082
rect 2072 13030 2084 13082
rect 2084 13030 2114 13082
rect 2138 13030 2148 13082
rect 2148 13030 2194 13082
rect 1898 13028 1954 13030
rect 1978 13028 2034 13030
rect 2058 13028 2114 13030
rect 2138 13028 2194 13030
rect 2841 13082 2897 13084
rect 2921 13082 2977 13084
rect 3001 13082 3057 13084
rect 3081 13082 3137 13084
rect 2841 13030 2887 13082
rect 2887 13030 2897 13082
rect 2921 13030 2951 13082
rect 2951 13030 2963 13082
rect 2963 13030 2977 13082
rect 3001 13030 3015 13082
rect 3015 13030 3027 13082
rect 3027 13030 3057 13082
rect 3081 13030 3091 13082
rect 3091 13030 3137 13082
rect 2841 13028 2897 13030
rect 2921 13028 2977 13030
rect 3001 13028 3057 13030
rect 3081 13028 3137 13030
rect 1427 12538 1483 12540
rect 1507 12538 1563 12540
rect 1587 12538 1643 12540
rect 1667 12538 1723 12540
rect 1427 12486 1473 12538
rect 1473 12486 1483 12538
rect 1507 12486 1537 12538
rect 1537 12486 1549 12538
rect 1549 12486 1563 12538
rect 1587 12486 1601 12538
rect 1601 12486 1613 12538
rect 1613 12486 1643 12538
rect 1667 12486 1677 12538
rect 1677 12486 1723 12538
rect 1427 12484 1483 12486
rect 1507 12484 1563 12486
rect 1587 12484 1643 12486
rect 1667 12484 1723 12486
rect 2370 12538 2426 12540
rect 2450 12538 2506 12540
rect 2530 12538 2586 12540
rect 2610 12538 2666 12540
rect 2370 12486 2416 12538
rect 2416 12486 2426 12538
rect 2450 12486 2480 12538
rect 2480 12486 2492 12538
rect 2492 12486 2506 12538
rect 2530 12486 2544 12538
rect 2544 12486 2556 12538
rect 2556 12486 2586 12538
rect 2610 12486 2620 12538
rect 2620 12486 2666 12538
rect 2370 12484 2426 12486
rect 2450 12484 2506 12486
rect 2530 12484 2586 12486
rect 2610 12484 2666 12486
rect 3313 12538 3369 12540
rect 3393 12538 3449 12540
rect 3473 12538 3529 12540
rect 3553 12538 3609 12540
rect 3313 12486 3359 12538
rect 3359 12486 3369 12538
rect 3393 12486 3423 12538
rect 3423 12486 3435 12538
rect 3435 12486 3449 12538
rect 3473 12486 3487 12538
rect 3487 12486 3499 12538
rect 3499 12486 3529 12538
rect 3553 12486 3563 12538
rect 3563 12486 3609 12538
rect 3313 12484 3369 12486
rect 3393 12484 3449 12486
rect 3473 12484 3529 12486
rect 3553 12484 3609 12486
rect 1898 11994 1954 11996
rect 1978 11994 2034 11996
rect 2058 11994 2114 11996
rect 2138 11994 2194 11996
rect 1898 11942 1944 11994
rect 1944 11942 1954 11994
rect 1978 11942 2008 11994
rect 2008 11942 2020 11994
rect 2020 11942 2034 11994
rect 2058 11942 2072 11994
rect 2072 11942 2084 11994
rect 2084 11942 2114 11994
rect 2138 11942 2148 11994
rect 2148 11942 2194 11994
rect 1898 11940 1954 11942
rect 1978 11940 2034 11942
rect 2058 11940 2114 11942
rect 2138 11940 2194 11942
rect 2841 11994 2897 11996
rect 2921 11994 2977 11996
rect 3001 11994 3057 11996
rect 3081 11994 3137 11996
rect 2841 11942 2887 11994
rect 2887 11942 2897 11994
rect 2921 11942 2951 11994
rect 2951 11942 2963 11994
rect 2963 11942 2977 11994
rect 3001 11942 3015 11994
rect 3015 11942 3027 11994
rect 3027 11942 3057 11994
rect 3081 11942 3091 11994
rect 3091 11942 3137 11994
rect 2841 11940 2897 11942
rect 2921 11940 2977 11942
rect 3001 11940 3057 11942
rect 3081 11940 3137 11942
rect 1427 11450 1483 11452
rect 1507 11450 1563 11452
rect 1587 11450 1643 11452
rect 1667 11450 1723 11452
rect 1427 11398 1473 11450
rect 1473 11398 1483 11450
rect 1507 11398 1537 11450
rect 1537 11398 1549 11450
rect 1549 11398 1563 11450
rect 1587 11398 1601 11450
rect 1601 11398 1613 11450
rect 1613 11398 1643 11450
rect 1667 11398 1677 11450
rect 1677 11398 1723 11450
rect 1427 11396 1483 11398
rect 1507 11396 1563 11398
rect 1587 11396 1643 11398
rect 1667 11396 1723 11398
rect 1427 10362 1483 10364
rect 1507 10362 1563 10364
rect 1587 10362 1643 10364
rect 1667 10362 1723 10364
rect 1427 10310 1473 10362
rect 1473 10310 1483 10362
rect 1507 10310 1537 10362
rect 1537 10310 1549 10362
rect 1549 10310 1563 10362
rect 1587 10310 1601 10362
rect 1601 10310 1613 10362
rect 1613 10310 1643 10362
rect 1667 10310 1677 10362
rect 1677 10310 1723 10362
rect 1427 10308 1483 10310
rect 1507 10308 1563 10310
rect 1587 10308 1643 10310
rect 1667 10308 1723 10310
rect 1427 9274 1483 9276
rect 1507 9274 1563 9276
rect 1587 9274 1643 9276
rect 1667 9274 1723 9276
rect 1427 9222 1473 9274
rect 1473 9222 1483 9274
rect 1507 9222 1537 9274
rect 1537 9222 1549 9274
rect 1549 9222 1563 9274
rect 1587 9222 1601 9274
rect 1601 9222 1613 9274
rect 1613 9222 1643 9274
rect 1667 9222 1677 9274
rect 1677 9222 1723 9274
rect 1427 9220 1483 9222
rect 1507 9220 1563 9222
rect 1587 9220 1643 9222
rect 1667 9220 1723 9222
rect 2370 11450 2426 11452
rect 2450 11450 2506 11452
rect 2530 11450 2586 11452
rect 2610 11450 2666 11452
rect 2370 11398 2416 11450
rect 2416 11398 2426 11450
rect 2450 11398 2480 11450
rect 2480 11398 2492 11450
rect 2492 11398 2506 11450
rect 2530 11398 2544 11450
rect 2544 11398 2556 11450
rect 2556 11398 2586 11450
rect 2610 11398 2620 11450
rect 2620 11398 2666 11450
rect 2370 11396 2426 11398
rect 2450 11396 2506 11398
rect 2530 11396 2586 11398
rect 2610 11396 2666 11398
rect 3313 11450 3369 11452
rect 3393 11450 3449 11452
rect 3473 11450 3529 11452
rect 3553 11450 3609 11452
rect 3313 11398 3359 11450
rect 3359 11398 3369 11450
rect 3393 11398 3423 11450
rect 3423 11398 3435 11450
rect 3435 11398 3449 11450
rect 3473 11398 3487 11450
rect 3487 11398 3499 11450
rect 3499 11398 3529 11450
rect 3553 11398 3563 11450
rect 3563 11398 3609 11450
rect 3313 11396 3369 11398
rect 3393 11396 3449 11398
rect 3473 11396 3529 11398
rect 3553 11396 3609 11398
rect 1898 10906 1954 10908
rect 1978 10906 2034 10908
rect 2058 10906 2114 10908
rect 2138 10906 2194 10908
rect 1898 10854 1944 10906
rect 1944 10854 1954 10906
rect 1978 10854 2008 10906
rect 2008 10854 2020 10906
rect 2020 10854 2034 10906
rect 2058 10854 2072 10906
rect 2072 10854 2084 10906
rect 2084 10854 2114 10906
rect 2138 10854 2148 10906
rect 2148 10854 2194 10906
rect 1898 10852 1954 10854
rect 1978 10852 2034 10854
rect 2058 10852 2114 10854
rect 2138 10852 2194 10854
rect 2370 10362 2426 10364
rect 2450 10362 2506 10364
rect 2530 10362 2586 10364
rect 2610 10362 2666 10364
rect 2370 10310 2416 10362
rect 2416 10310 2426 10362
rect 2450 10310 2480 10362
rect 2480 10310 2492 10362
rect 2492 10310 2506 10362
rect 2530 10310 2544 10362
rect 2544 10310 2556 10362
rect 2556 10310 2586 10362
rect 2610 10310 2620 10362
rect 2620 10310 2666 10362
rect 2370 10308 2426 10310
rect 2450 10308 2506 10310
rect 2530 10308 2586 10310
rect 2610 10308 2666 10310
rect 1898 9818 1954 9820
rect 1978 9818 2034 9820
rect 2058 9818 2114 9820
rect 2138 9818 2194 9820
rect 1898 9766 1944 9818
rect 1944 9766 1954 9818
rect 1978 9766 2008 9818
rect 2008 9766 2020 9818
rect 2020 9766 2034 9818
rect 2058 9766 2072 9818
rect 2072 9766 2084 9818
rect 2084 9766 2114 9818
rect 2138 9766 2148 9818
rect 2148 9766 2194 9818
rect 1898 9764 1954 9766
rect 1978 9764 2034 9766
rect 2058 9764 2114 9766
rect 2138 9764 2194 9766
rect 1427 8186 1483 8188
rect 1507 8186 1563 8188
rect 1587 8186 1643 8188
rect 1667 8186 1723 8188
rect 1427 8134 1473 8186
rect 1473 8134 1483 8186
rect 1507 8134 1537 8186
rect 1537 8134 1549 8186
rect 1549 8134 1563 8186
rect 1587 8134 1601 8186
rect 1601 8134 1613 8186
rect 1613 8134 1643 8186
rect 1667 8134 1677 8186
rect 1677 8134 1723 8186
rect 1427 8132 1483 8134
rect 1507 8132 1563 8134
rect 1587 8132 1643 8134
rect 1667 8132 1723 8134
rect 1898 8730 1954 8732
rect 1978 8730 2034 8732
rect 2058 8730 2114 8732
rect 2138 8730 2194 8732
rect 1898 8678 1944 8730
rect 1944 8678 1954 8730
rect 1978 8678 2008 8730
rect 2008 8678 2020 8730
rect 2020 8678 2034 8730
rect 2058 8678 2072 8730
rect 2072 8678 2084 8730
rect 2084 8678 2114 8730
rect 2138 8678 2148 8730
rect 2148 8678 2194 8730
rect 1898 8676 1954 8678
rect 1978 8676 2034 8678
rect 2058 8676 2114 8678
rect 2138 8676 2194 8678
rect 2841 10906 2897 10908
rect 2921 10906 2977 10908
rect 3001 10906 3057 10908
rect 3081 10906 3137 10908
rect 2841 10854 2887 10906
rect 2887 10854 2897 10906
rect 2921 10854 2951 10906
rect 2951 10854 2963 10906
rect 2963 10854 2977 10906
rect 3001 10854 3015 10906
rect 3015 10854 3027 10906
rect 3027 10854 3057 10906
rect 3081 10854 3091 10906
rect 3091 10854 3137 10906
rect 2841 10852 2897 10854
rect 2921 10852 2977 10854
rect 3001 10852 3057 10854
rect 3081 10852 3137 10854
rect 3422 11228 3424 11248
rect 3424 11228 3476 11248
rect 3476 11228 3478 11248
rect 3422 11192 3478 11228
rect 3313 10362 3369 10364
rect 3393 10362 3449 10364
rect 3473 10362 3529 10364
rect 3553 10362 3609 10364
rect 3313 10310 3359 10362
rect 3359 10310 3369 10362
rect 3393 10310 3423 10362
rect 3423 10310 3435 10362
rect 3435 10310 3449 10362
rect 3473 10310 3487 10362
rect 3487 10310 3499 10362
rect 3499 10310 3529 10362
rect 3553 10310 3563 10362
rect 3563 10310 3609 10362
rect 3313 10308 3369 10310
rect 3393 10308 3449 10310
rect 3473 10308 3529 10310
rect 3553 10308 3609 10310
rect 2841 9818 2897 9820
rect 2921 9818 2977 9820
rect 3001 9818 3057 9820
rect 3081 9818 3137 9820
rect 2841 9766 2887 9818
rect 2887 9766 2897 9818
rect 2921 9766 2951 9818
rect 2951 9766 2963 9818
rect 2963 9766 2977 9818
rect 3001 9766 3015 9818
rect 3015 9766 3027 9818
rect 3027 9766 3057 9818
rect 3081 9766 3091 9818
rect 3091 9766 3137 9818
rect 2841 9764 2897 9766
rect 2921 9764 2977 9766
rect 3001 9764 3057 9766
rect 3081 9764 3137 9766
rect 2370 9274 2426 9276
rect 2450 9274 2506 9276
rect 2530 9274 2586 9276
rect 2610 9274 2666 9276
rect 2370 9222 2416 9274
rect 2416 9222 2426 9274
rect 2450 9222 2480 9274
rect 2480 9222 2492 9274
rect 2492 9222 2506 9274
rect 2530 9222 2544 9274
rect 2544 9222 2556 9274
rect 2556 9222 2586 9274
rect 2610 9222 2620 9274
rect 2620 9222 2666 9274
rect 2370 9220 2426 9222
rect 2450 9220 2506 9222
rect 2530 9220 2586 9222
rect 2610 9220 2666 9222
rect 2370 8186 2426 8188
rect 2450 8186 2506 8188
rect 2530 8186 2586 8188
rect 2610 8186 2666 8188
rect 2370 8134 2416 8186
rect 2416 8134 2426 8186
rect 2450 8134 2480 8186
rect 2480 8134 2492 8186
rect 2492 8134 2506 8186
rect 2530 8134 2544 8186
rect 2544 8134 2556 8186
rect 2556 8134 2586 8186
rect 2610 8134 2620 8186
rect 2620 8134 2666 8186
rect 2370 8132 2426 8134
rect 2450 8132 2506 8134
rect 2530 8132 2586 8134
rect 2610 8132 2666 8134
rect 1898 7642 1954 7644
rect 1978 7642 2034 7644
rect 2058 7642 2114 7644
rect 2138 7642 2194 7644
rect 1898 7590 1944 7642
rect 1944 7590 1954 7642
rect 1978 7590 2008 7642
rect 2008 7590 2020 7642
rect 2020 7590 2034 7642
rect 2058 7590 2072 7642
rect 2072 7590 2084 7642
rect 2084 7590 2114 7642
rect 2138 7590 2148 7642
rect 2148 7590 2194 7642
rect 1898 7588 1954 7590
rect 1978 7588 2034 7590
rect 2058 7588 2114 7590
rect 2138 7588 2194 7590
rect 1427 7098 1483 7100
rect 1507 7098 1563 7100
rect 1587 7098 1643 7100
rect 1667 7098 1723 7100
rect 1427 7046 1473 7098
rect 1473 7046 1483 7098
rect 1507 7046 1537 7098
rect 1537 7046 1549 7098
rect 1549 7046 1563 7098
rect 1587 7046 1601 7098
rect 1601 7046 1613 7098
rect 1613 7046 1643 7098
rect 1667 7046 1677 7098
rect 1677 7046 1723 7098
rect 1427 7044 1483 7046
rect 1507 7044 1563 7046
rect 1587 7044 1643 7046
rect 1667 7044 1723 7046
rect 1898 6554 1954 6556
rect 1978 6554 2034 6556
rect 2058 6554 2114 6556
rect 2138 6554 2194 6556
rect 1898 6502 1944 6554
rect 1944 6502 1954 6554
rect 1978 6502 2008 6554
rect 2008 6502 2020 6554
rect 2020 6502 2034 6554
rect 2058 6502 2072 6554
rect 2072 6502 2084 6554
rect 2084 6502 2114 6554
rect 2138 6502 2148 6554
rect 2148 6502 2194 6554
rect 1898 6500 1954 6502
rect 1978 6500 2034 6502
rect 2058 6500 2114 6502
rect 2138 6500 2194 6502
rect 2370 7098 2426 7100
rect 2450 7098 2506 7100
rect 2530 7098 2586 7100
rect 2610 7098 2666 7100
rect 2370 7046 2416 7098
rect 2416 7046 2426 7098
rect 2450 7046 2480 7098
rect 2480 7046 2492 7098
rect 2492 7046 2506 7098
rect 2530 7046 2544 7098
rect 2544 7046 2556 7098
rect 2556 7046 2586 7098
rect 2610 7046 2620 7098
rect 2620 7046 2666 7098
rect 2370 7044 2426 7046
rect 2450 7044 2506 7046
rect 2530 7044 2586 7046
rect 2610 7044 2666 7046
rect 3313 9274 3369 9276
rect 3393 9274 3449 9276
rect 3473 9274 3529 9276
rect 3553 9274 3609 9276
rect 3313 9222 3359 9274
rect 3359 9222 3369 9274
rect 3393 9222 3423 9274
rect 3423 9222 3435 9274
rect 3435 9222 3449 9274
rect 3473 9222 3487 9274
rect 3487 9222 3499 9274
rect 3499 9222 3529 9274
rect 3553 9222 3563 9274
rect 3563 9222 3609 9274
rect 3313 9220 3369 9222
rect 3393 9220 3449 9222
rect 3473 9220 3529 9222
rect 3553 9220 3609 9222
rect 2841 8730 2897 8732
rect 2921 8730 2977 8732
rect 3001 8730 3057 8732
rect 3081 8730 3137 8732
rect 2841 8678 2887 8730
rect 2887 8678 2897 8730
rect 2921 8678 2951 8730
rect 2951 8678 2963 8730
rect 2963 8678 2977 8730
rect 3001 8678 3015 8730
rect 3015 8678 3027 8730
rect 3027 8678 3057 8730
rect 3081 8678 3091 8730
rect 3091 8678 3137 8730
rect 2841 8676 2897 8678
rect 2921 8676 2977 8678
rect 3001 8676 3057 8678
rect 3081 8676 3137 8678
rect 3784 15258 3840 15260
rect 3864 15258 3920 15260
rect 3944 15258 4000 15260
rect 4024 15258 4080 15260
rect 3784 15206 3830 15258
rect 3830 15206 3840 15258
rect 3864 15206 3894 15258
rect 3894 15206 3906 15258
rect 3906 15206 3920 15258
rect 3944 15206 3958 15258
rect 3958 15206 3970 15258
rect 3970 15206 4000 15258
rect 4024 15206 4034 15258
rect 4034 15206 4080 15258
rect 3784 15204 3840 15206
rect 3864 15204 3920 15206
rect 3944 15204 4000 15206
rect 4024 15204 4080 15206
rect 4256 14714 4312 14716
rect 4336 14714 4392 14716
rect 4416 14714 4472 14716
rect 4496 14714 4552 14716
rect 4256 14662 4302 14714
rect 4302 14662 4312 14714
rect 4336 14662 4366 14714
rect 4366 14662 4378 14714
rect 4378 14662 4392 14714
rect 4416 14662 4430 14714
rect 4430 14662 4442 14714
rect 4442 14662 4472 14714
rect 4496 14662 4506 14714
rect 4506 14662 4552 14714
rect 4256 14660 4312 14662
rect 4336 14660 4392 14662
rect 4416 14660 4472 14662
rect 4496 14660 4552 14662
rect 3784 14170 3840 14172
rect 3864 14170 3920 14172
rect 3944 14170 4000 14172
rect 4024 14170 4080 14172
rect 3784 14118 3830 14170
rect 3830 14118 3840 14170
rect 3864 14118 3894 14170
rect 3894 14118 3906 14170
rect 3906 14118 3920 14170
rect 3944 14118 3958 14170
rect 3958 14118 3970 14170
rect 3970 14118 4000 14170
rect 4024 14118 4034 14170
rect 4034 14118 4080 14170
rect 3784 14116 3840 14118
rect 3864 14116 3920 14118
rect 3944 14116 4000 14118
rect 4024 14116 4080 14118
rect 4256 13626 4312 13628
rect 4336 13626 4392 13628
rect 4416 13626 4472 13628
rect 4496 13626 4552 13628
rect 4256 13574 4302 13626
rect 4302 13574 4312 13626
rect 4336 13574 4366 13626
rect 4366 13574 4378 13626
rect 4378 13574 4392 13626
rect 4416 13574 4430 13626
rect 4430 13574 4442 13626
rect 4442 13574 4472 13626
rect 4496 13574 4506 13626
rect 4506 13574 4552 13626
rect 4256 13572 4312 13574
rect 4336 13572 4392 13574
rect 4416 13572 4472 13574
rect 4496 13572 4552 13574
rect 3784 13082 3840 13084
rect 3864 13082 3920 13084
rect 3944 13082 4000 13084
rect 4024 13082 4080 13084
rect 3784 13030 3830 13082
rect 3830 13030 3840 13082
rect 3864 13030 3894 13082
rect 3894 13030 3906 13082
rect 3906 13030 3920 13082
rect 3944 13030 3958 13082
rect 3958 13030 3970 13082
rect 3970 13030 4000 13082
rect 4024 13030 4034 13082
rect 4034 13030 4080 13082
rect 3784 13028 3840 13030
rect 3864 13028 3920 13030
rect 3944 13028 4000 13030
rect 4024 13028 4080 13030
rect 4256 12538 4312 12540
rect 4336 12538 4392 12540
rect 4416 12538 4472 12540
rect 4496 12538 4552 12540
rect 4256 12486 4302 12538
rect 4302 12486 4312 12538
rect 4336 12486 4366 12538
rect 4366 12486 4378 12538
rect 4378 12486 4392 12538
rect 4416 12486 4430 12538
rect 4430 12486 4442 12538
rect 4442 12486 4472 12538
rect 4496 12486 4506 12538
rect 4506 12486 4552 12538
rect 4256 12484 4312 12486
rect 4336 12484 4392 12486
rect 4416 12484 4472 12486
rect 4496 12484 4552 12486
rect 3784 11994 3840 11996
rect 3864 11994 3920 11996
rect 3944 11994 4000 11996
rect 4024 11994 4080 11996
rect 3784 11942 3830 11994
rect 3830 11942 3840 11994
rect 3864 11942 3894 11994
rect 3894 11942 3906 11994
rect 3906 11942 3920 11994
rect 3944 11942 3958 11994
rect 3958 11942 3970 11994
rect 3970 11942 4000 11994
rect 4024 11942 4034 11994
rect 4034 11942 4080 11994
rect 3784 11940 3840 11942
rect 3864 11940 3920 11942
rect 3944 11940 4000 11942
rect 4024 11940 4080 11942
rect 3784 10906 3840 10908
rect 3864 10906 3920 10908
rect 3944 10906 4000 10908
rect 4024 10906 4080 10908
rect 3784 10854 3830 10906
rect 3830 10854 3840 10906
rect 3864 10854 3894 10906
rect 3894 10854 3906 10906
rect 3906 10854 3920 10906
rect 3944 10854 3958 10906
rect 3958 10854 3970 10906
rect 3970 10854 4000 10906
rect 4024 10854 4034 10906
rect 4034 10854 4080 10906
rect 3784 10852 3840 10854
rect 3864 10852 3920 10854
rect 3944 10852 4000 10854
rect 4024 10852 4080 10854
rect 4256 11450 4312 11452
rect 4336 11450 4392 11452
rect 4416 11450 4472 11452
rect 4496 11450 4552 11452
rect 4256 11398 4302 11450
rect 4302 11398 4312 11450
rect 4336 11398 4366 11450
rect 4366 11398 4378 11450
rect 4378 11398 4392 11450
rect 4416 11398 4430 11450
rect 4430 11398 4442 11450
rect 4442 11398 4472 11450
rect 4496 11398 4506 11450
rect 4506 11398 4552 11450
rect 4256 11396 4312 11398
rect 4336 11396 4392 11398
rect 4416 11396 4472 11398
rect 4496 11396 4552 11398
rect 3784 9818 3840 9820
rect 3864 9818 3920 9820
rect 3944 9818 4000 9820
rect 4024 9818 4080 9820
rect 3784 9766 3830 9818
rect 3830 9766 3840 9818
rect 3864 9766 3894 9818
rect 3894 9766 3906 9818
rect 3906 9766 3920 9818
rect 3944 9766 3958 9818
rect 3958 9766 3970 9818
rect 3970 9766 4000 9818
rect 4024 9766 4034 9818
rect 4034 9766 4080 9818
rect 3784 9764 3840 9766
rect 3864 9764 3920 9766
rect 3944 9764 4000 9766
rect 4024 9764 4080 9766
rect 4256 10362 4312 10364
rect 4336 10362 4392 10364
rect 4416 10362 4472 10364
rect 4496 10362 4552 10364
rect 4256 10310 4302 10362
rect 4302 10310 4312 10362
rect 4336 10310 4366 10362
rect 4366 10310 4378 10362
rect 4378 10310 4392 10362
rect 4416 10310 4430 10362
rect 4430 10310 4442 10362
rect 4442 10310 4472 10362
rect 4496 10310 4506 10362
rect 4506 10310 4552 10362
rect 4256 10308 4312 10310
rect 4336 10308 4392 10310
rect 4416 10308 4472 10310
rect 4496 10308 4552 10310
rect 4727 18522 4783 18524
rect 4807 18522 4863 18524
rect 4887 18522 4943 18524
rect 4967 18522 5023 18524
rect 4727 18470 4773 18522
rect 4773 18470 4783 18522
rect 4807 18470 4837 18522
rect 4837 18470 4849 18522
rect 4849 18470 4863 18522
rect 4887 18470 4901 18522
rect 4901 18470 4913 18522
rect 4913 18470 4943 18522
rect 4967 18470 4977 18522
rect 4977 18470 5023 18522
rect 4727 18468 4783 18470
rect 4807 18468 4863 18470
rect 4887 18468 4943 18470
rect 4967 18468 5023 18470
rect 4727 17434 4783 17436
rect 4807 17434 4863 17436
rect 4887 17434 4943 17436
rect 4967 17434 5023 17436
rect 4727 17382 4773 17434
rect 4773 17382 4783 17434
rect 4807 17382 4837 17434
rect 4837 17382 4849 17434
rect 4849 17382 4863 17434
rect 4887 17382 4901 17434
rect 4901 17382 4913 17434
rect 4913 17382 4943 17434
rect 4967 17382 4977 17434
rect 4977 17382 5023 17434
rect 4727 17380 4783 17382
rect 4807 17380 4863 17382
rect 4887 17380 4943 17382
rect 4967 17380 5023 17382
rect 5078 17176 5134 17232
rect 4727 16346 4783 16348
rect 4807 16346 4863 16348
rect 4887 16346 4943 16348
rect 4967 16346 5023 16348
rect 4727 16294 4773 16346
rect 4773 16294 4783 16346
rect 4807 16294 4837 16346
rect 4837 16294 4849 16346
rect 4849 16294 4863 16346
rect 4887 16294 4901 16346
rect 4901 16294 4913 16346
rect 4913 16294 4943 16346
rect 4967 16294 4977 16346
rect 4977 16294 5023 16346
rect 4727 16292 4783 16294
rect 4807 16292 4863 16294
rect 4887 16292 4943 16294
rect 4967 16292 5023 16294
rect 4727 15258 4783 15260
rect 4807 15258 4863 15260
rect 4887 15258 4943 15260
rect 4967 15258 5023 15260
rect 4727 15206 4773 15258
rect 4773 15206 4783 15258
rect 4807 15206 4837 15258
rect 4837 15206 4849 15258
rect 4849 15206 4863 15258
rect 4887 15206 4901 15258
rect 4901 15206 4913 15258
rect 4913 15206 4943 15258
rect 4967 15206 4977 15258
rect 4977 15206 5023 15258
rect 4727 15204 4783 15206
rect 4807 15204 4863 15206
rect 4887 15204 4943 15206
rect 4967 15204 5023 15206
rect 4727 14170 4783 14172
rect 4807 14170 4863 14172
rect 4887 14170 4943 14172
rect 4967 14170 5023 14172
rect 4727 14118 4773 14170
rect 4773 14118 4783 14170
rect 4807 14118 4837 14170
rect 4837 14118 4849 14170
rect 4849 14118 4863 14170
rect 4887 14118 4901 14170
rect 4901 14118 4913 14170
rect 4913 14118 4943 14170
rect 4967 14118 4977 14170
rect 4977 14118 5023 14170
rect 4727 14116 4783 14118
rect 4807 14116 4863 14118
rect 4887 14116 4943 14118
rect 4967 14116 5023 14118
rect 4727 13082 4783 13084
rect 4807 13082 4863 13084
rect 4887 13082 4943 13084
rect 4967 13082 5023 13084
rect 4727 13030 4773 13082
rect 4773 13030 4783 13082
rect 4807 13030 4837 13082
rect 4837 13030 4849 13082
rect 4849 13030 4863 13082
rect 4887 13030 4901 13082
rect 4901 13030 4913 13082
rect 4913 13030 4943 13082
rect 4967 13030 4977 13082
rect 4977 13030 5023 13082
rect 4727 13028 4783 13030
rect 4807 13028 4863 13030
rect 4887 13028 4943 13030
rect 4967 13028 5023 13030
rect 4727 11994 4783 11996
rect 4807 11994 4863 11996
rect 4887 11994 4943 11996
rect 4967 11994 5023 11996
rect 4727 11942 4773 11994
rect 4773 11942 4783 11994
rect 4807 11942 4837 11994
rect 4837 11942 4849 11994
rect 4849 11942 4863 11994
rect 4887 11942 4901 11994
rect 4901 11942 4913 11994
rect 4913 11942 4943 11994
rect 4967 11942 4977 11994
rect 4977 11942 5023 11994
rect 4727 11940 4783 11942
rect 4807 11940 4863 11942
rect 4887 11940 4943 11942
rect 4967 11940 5023 11942
rect 4727 10906 4783 10908
rect 4807 10906 4863 10908
rect 4887 10906 4943 10908
rect 4967 10906 5023 10908
rect 4727 10854 4773 10906
rect 4773 10854 4783 10906
rect 4807 10854 4837 10906
rect 4837 10854 4849 10906
rect 4849 10854 4863 10906
rect 4887 10854 4901 10906
rect 4901 10854 4913 10906
rect 4913 10854 4943 10906
rect 4967 10854 4977 10906
rect 4977 10854 5023 10906
rect 4727 10852 4783 10854
rect 4807 10852 4863 10854
rect 4887 10852 4943 10854
rect 4967 10852 5023 10854
rect 3784 8730 3840 8732
rect 3864 8730 3920 8732
rect 3944 8730 4000 8732
rect 4024 8730 4080 8732
rect 3784 8678 3830 8730
rect 3830 8678 3840 8730
rect 3864 8678 3894 8730
rect 3894 8678 3906 8730
rect 3906 8678 3920 8730
rect 3944 8678 3958 8730
rect 3958 8678 3970 8730
rect 3970 8678 4000 8730
rect 4024 8678 4034 8730
rect 4034 8678 4080 8730
rect 3784 8676 3840 8678
rect 3864 8676 3920 8678
rect 3944 8676 4000 8678
rect 4024 8676 4080 8678
rect 4256 9274 4312 9276
rect 4336 9274 4392 9276
rect 4416 9274 4472 9276
rect 4496 9274 4552 9276
rect 4256 9222 4302 9274
rect 4302 9222 4312 9274
rect 4336 9222 4366 9274
rect 4366 9222 4378 9274
rect 4378 9222 4392 9274
rect 4416 9222 4430 9274
rect 4430 9222 4442 9274
rect 4442 9222 4472 9274
rect 4496 9222 4506 9274
rect 4506 9222 4552 9274
rect 4256 9220 4312 9222
rect 4336 9220 4392 9222
rect 4416 9220 4472 9222
rect 4496 9220 4552 9222
rect 3313 8186 3369 8188
rect 3393 8186 3449 8188
rect 3473 8186 3529 8188
rect 3553 8186 3609 8188
rect 3313 8134 3359 8186
rect 3359 8134 3369 8186
rect 3393 8134 3423 8186
rect 3423 8134 3435 8186
rect 3435 8134 3449 8186
rect 3473 8134 3487 8186
rect 3487 8134 3499 8186
rect 3499 8134 3529 8186
rect 3553 8134 3563 8186
rect 3563 8134 3609 8186
rect 3313 8132 3369 8134
rect 3393 8132 3449 8134
rect 3473 8132 3529 8134
rect 3553 8132 3609 8134
rect 2841 7642 2897 7644
rect 2921 7642 2977 7644
rect 3001 7642 3057 7644
rect 3081 7642 3137 7644
rect 2841 7590 2887 7642
rect 2887 7590 2897 7642
rect 2921 7590 2951 7642
rect 2951 7590 2963 7642
rect 2963 7590 2977 7642
rect 3001 7590 3015 7642
rect 3015 7590 3027 7642
rect 3027 7590 3057 7642
rect 3081 7590 3091 7642
rect 3091 7590 3137 7642
rect 2841 7588 2897 7590
rect 2921 7588 2977 7590
rect 3001 7588 3057 7590
rect 3081 7588 3137 7590
rect 3784 7642 3840 7644
rect 3864 7642 3920 7644
rect 3944 7642 4000 7644
rect 4024 7642 4080 7644
rect 3784 7590 3830 7642
rect 3830 7590 3840 7642
rect 3864 7590 3894 7642
rect 3894 7590 3906 7642
rect 3906 7590 3920 7642
rect 3944 7590 3958 7642
rect 3958 7590 3970 7642
rect 3970 7590 4000 7642
rect 4024 7590 4034 7642
rect 4034 7590 4080 7642
rect 3784 7588 3840 7590
rect 3864 7588 3920 7590
rect 3944 7588 4000 7590
rect 4024 7588 4080 7590
rect 4256 8186 4312 8188
rect 4336 8186 4392 8188
rect 4416 8186 4472 8188
rect 4496 8186 4552 8188
rect 4256 8134 4302 8186
rect 4302 8134 4312 8186
rect 4336 8134 4366 8186
rect 4366 8134 4378 8186
rect 4378 8134 4392 8186
rect 4416 8134 4430 8186
rect 4430 8134 4442 8186
rect 4442 8134 4472 8186
rect 4496 8134 4506 8186
rect 4506 8134 4552 8186
rect 4256 8132 4312 8134
rect 4336 8132 4392 8134
rect 4416 8132 4472 8134
rect 4496 8132 4552 8134
rect 3313 7098 3369 7100
rect 3393 7098 3449 7100
rect 3473 7098 3529 7100
rect 3553 7098 3609 7100
rect 3313 7046 3359 7098
rect 3359 7046 3369 7098
rect 3393 7046 3423 7098
rect 3423 7046 3435 7098
rect 3435 7046 3449 7098
rect 3473 7046 3487 7098
rect 3487 7046 3499 7098
rect 3499 7046 3529 7098
rect 3553 7046 3563 7098
rect 3563 7046 3609 7098
rect 3313 7044 3369 7046
rect 3393 7044 3449 7046
rect 3473 7044 3529 7046
rect 3553 7044 3609 7046
rect 2841 6554 2897 6556
rect 2921 6554 2977 6556
rect 3001 6554 3057 6556
rect 3081 6554 3137 6556
rect 2841 6502 2887 6554
rect 2887 6502 2897 6554
rect 2921 6502 2951 6554
rect 2951 6502 2963 6554
rect 2963 6502 2977 6554
rect 3001 6502 3015 6554
rect 3015 6502 3027 6554
rect 3027 6502 3057 6554
rect 3081 6502 3091 6554
rect 3091 6502 3137 6554
rect 2841 6500 2897 6502
rect 2921 6500 2977 6502
rect 3001 6500 3057 6502
rect 3081 6500 3137 6502
rect 3606 6704 3662 6760
rect 3514 6296 3570 6352
rect 3784 6554 3840 6556
rect 3864 6554 3920 6556
rect 3944 6554 4000 6556
rect 4024 6554 4080 6556
rect 3784 6502 3830 6554
rect 3830 6502 3840 6554
rect 3864 6502 3894 6554
rect 3894 6502 3906 6554
rect 3906 6502 3920 6554
rect 3944 6502 3958 6554
rect 3958 6502 3970 6554
rect 3970 6502 4000 6554
rect 4024 6502 4034 6554
rect 4034 6502 4080 6554
rect 3784 6500 3840 6502
rect 3864 6500 3920 6502
rect 3944 6500 4000 6502
rect 4024 6500 4080 6502
rect 3790 6296 3846 6352
rect 1427 6010 1483 6012
rect 1507 6010 1563 6012
rect 1587 6010 1643 6012
rect 1667 6010 1723 6012
rect 1427 5958 1473 6010
rect 1473 5958 1483 6010
rect 1507 5958 1537 6010
rect 1537 5958 1549 6010
rect 1549 5958 1563 6010
rect 1587 5958 1601 6010
rect 1601 5958 1613 6010
rect 1613 5958 1643 6010
rect 1667 5958 1677 6010
rect 1677 5958 1723 6010
rect 1427 5956 1483 5958
rect 1507 5956 1563 5958
rect 1587 5956 1643 5958
rect 1667 5956 1723 5958
rect 1898 5466 1954 5468
rect 1978 5466 2034 5468
rect 2058 5466 2114 5468
rect 2138 5466 2194 5468
rect 1898 5414 1944 5466
rect 1944 5414 1954 5466
rect 1978 5414 2008 5466
rect 2008 5414 2020 5466
rect 2020 5414 2034 5466
rect 2058 5414 2072 5466
rect 2072 5414 2084 5466
rect 2084 5414 2114 5466
rect 2138 5414 2148 5466
rect 2148 5414 2194 5466
rect 1898 5412 1954 5414
rect 1978 5412 2034 5414
rect 2058 5412 2114 5414
rect 2138 5412 2194 5414
rect 2370 6010 2426 6012
rect 2450 6010 2506 6012
rect 2530 6010 2586 6012
rect 2610 6010 2666 6012
rect 2370 5958 2416 6010
rect 2416 5958 2426 6010
rect 2450 5958 2480 6010
rect 2480 5958 2492 6010
rect 2492 5958 2506 6010
rect 2530 5958 2544 6010
rect 2544 5958 2556 6010
rect 2556 5958 2586 6010
rect 2610 5958 2620 6010
rect 2620 5958 2666 6010
rect 2370 5956 2426 5958
rect 2450 5956 2506 5958
rect 2530 5956 2586 5958
rect 2610 5956 2666 5958
rect 3313 6010 3369 6012
rect 3393 6010 3449 6012
rect 3473 6010 3529 6012
rect 3553 6010 3609 6012
rect 3313 5958 3359 6010
rect 3359 5958 3369 6010
rect 3393 5958 3423 6010
rect 3423 5958 3435 6010
rect 3435 5958 3449 6010
rect 3473 5958 3487 6010
rect 3487 5958 3499 6010
rect 3499 5958 3529 6010
rect 3553 5958 3563 6010
rect 3563 5958 3609 6010
rect 3313 5956 3369 5958
rect 3393 5956 3449 5958
rect 3473 5956 3529 5958
rect 3553 5956 3609 5958
rect 2841 5466 2897 5468
rect 2921 5466 2977 5468
rect 3001 5466 3057 5468
rect 3081 5466 3137 5468
rect 2841 5414 2887 5466
rect 2887 5414 2897 5466
rect 2921 5414 2951 5466
rect 2951 5414 2963 5466
rect 2963 5414 2977 5466
rect 3001 5414 3015 5466
rect 3015 5414 3027 5466
rect 3027 5414 3057 5466
rect 3081 5414 3091 5466
rect 3091 5414 3137 5466
rect 2841 5412 2897 5414
rect 2921 5412 2977 5414
rect 3001 5412 3057 5414
rect 3081 5412 3137 5414
rect 4256 7098 4312 7100
rect 4336 7098 4392 7100
rect 4416 7098 4472 7100
rect 4496 7098 4552 7100
rect 4256 7046 4302 7098
rect 4302 7046 4312 7098
rect 4336 7046 4366 7098
rect 4366 7046 4378 7098
rect 4378 7046 4392 7098
rect 4416 7046 4430 7098
rect 4430 7046 4442 7098
rect 4442 7046 4472 7098
rect 4496 7046 4506 7098
rect 4506 7046 4552 7098
rect 4256 7044 4312 7046
rect 4336 7044 4392 7046
rect 4416 7044 4472 7046
rect 4496 7044 4552 7046
rect 4727 9818 4783 9820
rect 4807 9818 4863 9820
rect 4887 9818 4943 9820
rect 4967 9818 5023 9820
rect 4727 9766 4773 9818
rect 4773 9766 4783 9818
rect 4807 9766 4837 9818
rect 4837 9766 4849 9818
rect 4849 9766 4863 9818
rect 4887 9766 4901 9818
rect 4901 9766 4913 9818
rect 4913 9766 4943 9818
rect 4967 9766 4977 9818
rect 4977 9766 5023 9818
rect 4727 9764 4783 9766
rect 4807 9764 4863 9766
rect 4887 9764 4943 9766
rect 4967 9764 5023 9766
rect 5538 19896 5594 19952
rect 5354 14456 5410 14512
rect 5170 9424 5226 9480
rect 4727 8730 4783 8732
rect 4807 8730 4863 8732
rect 4887 8730 4943 8732
rect 4967 8730 5023 8732
rect 4727 8678 4773 8730
rect 4773 8678 4783 8730
rect 4807 8678 4837 8730
rect 4837 8678 4849 8730
rect 4849 8678 4863 8730
rect 4887 8678 4901 8730
rect 4901 8678 4913 8730
rect 4913 8678 4943 8730
rect 4967 8678 4977 8730
rect 4977 8678 5023 8730
rect 4727 8676 4783 8678
rect 4807 8676 4863 8678
rect 4887 8676 4943 8678
rect 4967 8676 5023 8678
rect 5078 8200 5134 8256
rect 4727 7642 4783 7644
rect 4807 7642 4863 7644
rect 4887 7642 4943 7644
rect 4967 7642 5023 7644
rect 4727 7590 4773 7642
rect 4773 7590 4783 7642
rect 4807 7590 4837 7642
rect 4837 7590 4849 7642
rect 4849 7590 4863 7642
rect 4887 7590 4901 7642
rect 4901 7590 4913 7642
rect 4913 7590 4943 7642
rect 4967 7590 4977 7642
rect 4977 7590 5023 7642
rect 4727 7588 4783 7590
rect 4807 7588 4863 7590
rect 4887 7588 4943 7590
rect 4967 7588 5023 7590
rect 4727 6554 4783 6556
rect 4807 6554 4863 6556
rect 4887 6554 4943 6556
rect 4967 6554 5023 6556
rect 4727 6502 4773 6554
rect 4773 6502 4783 6554
rect 4807 6502 4837 6554
rect 4837 6502 4849 6554
rect 4849 6502 4863 6554
rect 4887 6502 4901 6554
rect 4901 6502 4913 6554
rect 4913 6502 4943 6554
rect 4967 6502 4977 6554
rect 4977 6502 5023 6554
rect 4727 6500 4783 6502
rect 4807 6500 4863 6502
rect 4887 6500 4943 6502
rect 4967 6500 5023 6502
rect 1427 4922 1483 4924
rect 1507 4922 1563 4924
rect 1587 4922 1643 4924
rect 1667 4922 1723 4924
rect 1427 4870 1473 4922
rect 1473 4870 1483 4922
rect 1507 4870 1537 4922
rect 1537 4870 1549 4922
rect 1549 4870 1563 4922
rect 1587 4870 1601 4922
rect 1601 4870 1613 4922
rect 1613 4870 1643 4922
rect 1667 4870 1677 4922
rect 1677 4870 1723 4922
rect 1427 4868 1483 4870
rect 1507 4868 1563 4870
rect 1587 4868 1643 4870
rect 1667 4868 1723 4870
rect 1898 4378 1954 4380
rect 1978 4378 2034 4380
rect 2058 4378 2114 4380
rect 2138 4378 2194 4380
rect 1898 4326 1944 4378
rect 1944 4326 1954 4378
rect 1978 4326 2008 4378
rect 2008 4326 2020 4378
rect 2020 4326 2034 4378
rect 2058 4326 2072 4378
rect 2072 4326 2084 4378
rect 2084 4326 2114 4378
rect 2138 4326 2148 4378
rect 2148 4326 2194 4378
rect 1898 4324 1954 4326
rect 1978 4324 2034 4326
rect 2058 4324 2114 4326
rect 2138 4324 2194 4326
rect 1427 3834 1483 3836
rect 1507 3834 1563 3836
rect 1587 3834 1643 3836
rect 1667 3834 1723 3836
rect 1427 3782 1473 3834
rect 1473 3782 1483 3834
rect 1507 3782 1537 3834
rect 1537 3782 1549 3834
rect 1549 3782 1563 3834
rect 1587 3782 1601 3834
rect 1601 3782 1613 3834
rect 1613 3782 1643 3834
rect 1667 3782 1677 3834
rect 1677 3782 1723 3834
rect 1427 3780 1483 3782
rect 1507 3780 1563 3782
rect 1587 3780 1643 3782
rect 1667 3780 1723 3782
rect 1898 3290 1954 3292
rect 1978 3290 2034 3292
rect 2058 3290 2114 3292
rect 2138 3290 2194 3292
rect 1898 3238 1944 3290
rect 1944 3238 1954 3290
rect 1978 3238 2008 3290
rect 2008 3238 2020 3290
rect 2020 3238 2034 3290
rect 2058 3238 2072 3290
rect 2072 3238 2084 3290
rect 2084 3238 2114 3290
rect 2138 3238 2148 3290
rect 2148 3238 2194 3290
rect 1898 3236 1954 3238
rect 1978 3236 2034 3238
rect 2058 3236 2114 3238
rect 2138 3236 2194 3238
rect 1427 2746 1483 2748
rect 1507 2746 1563 2748
rect 1587 2746 1643 2748
rect 1667 2746 1723 2748
rect 1427 2694 1473 2746
rect 1473 2694 1483 2746
rect 1507 2694 1537 2746
rect 1537 2694 1549 2746
rect 1549 2694 1563 2746
rect 1587 2694 1601 2746
rect 1601 2694 1613 2746
rect 1613 2694 1643 2746
rect 1667 2694 1677 2746
rect 1677 2694 1723 2746
rect 1427 2692 1483 2694
rect 1507 2692 1563 2694
rect 1587 2692 1643 2694
rect 1667 2692 1723 2694
rect 1898 2202 1954 2204
rect 1978 2202 2034 2204
rect 2058 2202 2114 2204
rect 2138 2202 2194 2204
rect 1898 2150 1944 2202
rect 1944 2150 1954 2202
rect 1978 2150 2008 2202
rect 2008 2150 2020 2202
rect 2020 2150 2034 2202
rect 2058 2150 2072 2202
rect 2072 2150 2084 2202
rect 2084 2150 2114 2202
rect 2138 2150 2148 2202
rect 2148 2150 2194 2202
rect 1898 2148 1954 2150
rect 1978 2148 2034 2150
rect 2058 2148 2114 2150
rect 2138 2148 2194 2150
rect 2370 4922 2426 4924
rect 2450 4922 2506 4924
rect 2530 4922 2586 4924
rect 2610 4922 2666 4924
rect 2370 4870 2416 4922
rect 2416 4870 2426 4922
rect 2450 4870 2480 4922
rect 2480 4870 2492 4922
rect 2492 4870 2506 4922
rect 2530 4870 2544 4922
rect 2544 4870 2556 4922
rect 2556 4870 2586 4922
rect 2610 4870 2620 4922
rect 2620 4870 2666 4922
rect 2370 4868 2426 4870
rect 2450 4868 2506 4870
rect 2530 4868 2586 4870
rect 2610 4868 2666 4870
rect 2370 3834 2426 3836
rect 2450 3834 2506 3836
rect 2530 3834 2586 3836
rect 2610 3834 2666 3836
rect 2370 3782 2416 3834
rect 2416 3782 2426 3834
rect 2450 3782 2480 3834
rect 2480 3782 2492 3834
rect 2492 3782 2506 3834
rect 2530 3782 2544 3834
rect 2544 3782 2556 3834
rect 2556 3782 2586 3834
rect 2610 3782 2620 3834
rect 2620 3782 2666 3834
rect 2370 3780 2426 3782
rect 2450 3780 2506 3782
rect 2530 3780 2586 3782
rect 2610 3780 2666 3782
rect 2370 2746 2426 2748
rect 2450 2746 2506 2748
rect 2530 2746 2586 2748
rect 2610 2746 2666 2748
rect 2370 2694 2416 2746
rect 2416 2694 2426 2746
rect 2450 2694 2480 2746
rect 2480 2694 2492 2746
rect 2492 2694 2506 2746
rect 2530 2694 2544 2746
rect 2544 2694 2556 2746
rect 2556 2694 2586 2746
rect 2610 2694 2620 2746
rect 2620 2694 2666 2746
rect 2370 2692 2426 2694
rect 2450 2692 2506 2694
rect 2530 2692 2586 2694
rect 2610 2692 2666 2694
rect 3313 4922 3369 4924
rect 3393 4922 3449 4924
rect 3473 4922 3529 4924
rect 3553 4922 3609 4924
rect 3313 4870 3359 4922
rect 3359 4870 3369 4922
rect 3393 4870 3423 4922
rect 3423 4870 3435 4922
rect 3435 4870 3449 4922
rect 3473 4870 3487 4922
rect 3487 4870 3499 4922
rect 3499 4870 3529 4922
rect 3553 4870 3563 4922
rect 3563 4870 3609 4922
rect 3313 4868 3369 4870
rect 3393 4868 3449 4870
rect 3473 4868 3529 4870
rect 3553 4868 3609 4870
rect 2841 4378 2897 4380
rect 2921 4378 2977 4380
rect 3001 4378 3057 4380
rect 3081 4378 3137 4380
rect 2841 4326 2887 4378
rect 2887 4326 2897 4378
rect 2921 4326 2951 4378
rect 2951 4326 2963 4378
rect 2963 4326 2977 4378
rect 3001 4326 3015 4378
rect 3015 4326 3027 4378
rect 3027 4326 3057 4378
rect 3081 4326 3091 4378
rect 3091 4326 3137 4378
rect 2841 4324 2897 4326
rect 2921 4324 2977 4326
rect 3001 4324 3057 4326
rect 3081 4324 3137 4326
rect 3313 3834 3369 3836
rect 3393 3834 3449 3836
rect 3473 3834 3529 3836
rect 3553 3834 3609 3836
rect 3313 3782 3359 3834
rect 3359 3782 3369 3834
rect 3393 3782 3423 3834
rect 3423 3782 3435 3834
rect 3435 3782 3449 3834
rect 3473 3782 3487 3834
rect 3487 3782 3499 3834
rect 3499 3782 3529 3834
rect 3553 3782 3563 3834
rect 3563 3782 3609 3834
rect 3313 3780 3369 3782
rect 3393 3780 3449 3782
rect 3473 3780 3529 3782
rect 3553 3780 3609 3782
rect 2841 3290 2897 3292
rect 2921 3290 2977 3292
rect 3001 3290 3057 3292
rect 3081 3290 3137 3292
rect 2841 3238 2887 3290
rect 2887 3238 2897 3290
rect 2921 3238 2951 3290
rect 2951 3238 2963 3290
rect 2963 3238 2977 3290
rect 3001 3238 3015 3290
rect 3015 3238 3027 3290
rect 3027 3238 3057 3290
rect 3081 3238 3091 3290
rect 3091 3238 3137 3290
rect 2841 3236 2897 3238
rect 2921 3236 2977 3238
rect 3001 3236 3057 3238
rect 3081 3236 3137 3238
rect 3784 5466 3840 5468
rect 3864 5466 3920 5468
rect 3944 5466 4000 5468
rect 4024 5466 4080 5468
rect 3784 5414 3830 5466
rect 3830 5414 3840 5466
rect 3864 5414 3894 5466
rect 3894 5414 3906 5466
rect 3906 5414 3920 5466
rect 3944 5414 3958 5466
rect 3958 5414 3970 5466
rect 3970 5414 4000 5466
rect 4024 5414 4034 5466
rect 4034 5414 4080 5466
rect 3784 5412 3840 5414
rect 3864 5412 3920 5414
rect 3944 5412 4000 5414
rect 4024 5412 4080 5414
rect 4256 6010 4312 6012
rect 4336 6010 4392 6012
rect 4416 6010 4472 6012
rect 4496 6010 4552 6012
rect 4256 5958 4302 6010
rect 4302 5958 4312 6010
rect 4336 5958 4366 6010
rect 4366 5958 4378 6010
rect 4378 5958 4392 6010
rect 4416 5958 4430 6010
rect 4430 5958 4442 6010
rect 4442 5958 4472 6010
rect 4496 5958 4506 6010
rect 4506 5958 4552 6010
rect 4256 5956 4312 5958
rect 4336 5956 4392 5958
rect 4416 5956 4472 5958
rect 4496 5956 4552 5958
rect 4256 4922 4312 4924
rect 4336 4922 4392 4924
rect 4416 4922 4472 4924
rect 4496 4922 4552 4924
rect 4256 4870 4302 4922
rect 4302 4870 4312 4922
rect 4336 4870 4366 4922
rect 4366 4870 4378 4922
rect 4378 4870 4392 4922
rect 4416 4870 4430 4922
rect 4430 4870 4442 4922
rect 4442 4870 4472 4922
rect 4496 4870 4506 4922
rect 4506 4870 4552 4922
rect 4256 4868 4312 4870
rect 4336 4868 4392 4870
rect 4416 4868 4472 4870
rect 4496 4868 4552 4870
rect 3784 4378 3840 4380
rect 3864 4378 3920 4380
rect 3944 4378 4000 4380
rect 4024 4378 4080 4380
rect 3784 4326 3830 4378
rect 3830 4326 3840 4378
rect 3864 4326 3894 4378
rect 3894 4326 3906 4378
rect 3906 4326 3920 4378
rect 3944 4326 3958 4378
rect 3958 4326 3970 4378
rect 3970 4326 4000 4378
rect 4024 4326 4034 4378
rect 4034 4326 4080 4378
rect 3784 4324 3840 4326
rect 3864 4324 3920 4326
rect 3944 4324 4000 4326
rect 4024 4324 4080 4326
rect 3784 3290 3840 3292
rect 3864 3290 3920 3292
rect 3944 3290 4000 3292
rect 4024 3290 4080 3292
rect 3784 3238 3830 3290
rect 3830 3238 3840 3290
rect 3864 3238 3894 3290
rect 3894 3238 3906 3290
rect 3906 3238 3920 3290
rect 3944 3238 3958 3290
rect 3958 3238 3970 3290
rect 3970 3238 4000 3290
rect 4024 3238 4034 3290
rect 4034 3238 4080 3290
rect 3784 3236 3840 3238
rect 3864 3236 3920 3238
rect 3944 3236 4000 3238
rect 4024 3236 4080 3238
rect 3313 2746 3369 2748
rect 3393 2746 3449 2748
rect 3473 2746 3529 2748
rect 3553 2746 3609 2748
rect 3313 2694 3359 2746
rect 3359 2694 3369 2746
rect 3393 2694 3423 2746
rect 3423 2694 3435 2746
rect 3435 2694 3449 2746
rect 3473 2694 3487 2746
rect 3487 2694 3499 2746
rect 3499 2694 3529 2746
rect 3553 2694 3563 2746
rect 3563 2694 3609 2746
rect 3313 2692 3369 2694
rect 3393 2692 3449 2694
rect 3473 2692 3529 2694
rect 3553 2692 3609 2694
rect 2686 2352 2742 2408
rect 2841 2202 2897 2204
rect 2921 2202 2977 2204
rect 3001 2202 3057 2204
rect 3081 2202 3137 2204
rect 2841 2150 2887 2202
rect 2887 2150 2897 2202
rect 2921 2150 2951 2202
rect 2951 2150 2963 2202
rect 2963 2150 2977 2202
rect 3001 2150 3015 2202
rect 3015 2150 3027 2202
rect 3027 2150 3057 2202
rect 3081 2150 3091 2202
rect 3091 2150 3137 2202
rect 2841 2148 2897 2150
rect 2921 2148 2977 2150
rect 3001 2148 3057 2150
rect 3081 2148 3137 2150
rect 3784 2202 3840 2204
rect 3864 2202 3920 2204
rect 3944 2202 4000 2204
rect 4024 2202 4080 2204
rect 3784 2150 3830 2202
rect 3830 2150 3840 2202
rect 3864 2150 3894 2202
rect 3894 2150 3906 2202
rect 3906 2150 3920 2202
rect 3944 2150 3958 2202
rect 3958 2150 3970 2202
rect 3970 2150 4000 2202
rect 4024 2150 4034 2202
rect 4034 2150 4080 2202
rect 3784 2148 3840 2150
rect 3864 2148 3920 2150
rect 3944 2148 4000 2150
rect 4024 2148 4080 2150
rect 4256 3834 4312 3836
rect 4336 3834 4392 3836
rect 4416 3834 4472 3836
rect 4496 3834 4552 3836
rect 4256 3782 4302 3834
rect 4302 3782 4312 3834
rect 4336 3782 4366 3834
rect 4366 3782 4378 3834
rect 4378 3782 4392 3834
rect 4416 3782 4430 3834
rect 4430 3782 4442 3834
rect 4442 3782 4472 3834
rect 4496 3782 4506 3834
rect 4506 3782 4552 3834
rect 4256 3780 4312 3782
rect 4336 3780 4392 3782
rect 4416 3780 4472 3782
rect 4496 3780 4552 3782
rect 4256 2746 4312 2748
rect 4336 2746 4392 2748
rect 4416 2746 4472 2748
rect 4496 2746 4552 2748
rect 4256 2694 4302 2746
rect 4302 2694 4312 2746
rect 4336 2694 4366 2746
rect 4366 2694 4378 2746
rect 4378 2694 4392 2746
rect 4416 2694 4430 2746
rect 4430 2694 4442 2746
rect 4442 2694 4472 2746
rect 4496 2694 4506 2746
rect 4506 2694 4552 2746
rect 4256 2692 4312 2694
rect 4336 2692 4392 2694
rect 4416 2692 4472 2694
rect 4496 2692 4552 2694
rect 1427 1658 1483 1660
rect 1507 1658 1563 1660
rect 1587 1658 1643 1660
rect 1667 1658 1723 1660
rect 1427 1606 1473 1658
rect 1473 1606 1483 1658
rect 1507 1606 1537 1658
rect 1537 1606 1549 1658
rect 1549 1606 1563 1658
rect 1587 1606 1601 1658
rect 1601 1606 1613 1658
rect 1613 1606 1643 1658
rect 1667 1606 1677 1658
rect 1677 1606 1723 1658
rect 1427 1604 1483 1606
rect 1507 1604 1563 1606
rect 1587 1604 1643 1606
rect 1667 1604 1723 1606
rect 2370 1658 2426 1660
rect 2450 1658 2506 1660
rect 2530 1658 2586 1660
rect 2610 1658 2666 1660
rect 2370 1606 2416 1658
rect 2416 1606 2426 1658
rect 2450 1606 2480 1658
rect 2480 1606 2492 1658
rect 2492 1606 2506 1658
rect 2530 1606 2544 1658
rect 2544 1606 2556 1658
rect 2556 1606 2586 1658
rect 2610 1606 2620 1658
rect 2620 1606 2666 1658
rect 2370 1604 2426 1606
rect 2450 1604 2506 1606
rect 2530 1604 2586 1606
rect 2610 1604 2666 1606
rect 3313 1658 3369 1660
rect 3393 1658 3449 1660
rect 3473 1658 3529 1660
rect 3553 1658 3609 1660
rect 3313 1606 3359 1658
rect 3359 1606 3369 1658
rect 3393 1606 3423 1658
rect 3423 1606 3435 1658
rect 3435 1606 3449 1658
rect 3473 1606 3487 1658
rect 3487 1606 3499 1658
rect 3499 1606 3529 1658
rect 3553 1606 3563 1658
rect 3563 1606 3609 1658
rect 3313 1604 3369 1606
rect 3393 1604 3449 1606
rect 3473 1604 3529 1606
rect 3553 1604 3609 1606
rect 1898 1114 1954 1116
rect 1978 1114 2034 1116
rect 2058 1114 2114 1116
rect 2138 1114 2194 1116
rect 1898 1062 1944 1114
rect 1944 1062 1954 1114
rect 1978 1062 2008 1114
rect 2008 1062 2020 1114
rect 2020 1062 2034 1114
rect 2058 1062 2072 1114
rect 2072 1062 2084 1114
rect 2084 1062 2114 1114
rect 2138 1062 2148 1114
rect 2148 1062 2194 1114
rect 1898 1060 1954 1062
rect 1978 1060 2034 1062
rect 2058 1060 2114 1062
rect 2138 1060 2194 1062
rect 2841 1114 2897 1116
rect 2921 1114 2977 1116
rect 3001 1114 3057 1116
rect 3081 1114 3137 1116
rect 2841 1062 2887 1114
rect 2887 1062 2897 1114
rect 2921 1062 2951 1114
rect 2951 1062 2963 1114
rect 2963 1062 2977 1114
rect 3001 1062 3015 1114
rect 3015 1062 3027 1114
rect 3027 1062 3057 1114
rect 3081 1062 3091 1114
rect 3091 1062 3137 1114
rect 2841 1060 2897 1062
rect 2921 1060 2977 1062
rect 3001 1060 3057 1062
rect 3081 1060 3137 1062
rect 3784 1114 3840 1116
rect 3864 1114 3920 1116
rect 3944 1114 4000 1116
rect 4024 1114 4080 1116
rect 3784 1062 3830 1114
rect 3830 1062 3840 1114
rect 3864 1062 3894 1114
rect 3894 1062 3906 1114
rect 3906 1062 3920 1114
rect 3944 1062 3958 1114
rect 3958 1062 3970 1114
rect 3970 1062 4000 1114
rect 4024 1062 4034 1114
rect 4034 1062 4080 1114
rect 3784 1060 3840 1062
rect 3864 1060 3920 1062
rect 3944 1060 4000 1062
rect 4024 1060 4080 1062
rect 4256 1658 4312 1660
rect 4336 1658 4392 1660
rect 4416 1658 4472 1660
rect 4496 1658 4552 1660
rect 4256 1606 4302 1658
rect 4302 1606 4312 1658
rect 4336 1606 4366 1658
rect 4366 1606 4378 1658
rect 4378 1606 4392 1658
rect 4416 1606 4430 1658
rect 4430 1606 4442 1658
rect 4442 1606 4472 1658
rect 4496 1606 4506 1658
rect 4506 1606 4552 1658
rect 4256 1604 4312 1606
rect 4336 1604 4392 1606
rect 4416 1604 4472 1606
rect 4496 1604 4552 1606
rect 4727 5466 4783 5468
rect 4807 5466 4863 5468
rect 4887 5466 4943 5468
rect 4967 5466 5023 5468
rect 4727 5414 4773 5466
rect 4773 5414 4783 5466
rect 4807 5414 4837 5466
rect 4837 5414 4849 5466
rect 4849 5414 4863 5466
rect 4887 5414 4901 5466
rect 4901 5414 4913 5466
rect 4913 5414 4943 5466
rect 4967 5414 4977 5466
rect 4977 5414 5023 5466
rect 4727 5412 4783 5414
rect 4807 5412 4863 5414
rect 4887 5412 4943 5414
rect 4967 5412 5023 5414
rect 5078 5208 5134 5264
rect 4727 4378 4783 4380
rect 4807 4378 4863 4380
rect 4887 4378 4943 4380
rect 4967 4378 5023 4380
rect 4727 4326 4773 4378
rect 4773 4326 4783 4378
rect 4807 4326 4837 4378
rect 4837 4326 4849 4378
rect 4849 4326 4863 4378
rect 4887 4326 4901 4378
rect 4901 4326 4913 4378
rect 4913 4326 4943 4378
rect 4967 4326 4977 4378
rect 4977 4326 5023 4378
rect 4727 4324 4783 4326
rect 4807 4324 4863 4326
rect 4887 4324 4943 4326
rect 4967 4324 5023 4326
rect 5446 12416 5502 12472
rect 5078 3712 5134 3768
rect 4727 3290 4783 3292
rect 4807 3290 4863 3292
rect 4887 3290 4943 3292
rect 4967 3290 5023 3292
rect 4727 3238 4773 3290
rect 4773 3238 4783 3290
rect 4807 3238 4837 3290
rect 4837 3238 4849 3290
rect 4849 3238 4863 3290
rect 4887 3238 4901 3290
rect 4901 3238 4913 3290
rect 4913 3238 4943 3290
rect 4967 3238 4977 3290
rect 4977 3238 5023 3290
rect 4727 3236 4783 3238
rect 4807 3236 4863 3238
rect 4887 3236 4943 3238
rect 4967 3236 5023 3238
rect 4727 2202 4783 2204
rect 4807 2202 4863 2204
rect 4887 2202 4943 2204
rect 4967 2202 5023 2204
rect 4727 2150 4773 2202
rect 4773 2150 4783 2202
rect 4807 2150 4837 2202
rect 4837 2150 4849 2202
rect 4849 2150 4863 2202
rect 4887 2150 4901 2202
rect 4901 2150 4913 2202
rect 4913 2150 4943 2202
rect 4967 2150 4977 2202
rect 4977 2150 5023 2202
rect 4727 2148 4783 2150
rect 4807 2148 4863 2150
rect 4887 2148 4943 2150
rect 4967 2148 5023 2150
rect 4727 1114 4783 1116
rect 4807 1114 4863 1116
rect 4887 1114 4943 1116
rect 4967 1114 5023 1116
rect 4727 1062 4773 1114
rect 4773 1062 4783 1114
rect 4807 1062 4837 1114
rect 4837 1062 4849 1114
rect 4849 1062 4863 1114
rect 4887 1062 4901 1114
rect 4901 1062 4913 1114
rect 4913 1062 4943 1114
rect 4967 1062 4977 1114
rect 4977 1062 5023 1114
rect 4727 1060 4783 1062
rect 4807 1060 4863 1062
rect 4887 1060 4943 1062
rect 4967 1060 5023 1062
rect 5078 720 5134 776
<< metal3 >>
rect 5073 23218 5139 23221
rect 5200 23218 6000 23248
rect 5073 23216 6000 23218
rect 5073 23160 5078 23216
rect 5134 23160 6000 23216
rect 5073 23158 6000 23160
rect 5073 23155 5139 23158
rect 5200 23128 6000 23158
rect 1888 22880 2204 22881
rect 1888 22816 1894 22880
rect 1958 22816 1974 22880
rect 2038 22816 2054 22880
rect 2118 22816 2134 22880
rect 2198 22816 2204 22880
rect 1888 22815 2204 22816
rect 2831 22880 3147 22881
rect 2831 22816 2837 22880
rect 2901 22816 2917 22880
rect 2981 22816 2997 22880
rect 3061 22816 3077 22880
rect 3141 22816 3147 22880
rect 2831 22815 3147 22816
rect 3774 22880 4090 22881
rect 3774 22816 3780 22880
rect 3844 22816 3860 22880
rect 3924 22816 3940 22880
rect 4004 22816 4020 22880
rect 4084 22816 4090 22880
rect 3774 22815 4090 22816
rect 4717 22880 5033 22881
rect 4717 22816 4723 22880
rect 4787 22816 4803 22880
rect 4867 22816 4883 22880
rect 4947 22816 4963 22880
rect 5027 22816 5033 22880
rect 4717 22815 5033 22816
rect 1417 22336 1733 22337
rect 1417 22272 1423 22336
rect 1487 22272 1503 22336
rect 1567 22272 1583 22336
rect 1647 22272 1663 22336
rect 1727 22272 1733 22336
rect 1417 22271 1733 22272
rect 2360 22336 2676 22337
rect 2360 22272 2366 22336
rect 2430 22272 2446 22336
rect 2510 22272 2526 22336
rect 2590 22272 2606 22336
rect 2670 22272 2676 22336
rect 2360 22271 2676 22272
rect 3303 22336 3619 22337
rect 3303 22272 3309 22336
rect 3373 22272 3389 22336
rect 3453 22272 3469 22336
rect 3533 22272 3549 22336
rect 3613 22272 3619 22336
rect 3303 22271 3619 22272
rect 4246 22336 4562 22337
rect 4246 22272 4252 22336
rect 4316 22272 4332 22336
rect 4396 22272 4412 22336
rect 4476 22272 4492 22336
rect 4556 22272 4562 22336
rect 4246 22271 4562 22272
rect 1888 21792 2204 21793
rect 1888 21728 1894 21792
rect 1958 21728 1974 21792
rect 2038 21728 2054 21792
rect 2118 21728 2134 21792
rect 2198 21728 2204 21792
rect 1888 21727 2204 21728
rect 2831 21792 3147 21793
rect 2831 21728 2837 21792
rect 2901 21728 2917 21792
rect 2981 21728 2997 21792
rect 3061 21728 3077 21792
rect 3141 21728 3147 21792
rect 2831 21727 3147 21728
rect 3774 21792 4090 21793
rect 3774 21728 3780 21792
rect 3844 21728 3860 21792
rect 3924 21728 3940 21792
rect 4004 21728 4020 21792
rect 4084 21728 4090 21792
rect 3774 21727 4090 21728
rect 4717 21792 5033 21793
rect 4717 21728 4723 21792
rect 4787 21728 4803 21792
rect 4867 21728 4883 21792
rect 4947 21728 4963 21792
rect 5027 21728 5033 21792
rect 4717 21727 5033 21728
rect 5200 21722 6000 21752
rect 5168 21632 6000 21722
rect 5168 21453 5228 21632
rect 5165 21448 5231 21453
rect 5165 21392 5170 21448
rect 5226 21392 5231 21448
rect 5165 21387 5231 21392
rect 1417 21248 1733 21249
rect 1417 21184 1423 21248
rect 1487 21184 1503 21248
rect 1567 21184 1583 21248
rect 1647 21184 1663 21248
rect 1727 21184 1733 21248
rect 1417 21183 1733 21184
rect 2360 21248 2676 21249
rect 2360 21184 2366 21248
rect 2430 21184 2446 21248
rect 2510 21184 2526 21248
rect 2590 21184 2606 21248
rect 2670 21184 2676 21248
rect 2360 21183 2676 21184
rect 3303 21248 3619 21249
rect 3303 21184 3309 21248
rect 3373 21184 3389 21248
rect 3453 21184 3469 21248
rect 3533 21184 3549 21248
rect 3613 21184 3619 21248
rect 3303 21183 3619 21184
rect 4246 21248 4562 21249
rect 4246 21184 4252 21248
rect 4316 21184 4332 21248
rect 4396 21184 4412 21248
rect 4476 21184 4492 21248
rect 4556 21184 4562 21248
rect 4246 21183 4562 21184
rect 1888 20704 2204 20705
rect 1888 20640 1894 20704
rect 1958 20640 1974 20704
rect 2038 20640 2054 20704
rect 2118 20640 2134 20704
rect 2198 20640 2204 20704
rect 1888 20639 2204 20640
rect 2831 20704 3147 20705
rect 2831 20640 2837 20704
rect 2901 20640 2917 20704
rect 2981 20640 2997 20704
rect 3061 20640 3077 20704
rect 3141 20640 3147 20704
rect 2831 20639 3147 20640
rect 3774 20704 4090 20705
rect 3774 20640 3780 20704
rect 3844 20640 3860 20704
rect 3924 20640 3940 20704
rect 4004 20640 4020 20704
rect 4084 20640 4090 20704
rect 3774 20639 4090 20640
rect 4717 20704 5033 20705
rect 4717 20640 4723 20704
rect 4787 20640 4803 20704
rect 4867 20640 4883 20704
rect 4947 20640 4963 20704
rect 5027 20640 5033 20704
rect 4717 20639 5033 20640
rect 5200 20226 6000 20256
rect 5030 20166 6000 20226
rect 1417 20160 1733 20161
rect 1417 20096 1423 20160
rect 1487 20096 1503 20160
rect 1567 20096 1583 20160
rect 1647 20096 1663 20160
rect 1727 20096 1733 20160
rect 1417 20095 1733 20096
rect 2360 20160 2676 20161
rect 2360 20096 2366 20160
rect 2430 20096 2446 20160
rect 2510 20096 2526 20160
rect 2590 20096 2606 20160
rect 2670 20096 2676 20160
rect 2360 20095 2676 20096
rect 3303 20160 3619 20161
rect 3303 20096 3309 20160
rect 3373 20096 3389 20160
rect 3453 20096 3469 20160
rect 3533 20096 3549 20160
rect 3613 20096 3619 20160
rect 3303 20095 3619 20096
rect 4246 20160 4562 20161
rect 4246 20096 4252 20160
rect 4316 20096 4332 20160
rect 4396 20096 4412 20160
rect 4476 20096 4492 20160
rect 4556 20096 4562 20160
rect 4246 20095 4562 20096
rect 5030 19954 5090 20166
rect 5200 20136 6000 20166
rect 5533 19954 5599 19957
rect 5030 19952 5599 19954
rect 5030 19896 5538 19952
rect 5594 19896 5599 19952
rect 5030 19894 5599 19896
rect 5533 19891 5599 19894
rect 1888 19616 2204 19617
rect 1888 19552 1894 19616
rect 1958 19552 1974 19616
rect 2038 19552 2054 19616
rect 2118 19552 2134 19616
rect 2198 19552 2204 19616
rect 1888 19551 2204 19552
rect 2831 19616 3147 19617
rect 2831 19552 2837 19616
rect 2901 19552 2917 19616
rect 2981 19552 2997 19616
rect 3061 19552 3077 19616
rect 3141 19552 3147 19616
rect 2831 19551 3147 19552
rect 3774 19616 4090 19617
rect 3774 19552 3780 19616
rect 3844 19552 3860 19616
rect 3924 19552 3940 19616
rect 4004 19552 4020 19616
rect 4084 19552 4090 19616
rect 3774 19551 4090 19552
rect 4717 19616 5033 19617
rect 4717 19552 4723 19616
rect 4787 19552 4803 19616
rect 4867 19552 4883 19616
rect 4947 19552 4963 19616
rect 5027 19552 5033 19616
rect 4717 19551 5033 19552
rect 1417 19072 1733 19073
rect 1417 19008 1423 19072
rect 1487 19008 1503 19072
rect 1567 19008 1583 19072
rect 1647 19008 1663 19072
rect 1727 19008 1733 19072
rect 1417 19007 1733 19008
rect 2360 19072 2676 19073
rect 2360 19008 2366 19072
rect 2430 19008 2446 19072
rect 2510 19008 2526 19072
rect 2590 19008 2606 19072
rect 2670 19008 2676 19072
rect 2360 19007 2676 19008
rect 3303 19072 3619 19073
rect 3303 19008 3309 19072
rect 3373 19008 3389 19072
rect 3453 19008 3469 19072
rect 3533 19008 3549 19072
rect 3613 19008 3619 19072
rect 3303 19007 3619 19008
rect 4246 19072 4562 19073
rect 4246 19008 4252 19072
rect 4316 19008 4332 19072
rect 4396 19008 4412 19072
rect 4476 19008 4492 19072
rect 4556 19008 4562 19072
rect 4246 19007 4562 19008
rect 4613 18730 4679 18733
rect 5200 18730 6000 18760
rect 4613 18728 6000 18730
rect 4613 18672 4618 18728
rect 4674 18672 6000 18728
rect 4613 18670 6000 18672
rect 4613 18667 4679 18670
rect 5200 18640 6000 18670
rect 1888 18528 2204 18529
rect 1888 18464 1894 18528
rect 1958 18464 1974 18528
rect 2038 18464 2054 18528
rect 2118 18464 2134 18528
rect 2198 18464 2204 18528
rect 1888 18463 2204 18464
rect 2831 18528 3147 18529
rect 2831 18464 2837 18528
rect 2901 18464 2917 18528
rect 2981 18464 2997 18528
rect 3061 18464 3077 18528
rect 3141 18464 3147 18528
rect 2831 18463 3147 18464
rect 3774 18528 4090 18529
rect 3774 18464 3780 18528
rect 3844 18464 3860 18528
rect 3924 18464 3940 18528
rect 4004 18464 4020 18528
rect 4084 18464 4090 18528
rect 3774 18463 4090 18464
rect 4717 18528 5033 18529
rect 4717 18464 4723 18528
rect 4787 18464 4803 18528
rect 4867 18464 4883 18528
rect 4947 18464 4963 18528
rect 5027 18464 5033 18528
rect 4717 18463 5033 18464
rect 1417 17984 1733 17985
rect 1417 17920 1423 17984
rect 1487 17920 1503 17984
rect 1567 17920 1583 17984
rect 1647 17920 1663 17984
rect 1727 17920 1733 17984
rect 1417 17919 1733 17920
rect 2360 17984 2676 17985
rect 2360 17920 2366 17984
rect 2430 17920 2446 17984
rect 2510 17920 2526 17984
rect 2590 17920 2606 17984
rect 2670 17920 2676 17984
rect 2360 17919 2676 17920
rect 3303 17984 3619 17985
rect 3303 17920 3309 17984
rect 3373 17920 3389 17984
rect 3453 17920 3469 17984
rect 3533 17920 3549 17984
rect 3613 17920 3619 17984
rect 3303 17919 3619 17920
rect 4246 17984 4562 17985
rect 4246 17920 4252 17984
rect 4316 17920 4332 17984
rect 4396 17920 4412 17984
rect 4476 17920 4492 17984
rect 4556 17920 4562 17984
rect 4246 17919 4562 17920
rect 1888 17440 2204 17441
rect 1888 17376 1894 17440
rect 1958 17376 1974 17440
rect 2038 17376 2054 17440
rect 2118 17376 2134 17440
rect 2198 17376 2204 17440
rect 1888 17375 2204 17376
rect 2831 17440 3147 17441
rect 2831 17376 2837 17440
rect 2901 17376 2917 17440
rect 2981 17376 2997 17440
rect 3061 17376 3077 17440
rect 3141 17376 3147 17440
rect 2831 17375 3147 17376
rect 3774 17440 4090 17441
rect 3774 17376 3780 17440
rect 3844 17376 3860 17440
rect 3924 17376 3940 17440
rect 4004 17376 4020 17440
rect 4084 17376 4090 17440
rect 3774 17375 4090 17376
rect 4717 17440 5033 17441
rect 4717 17376 4723 17440
rect 4787 17376 4803 17440
rect 4867 17376 4883 17440
rect 4947 17376 4963 17440
rect 5027 17376 5033 17440
rect 4717 17375 5033 17376
rect 5073 17234 5139 17237
rect 5200 17234 6000 17264
rect 5073 17232 6000 17234
rect 5073 17176 5078 17232
rect 5134 17176 6000 17232
rect 5073 17174 6000 17176
rect 5073 17171 5139 17174
rect 5200 17144 6000 17174
rect 1417 16896 1733 16897
rect 1417 16832 1423 16896
rect 1487 16832 1503 16896
rect 1567 16832 1583 16896
rect 1647 16832 1663 16896
rect 1727 16832 1733 16896
rect 1417 16831 1733 16832
rect 2360 16896 2676 16897
rect 2360 16832 2366 16896
rect 2430 16832 2446 16896
rect 2510 16832 2526 16896
rect 2590 16832 2606 16896
rect 2670 16832 2676 16896
rect 2360 16831 2676 16832
rect 3303 16896 3619 16897
rect 3303 16832 3309 16896
rect 3373 16832 3389 16896
rect 3453 16832 3469 16896
rect 3533 16832 3549 16896
rect 3613 16832 3619 16896
rect 3303 16831 3619 16832
rect 4246 16896 4562 16897
rect 4246 16832 4252 16896
rect 4316 16832 4332 16896
rect 4396 16832 4412 16896
rect 4476 16832 4492 16896
rect 4556 16832 4562 16896
rect 4246 16831 4562 16832
rect 1888 16352 2204 16353
rect 1888 16288 1894 16352
rect 1958 16288 1974 16352
rect 2038 16288 2054 16352
rect 2118 16288 2134 16352
rect 2198 16288 2204 16352
rect 1888 16287 2204 16288
rect 2831 16352 3147 16353
rect 2831 16288 2837 16352
rect 2901 16288 2917 16352
rect 2981 16288 2997 16352
rect 3061 16288 3077 16352
rect 3141 16288 3147 16352
rect 2831 16287 3147 16288
rect 3774 16352 4090 16353
rect 3774 16288 3780 16352
rect 3844 16288 3860 16352
rect 3924 16288 3940 16352
rect 4004 16288 4020 16352
rect 4084 16288 4090 16352
rect 3774 16287 4090 16288
rect 4717 16352 5033 16353
rect 4717 16288 4723 16352
rect 4787 16288 4803 16352
rect 4867 16288 4883 16352
rect 4947 16288 4963 16352
rect 5027 16288 5033 16352
rect 4717 16287 5033 16288
rect 1417 15808 1733 15809
rect 1417 15744 1423 15808
rect 1487 15744 1503 15808
rect 1567 15744 1583 15808
rect 1647 15744 1663 15808
rect 1727 15744 1733 15808
rect 1417 15743 1733 15744
rect 2360 15808 2676 15809
rect 2360 15744 2366 15808
rect 2430 15744 2446 15808
rect 2510 15744 2526 15808
rect 2590 15744 2606 15808
rect 2670 15744 2676 15808
rect 2360 15743 2676 15744
rect 3303 15808 3619 15809
rect 3303 15744 3309 15808
rect 3373 15744 3389 15808
rect 3453 15744 3469 15808
rect 3533 15744 3549 15808
rect 3613 15744 3619 15808
rect 3303 15743 3619 15744
rect 4246 15808 4562 15809
rect 4246 15744 4252 15808
rect 4316 15744 4332 15808
rect 4396 15744 4412 15808
rect 4476 15744 4492 15808
rect 4556 15744 4562 15808
rect 4246 15743 4562 15744
rect 5200 15738 6000 15768
rect 4662 15678 6000 15738
rect 3693 15602 3759 15605
rect 4662 15602 4722 15678
rect 5200 15648 6000 15678
rect 3693 15600 4722 15602
rect 3693 15544 3698 15600
rect 3754 15544 4722 15600
rect 3693 15542 4722 15544
rect 3693 15539 3759 15542
rect 1888 15264 2204 15265
rect 1888 15200 1894 15264
rect 1958 15200 1974 15264
rect 2038 15200 2054 15264
rect 2118 15200 2134 15264
rect 2198 15200 2204 15264
rect 1888 15199 2204 15200
rect 2831 15264 3147 15265
rect 2831 15200 2837 15264
rect 2901 15200 2917 15264
rect 2981 15200 2997 15264
rect 3061 15200 3077 15264
rect 3141 15200 3147 15264
rect 2831 15199 3147 15200
rect 3774 15264 4090 15265
rect 3774 15200 3780 15264
rect 3844 15200 3860 15264
rect 3924 15200 3940 15264
rect 4004 15200 4020 15264
rect 4084 15200 4090 15264
rect 3774 15199 4090 15200
rect 4717 15264 5033 15265
rect 4717 15200 4723 15264
rect 4787 15200 4803 15264
rect 4867 15200 4883 15264
rect 4947 15200 4963 15264
rect 5027 15200 5033 15264
rect 4717 15199 5033 15200
rect 1417 14720 1733 14721
rect 1417 14656 1423 14720
rect 1487 14656 1503 14720
rect 1567 14656 1583 14720
rect 1647 14656 1663 14720
rect 1727 14656 1733 14720
rect 1417 14655 1733 14656
rect 2360 14720 2676 14721
rect 2360 14656 2366 14720
rect 2430 14656 2446 14720
rect 2510 14656 2526 14720
rect 2590 14656 2606 14720
rect 2670 14656 2676 14720
rect 2360 14655 2676 14656
rect 3303 14720 3619 14721
rect 3303 14656 3309 14720
rect 3373 14656 3389 14720
rect 3453 14656 3469 14720
rect 3533 14656 3549 14720
rect 3613 14656 3619 14720
rect 3303 14655 3619 14656
rect 4246 14720 4562 14721
rect 4246 14656 4252 14720
rect 4316 14656 4332 14720
rect 4396 14656 4412 14720
rect 4476 14656 4492 14720
rect 4556 14656 4562 14720
rect 4246 14655 4562 14656
rect 5349 14514 5415 14517
rect 5168 14512 5415 14514
rect 5168 14456 5354 14512
rect 5410 14456 5415 14512
rect 5168 14454 5415 14456
rect 5168 14272 5228 14454
rect 5349 14451 5415 14454
rect 5168 14182 6000 14272
rect 1888 14176 2204 14177
rect 1888 14112 1894 14176
rect 1958 14112 1974 14176
rect 2038 14112 2054 14176
rect 2118 14112 2134 14176
rect 2198 14112 2204 14176
rect 1888 14111 2204 14112
rect 2831 14176 3147 14177
rect 2831 14112 2837 14176
rect 2901 14112 2917 14176
rect 2981 14112 2997 14176
rect 3061 14112 3077 14176
rect 3141 14112 3147 14176
rect 2831 14111 3147 14112
rect 3774 14176 4090 14177
rect 3774 14112 3780 14176
rect 3844 14112 3860 14176
rect 3924 14112 3940 14176
rect 4004 14112 4020 14176
rect 4084 14112 4090 14176
rect 3774 14111 4090 14112
rect 4717 14176 5033 14177
rect 4717 14112 4723 14176
rect 4787 14112 4803 14176
rect 4867 14112 4883 14176
rect 4947 14112 4963 14176
rect 5027 14112 5033 14176
rect 5200 14152 6000 14182
rect 4717 14111 5033 14112
rect 1417 13632 1733 13633
rect 1417 13568 1423 13632
rect 1487 13568 1503 13632
rect 1567 13568 1583 13632
rect 1647 13568 1663 13632
rect 1727 13568 1733 13632
rect 1417 13567 1733 13568
rect 2360 13632 2676 13633
rect 2360 13568 2366 13632
rect 2430 13568 2446 13632
rect 2510 13568 2526 13632
rect 2590 13568 2606 13632
rect 2670 13568 2676 13632
rect 2360 13567 2676 13568
rect 3303 13632 3619 13633
rect 3303 13568 3309 13632
rect 3373 13568 3389 13632
rect 3453 13568 3469 13632
rect 3533 13568 3549 13632
rect 3613 13568 3619 13632
rect 3303 13567 3619 13568
rect 4246 13632 4562 13633
rect 4246 13568 4252 13632
rect 4316 13568 4332 13632
rect 4396 13568 4412 13632
rect 4476 13568 4492 13632
rect 4556 13568 4562 13632
rect 4246 13567 4562 13568
rect 1888 13088 2204 13089
rect 1888 13024 1894 13088
rect 1958 13024 1974 13088
rect 2038 13024 2054 13088
rect 2118 13024 2134 13088
rect 2198 13024 2204 13088
rect 1888 13023 2204 13024
rect 2831 13088 3147 13089
rect 2831 13024 2837 13088
rect 2901 13024 2917 13088
rect 2981 13024 2997 13088
rect 3061 13024 3077 13088
rect 3141 13024 3147 13088
rect 2831 13023 3147 13024
rect 3774 13088 4090 13089
rect 3774 13024 3780 13088
rect 3844 13024 3860 13088
rect 3924 13024 3940 13088
rect 4004 13024 4020 13088
rect 4084 13024 4090 13088
rect 3774 13023 4090 13024
rect 4717 13088 5033 13089
rect 4717 13024 4723 13088
rect 4787 13024 4803 13088
rect 4867 13024 4883 13088
rect 4947 13024 4963 13088
rect 5027 13024 5033 13088
rect 4717 13023 5033 13024
rect 5200 12746 6000 12776
rect 5076 12686 6000 12746
rect 1417 12544 1733 12545
rect 1417 12480 1423 12544
rect 1487 12480 1503 12544
rect 1567 12480 1583 12544
rect 1647 12480 1663 12544
rect 1727 12480 1733 12544
rect 1417 12479 1733 12480
rect 2360 12544 2676 12545
rect 2360 12480 2366 12544
rect 2430 12480 2446 12544
rect 2510 12480 2526 12544
rect 2590 12480 2606 12544
rect 2670 12480 2676 12544
rect 2360 12479 2676 12480
rect 3303 12544 3619 12545
rect 3303 12480 3309 12544
rect 3373 12480 3389 12544
rect 3453 12480 3469 12544
rect 3533 12480 3549 12544
rect 3613 12480 3619 12544
rect 3303 12479 3619 12480
rect 4246 12544 4562 12545
rect 4246 12480 4252 12544
rect 4316 12480 4332 12544
rect 4396 12480 4412 12544
rect 4476 12480 4492 12544
rect 4556 12480 4562 12544
rect 4246 12479 4562 12480
rect 5076 12474 5136 12686
rect 5200 12656 6000 12686
rect 5441 12474 5507 12477
rect 5076 12472 5507 12474
rect 5076 12416 5446 12472
rect 5502 12416 5507 12472
rect 5076 12414 5507 12416
rect 5441 12411 5507 12414
rect 1888 12000 2204 12001
rect 1888 11936 1894 12000
rect 1958 11936 1974 12000
rect 2038 11936 2054 12000
rect 2118 11936 2134 12000
rect 2198 11936 2204 12000
rect 1888 11935 2204 11936
rect 2831 12000 3147 12001
rect 2831 11936 2837 12000
rect 2901 11936 2917 12000
rect 2981 11936 2997 12000
rect 3061 11936 3077 12000
rect 3141 11936 3147 12000
rect 2831 11935 3147 11936
rect 3774 12000 4090 12001
rect 3774 11936 3780 12000
rect 3844 11936 3860 12000
rect 3924 11936 3940 12000
rect 4004 11936 4020 12000
rect 4084 11936 4090 12000
rect 3774 11935 4090 11936
rect 4717 12000 5033 12001
rect 4717 11936 4723 12000
rect 4787 11936 4803 12000
rect 4867 11936 4883 12000
rect 4947 11936 4963 12000
rect 5027 11936 5033 12000
rect 4717 11935 5033 11936
rect 1417 11456 1733 11457
rect 1417 11392 1423 11456
rect 1487 11392 1503 11456
rect 1567 11392 1583 11456
rect 1647 11392 1663 11456
rect 1727 11392 1733 11456
rect 1417 11391 1733 11392
rect 2360 11456 2676 11457
rect 2360 11392 2366 11456
rect 2430 11392 2446 11456
rect 2510 11392 2526 11456
rect 2590 11392 2606 11456
rect 2670 11392 2676 11456
rect 2360 11391 2676 11392
rect 3303 11456 3619 11457
rect 3303 11392 3309 11456
rect 3373 11392 3389 11456
rect 3453 11392 3469 11456
rect 3533 11392 3549 11456
rect 3613 11392 3619 11456
rect 3303 11391 3619 11392
rect 4246 11456 4562 11457
rect 4246 11392 4252 11456
rect 4316 11392 4332 11456
rect 4396 11392 4412 11456
rect 4476 11392 4492 11456
rect 4556 11392 4562 11456
rect 4246 11391 4562 11392
rect 3417 11250 3483 11253
rect 5200 11250 6000 11280
rect 3417 11248 6000 11250
rect 3417 11192 3422 11248
rect 3478 11192 6000 11248
rect 3417 11190 6000 11192
rect 3417 11187 3483 11190
rect 5200 11160 6000 11190
rect 1888 10912 2204 10913
rect 1888 10848 1894 10912
rect 1958 10848 1974 10912
rect 2038 10848 2054 10912
rect 2118 10848 2134 10912
rect 2198 10848 2204 10912
rect 1888 10847 2204 10848
rect 2831 10912 3147 10913
rect 2831 10848 2837 10912
rect 2901 10848 2917 10912
rect 2981 10848 2997 10912
rect 3061 10848 3077 10912
rect 3141 10848 3147 10912
rect 2831 10847 3147 10848
rect 3774 10912 4090 10913
rect 3774 10848 3780 10912
rect 3844 10848 3860 10912
rect 3924 10848 3940 10912
rect 4004 10848 4020 10912
rect 4084 10848 4090 10912
rect 3774 10847 4090 10848
rect 4717 10912 5033 10913
rect 4717 10848 4723 10912
rect 4787 10848 4803 10912
rect 4867 10848 4883 10912
rect 4947 10848 4963 10912
rect 5027 10848 5033 10912
rect 4717 10847 5033 10848
rect 1417 10368 1733 10369
rect 1417 10304 1423 10368
rect 1487 10304 1503 10368
rect 1567 10304 1583 10368
rect 1647 10304 1663 10368
rect 1727 10304 1733 10368
rect 1417 10303 1733 10304
rect 2360 10368 2676 10369
rect 2360 10304 2366 10368
rect 2430 10304 2446 10368
rect 2510 10304 2526 10368
rect 2590 10304 2606 10368
rect 2670 10304 2676 10368
rect 2360 10303 2676 10304
rect 3303 10368 3619 10369
rect 3303 10304 3309 10368
rect 3373 10304 3389 10368
rect 3453 10304 3469 10368
rect 3533 10304 3549 10368
rect 3613 10304 3619 10368
rect 3303 10303 3619 10304
rect 4246 10368 4562 10369
rect 4246 10304 4252 10368
rect 4316 10304 4332 10368
rect 4396 10304 4412 10368
rect 4476 10304 4492 10368
rect 4556 10304 4562 10368
rect 4246 10303 4562 10304
rect 1888 9824 2204 9825
rect 1888 9760 1894 9824
rect 1958 9760 1974 9824
rect 2038 9760 2054 9824
rect 2118 9760 2134 9824
rect 2198 9760 2204 9824
rect 1888 9759 2204 9760
rect 2831 9824 3147 9825
rect 2831 9760 2837 9824
rect 2901 9760 2917 9824
rect 2981 9760 2997 9824
rect 3061 9760 3077 9824
rect 3141 9760 3147 9824
rect 2831 9759 3147 9760
rect 3774 9824 4090 9825
rect 3774 9760 3780 9824
rect 3844 9760 3860 9824
rect 3924 9760 3940 9824
rect 4004 9760 4020 9824
rect 4084 9760 4090 9824
rect 3774 9759 4090 9760
rect 4717 9824 5033 9825
rect 4717 9760 4723 9824
rect 4787 9760 4803 9824
rect 4867 9760 4883 9824
rect 4947 9760 4963 9824
rect 5027 9760 5033 9824
rect 4717 9759 5033 9760
rect 5200 9754 6000 9784
rect 5168 9690 6000 9754
rect 5030 9664 6000 9690
rect 5030 9630 5228 9664
rect 5030 9482 5090 9630
rect 5165 9482 5231 9485
rect 5030 9480 5231 9482
rect 5030 9424 5170 9480
rect 5226 9424 5231 9480
rect 5030 9422 5231 9424
rect 5165 9419 5231 9422
rect 1417 9280 1733 9281
rect 1417 9216 1423 9280
rect 1487 9216 1503 9280
rect 1567 9216 1583 9280
rect 1647 9216 1663 9280
rect 1727 9216 1733 9280
rect 1417 9215 1733 9216
rect 2360 9280 2676 9281
rect 2360 9216 2366 9280
rect 2430 9216 2446 9280
rect 2510 9216 2526 9280
rect 2590 9216 2606 9280
rect 2670 9216 2676 9280
rect 2360 9215 2676 9216
rect 3303 9280 3619 9281
rect 3303 9216 3309 9280
rect 3373 9216 3389 9280
rect 3453 9216 3469 9280
rect 3533 9216 3549 9280
rect 3613 9216 3619 9280
rect 3303 9215 3619 9216
rect 4246 9280 4562 9281
rect 4246 9216 4252 9280
rect 4316 9216 4332 9280
rect 4396 9216 4412 9280
rect 4476 9216 4492 9280
rect 4556 9216 4562 9280
rect 4246 9215 4562 9216
rect 1888 8736 2204 8737
rect 1888 8672 1894 8736
rect 1958 8672 1974 8736
rect 2038 8672 2054 8736
rect 2118 8672 2134 8736
rect 2198 8672 2204 8736
rect 1888 8671 2204 8672
rect 2831 8736 3147 8737
rect 2831 8672 2837 8736
rect 2901 8672 2917 8736
rect 2981 8672 2997 8736
rect 3061 8672 3077 8736
rect 3141 8672 3147 8736
rect 2831 8671 3147 8672
rect 3774 8736 4090 8737
rect 3774 8672 3780 8736
rect 3844 8672 3860 8736
rect 3924 8672 3940 8736
rect 4004 8672 4020 8736
rect 4084 8672 4090 8736
rect 3774 8671 4090 8672
rect 4717 8736 5033 8737
rect 4717 8672 4723 8736
rect 4787 8672 4803 8736
rect 4867 8672 4883 8736
rect 4947 8672 4963 8736
rect 5027 8672 5033 8736
rect 4717 8671 5033 8672
rect 5073 8258 5139 8261
rect 5200 8258 6000 8288
rect 5073 8256 6000 8258
rect 5073 8200 5078 8256
rect 5134 8200 6000 8256
rect 5073 8198 6000 8200
rect 5073 8195 5139 8198
rect 1417 8192 1733 8193
rect 1417 8128 1423 8192
rect 1487 8128 1503 8192
rect 1567 8128 1583 8192
rect 1647 8128 1663 8192
rect 1727 8128 1733 8192
rect 1417 8127 1733 8128
rect 2360 8192 2676 8193
rect 2360 8128 2366 8192
rect 2430 8128 2446 8192
rect 2510 8128 2526 8192
rect 2590 8128 2606 8192
rect 2670 8128 2676 8192
rect 2360 8127 2676 8128
rect 3303 8192 3619 8193
rect 3303 8128 3309 8192
rect 3373 8128 3389 8192
rect 3453 8128 3469 8192
rect 3533 8128 3549 8192
rect 3613 8128 3619 8192
rect 3303 8127 3619 8128
rect 4246 8192 4562 8193
rect 4246 8128 4252 8192
rect 4316 8128 4332 8192
rect 4396 8128 4412 8192
rect 4476 8128 4492 8192
rect 4556 8128 4562 8192
rect 5200 8168 6000 8198
rect 4246 8127 4562 8128
rect 1888 7648 2204 7649
rect 1888 7584 1894 7648
rect 1958 7584 1974 7648
rect 2038 7584 2054 7648
rect 2118 7584 2134 7648
rect 2198 7584 2204 7648
rect 1888 7583 2204 7584
rect 2831 7648 3147 7649
rect 2831 7584 2837 7648
rect 2901 7584 2917 7648
rect 2981 7584 2997 7648
rect 3061 7584 3077 7648
rect 3141 7584 3147 7648
rect 2831 7583 3147 7584
rect 3774 7648 4090 7649
rect 3774 7584 3780 7648
rect 3844 7584 3860 7648
rect 3924 7584 3940 7648
rect 4004 7584 4020 7648
rect 4084 7584 4090 7648
rect 3774 7583 4090 7584
rect 4717 7648 5033 7649
rect 4717 7584 4723 7648
rect 4787 7584 4803 7648
rect 4867 7584 4883 7648
rect 4947 7584 4963 7648
rect 5027 7584 5033 7648
rect 4717 7583 5033 7584
rect 1417 7104 1733 7105
rect 1417 7040 1423 7104
rect 1487 7040 1503 7104
rect 1567 7040 1583 7104
rect 1647 7040 1663 7104
rect 1727 7040 1733 7104
rect 1417 7039 1733 7040
rect 2360 7104 2676 7105
rect 2360 7040 2366 7104
rect 2430 7040 2446 7104
rect 2510 7040 2526 7104
rect 2590 7040 2606 7104
rect 2670 7040 2676 7104
rect 2360 7039 2676 7040
rect 3303 7104 3619 7105
rect 3303 7040 3309 7104
rect 3373 7040 3389 7104
rect 3453 7040 3469 7104
rect 3533 7040 3549 7104
rect 3613 7040 3619 7104
rect 3303 7039 3619 7040
rect 4246 7104 4562 7105
rect 4246 7040 4252 7104
rect 4316 7040 4332 7104
rect 4396 7040 4412 7104
rect 4476 7040 4492 7104
rect 4556 7040 4562 7104
rect 4246 7039 4562 7040
rect 3601 6762 3667 6765
rect 5200 6762 6000 6792
rect 3601 6760 6000 6762
rect 3601 6704 3606 6760
rect 3662 6704 6000 6760
rect 3601 6702 6000 6704
rect 3601 6699 3667 6702
rect 5200 6672 6000 6702
rect 1888 6560 2204 6561
rect 1888 6496 1894 6560
rect 1958 6496 1974 6560
rect 2038 6496 2054 6560
rect 2118 6496 2134 6560
rect 2198 6496 2204 6560
rect 1888 6495 2204 6496
rect 2831 6560 3147 6561
rect 2831 6496 2837 6560
rect 2901 6496 2917 6560
rect 2981 6496 2997 6560
rect 3061 6496 3077 6560
rect 3141 6496 3147 6560
rect 2831 6495 3147 6496
rect 3774 6560 4090 6561
rect 3774 6496 3780 6560
rect 3844 6496 3860 6560
rect 3924 6496 3940 6560
rect 4004 6496 4020 6560
rect 4084 6496 4090 6560
rect 3774 6495 4090 6496
rect 4717 6560 5033 6561
rect 4717 6496 4723 6560
rect 4787 6496 4803 6560
rect 4867 6496 4883 6560
rect 4947 6496 4963 6560
rect 5027 6496 5033 6560
rect 4717 6495 5033 6496
rect 3509 6354 3575 6357
rect 3785 6354 3851 6357
rect 3509 6352 3851 6354
rect 3509 6296 3514 6352
rect 3570 6296 3790 6352
rect 3846 6296 3851 6352
rect 3509 6294 3851 6296
rect 3509 6291 3575 6294
rect 3785 6291 3851 6294
rect 1417 6016 1733 6017
rect 1417 5952 1423 6016
rect 1487 5952 1503 6016
rect 1567 5952 1583 6016
rect 1647 5952 1663 6016
rect 1727 5952 1733 6016
rect 1417 5951 1733 5952
rect 2360 6016 2676 6017
rect 2360 5952 2366 6016
rect 2430 5952 2446 6016
rect 2510 5952 2526 6016
rect 2590 5952 2606 6016
rect 2670 5952 2676 6016
rect 2360 5951 2676 5952
rect 3303 6016 3619 6017
rect 3303 5952 3309 6016
rect 3373 5952 3389 6016
rect 3453 5952 3469 6016
rect 3533 5952 3549 6016
rect 3613 5952 3619 6016
rect 3303 5951 3619 5952
rect 4246 6016 4562 6017
rect 4246 5952 4252 6016
rect 4316 5952 4332 6016
rect 4396 5952 4412 6016
rect 4476 5952 4492 6016
rect 4556 5952 4562 6016
rect 4246 5951 4562 5952
rect 1888 5472 2204 5473
rect 1888 5408 1894 5472
rect 1958 5408 1974 5472
rect 2038 5408 2054 5472
rect 2118 5408 2134 5472
rect 2198 5408 2204 5472
rect 1888 5407 2204 5408
rect 2831 5472 3147 5473
rect 2831 5408 2837 5472
rect 2901 5408 2917 5472
rect 2981 5408 2997 5472
rect 3061 5408 3077 5472
rect 3141 5408 3147 5472
rect 2831 5407 3147 5408
rect 3774 5472 4090 5473
rect 3774 5408 3780 5472
rect 3844 5408 3860 5472
rect 3924 5408 3940 5472
rect 4004 5408 4020 5472
rect 4084 5408 4090 5472
rect 3774 5407 4090 5408
rect 4717 5472 5033 5473
rect 4717 5408 4723 5472
rect 4787 5408 4803 5472
rect 4867 5408 4883 5472
rect 4947 5408 4963 5472
rect 5027 5408 5033 5472
rect 4717 5407 5033 5408
rect 5073 5266 5139 5269
rect 5200 5266 6000 5296
rect 5073 5264 6000 5266
rect 5073 5208 5078 5264
rect 5134 5208 6000 5264
rect 5073 5206 6000 5208
rect 5073 5203 5139 5206
rect 5200 5176 6000 5206
rect 1417 4928 1733 4929
rect 1417 4864 1423 4928
rect 1487 4864 1503 4928
rect 1567 4864 1583 4928
rect 1647 4864 1663 4928
rect 1727 4864 1733 4928
rect 1417 4863 1733 4864
rect 2360 4928 2676 4929
rect 2360 4864 2366 4928
rect 2430 4864 2446 4928
rect 2510 4864 2526 4928
rect 2590 4864 2606 4928
rect 2670 4864 2676 4928
rect 2360 4863 2676 4864
rect 3303 4928 3619 4929
rect 3303 4864 3309 4928
rect 3373 4864 3389 4928
rect 3453 4864 3469 4928
rect 3533 4864 3549 4928
rect 3613 4864 3619 4928
rect 3303 4863 3619 4864
rect 4246 4928 4562 4929
rect 4246 4864 4252 4928
rect 4316 4864 4332 4928
rect 4396 4864 4412 4928
rect 4476 4864 4492 4928
rect 4556 4864 4562 4928
rect 4246 4863 4562 4864
rect 1888 4384 2204 4385
rect 1888 4320 1894 4384
rect 1958 4320 1974 4384
rect 2038 4320 2054 4384
rect 2118 4320 2134 4384
rect 2198 4320 2204 4384
rect 1888 4319 2204 4320
rect 2831 4384 3147 4385
rect 2831 4320 2837 4384
rect 2901 4320 2917 4384
rect 2981 4320 2997 4384
rect 3061 4320 3077 4384
rect 3141 4320 3147 4384
rect 2831 4319 3147 4320
rect 3774 4384 4090 4385
rect 3774 4320 3780 4384
rect 3844 4320 3860 4384
rect 3924 4320 3940 4384
rect 4004 4320 4020 4384
rect 4084 4320 4090 4384
rect 3774 4319 4090 4320
rect 4717 4384 5033 4385
rect 4717 4320 4723 4384
rect 4787 4320 4803 4384
rect 4867 4320 4883 4384
rect 4947 4320 4963 4384
rect 5027 4320 5033 4384
rect 4717 4319 5033 4320
rect 1417 3840 1733 3841
rect 1417 3776 1423 3840
rect 1487 3776 1503 3840
rect 1567 3776 1583 3840
rect 1647 3776 1663 3840
rect 1727 3776 1733 3840
rect 1417 3775 1733 3776
rect 2360 3840 2676 3841
rect 2360 3776 2366 3840
rect 2430 3776 2446 3840
rect 2510 3776 2526 3840
rect 2590 3776 2606 3840
rect 2670 3776 2676 3840
rect 2360 3775 2676 3776
rect 3303 3840 3619 3841
rect 3303 3776 3309 3840
rect 3373 3776 3389 3840
rect 3453 3776 3469 3840
rect 3533 3776 3549 3840
rect 3613 3776 3619 3840
rect 3303 3775 3619 3776
rect 4246 3840 4562 3841
rect 4246 3776 4252 3840
rect 4316 3776 4332 3840
rect 4396 3776 4412 3840
rect 4476 3776 4492 3840
rect 4556 3776 4562 3840
rect 4246 3775 4562 3776
rect 5073 3770 5139 3773
rect 5200 3770 6000 3800
rect 5073 3768 6000 3770
rect 5073 3712 5078 3768
rect 5134 3712 6000 3768
rect 5073 3710 6000 3712
rect 5073 3707 5139 3710
rect 5200 3680 6000 3710
rect 1888 3296 2204 3297
rect 1888 3232 1894 3296
rect 1958 3232 1974 3296
rect 2038 3232 2054 3296
rect 2118 3232 2134 3296
rect 2198 3232 2204 3296
rect 1888 3231 2204 3232
rect 2831 3296 3147 3297
rect 2831 3232 2837 3296
rect 2901 3232 2917 3296
rect 2981 3232 2997 3296
rect 3061 3232 3077 3296
rect 3141 3232 3147 3296
rect 2831 3231 3147 3232
rect 3774 3296 4090 3297
rect 3774 3232 3780 3296
rect 3844 3232 3860 3296
rect 3924 3232 3940 3296
rect 4004 3232 4020 3296
rect 4084 3232 4090 3296
rect 3774 3231 4090 3232
rect 4717 3296 5033 3297
rect 4717 3232 4723 3296
rect 4787 3232 4803 3296
rect 4867 3232 4883 3296
rect 4947 3232 4963 3296
rect 5027 3232 5033 3296
rect 4717 3231 5033 3232
rect 1417 2752 1733 2753
rect 1417 2688 1423 2752
rect 1487 2688 1503 2752
rect 1567 2688 1583 2752
rect 1647 2688 1663 2752
rect 1727 2688 1733 2752
rect 1417 2687 1733 2688
rect 2360 2752 2676 2753
rect 2360 2688 2366 2752
rect 2430 2688 2446 2752
rect 2510 2688 2526 2752
rect 2590 2688 2606 2752
rect 2670 2688 2676 2752
rect 2360 2687 2676 2688
rect 3303 2752 3619 2753
rect 3303 2688 3309 2752
rect 3373 2688 3389 2752
rect 3453 2688 3469 2752
rect 3533 2688 3549 2752
rect 3613 2688 3619 2752
rect 3303 2687 3619 2688
rect 4246 2752 4562 2753
rect 4246 2688 4252 2752
rect 4316 2688 4332 2752
rect 4396 2688 4412 2752
rect 4476 2688 4492 2752
rect 4556 2688 4562 2752
rect 4246 2687 4562 2688
rect 2681 2410 2747 2413
rect 2681 2408 5228 2410
rect 2681 2352 2686 2408
rect 2742 2352 5228 2408
rect 2681 2350 5228 2352
rect 2681 2347 2747 2350
rect 5168 2304 5228 2350
rect 5168 2214 6000 2304
rect 1888 2208 2204 2209
rect 1888 2144 1894 2208
rect 1958 2144 1974 2208
rect 2038 2144 2054 2208
rect 2118 2144 2134 2208
rect 2198 2144 2204 2208
rect 1888 2143 2204 2144
rect 2831 2208 3147 2209
rect 2831 2144 2837 2208
rect 2901 2144 2917 2208
rect 2981 2144 2997 2208
rect 3061 2144 3077 2208
rect 3141 2144 3147 2208
rect 2831 2143 3147 2144
rect 3774 2208 4090 2209
rect 3774 2144 3780 2208
rect 3844 2144 3860 2208
rect 3924 2144 3940 2208
rect 4004 2144 4020 2208
rect 4084 2144 4090 2208
rect 3774 2143 4090 2144
rect 4717 2208 5033 2209
rect 4717 2144 4723 2208
rect 4787 2144 4803 2208
rect 4867 2144 4883 2208
rect 4947 2144 4963 2208
rect 5027 2144 5033 2208
rect 5200 2184 6000 2214
rect 4717 2143 5033 2144
rect 1417 1664 1733 1665
rect 1417 1600 1423 1664
rect 1487 1600 1503 1664
rect 1567 1600 1583 1664
rect 1647 1600 1663 1664
rect 1727 1600 1733 1664
rect 1417 1599 1733 1600
rect 2360 1664 2676 1665
rect 2360 1600 2366 1664
rect 2430 1600 2446 1664
rect 2510 1600 2526 1664
rect 2590 1600 2606 1664
rect 2670 1600 2676 1664
rect 2360 1599 2676 1600
rect 3303 1664 3619 1665
rect 3303 1600 3309 1664
rect 3373 1600 3389 1664
rect 3453 1600 3469 1664
rect 3533 1600 3549 1664
rect 3613 1600 3619 1664
rect 3303 1599 3619 1600
rect 4246 1664 4562 1665
rect 4246 1600 4252 1664
rect 4316 1600 4332 1664
rect 4396 1600 4412 1664
rect 4476 1600 4492 1664
rect 4556 1600 4562 1664
rect 4246 1599 4562 1600
rect 1888 1120 2204 1121
rect 1888 1056 1894 1120
rect 1958 1056 1974 1120
rect 2038 1056 2054 1120
rect 2118 1056 2134 1120
rect 2198 1056 2204 1120
rect 1888 1055 2204 1056
rect 2831 1120 3147 1121
rect 2831 1056 2837 1120
rect 2901 1056 2917 1120
rect 2981 1056 2997 1120
rect 3061 1056 3077 1120
rect 3141 1056 3147 1120
rect 2831 1055 3147 1056
rect 3774 1120 4090 1121
rect 3774 1056 3780 1120
rect 3844 1056 3860 1120
rect 3924 1056 3940 1120
rect 4004 1056 4020 1120
rect 4084 1056 4090 1120
rect 3774 1055 4090 1056
rect 4717 1120 5033 1121
rect 4717 1056 4723 1120
rect 4787 1056 4803 1120
rect 4867 1056 4883 1120
rect 4947 1056 4963 1120
rect 5027 1056 5033 1120
rect 4717 1055 5033 1056
rect 5073 778 5139 781
rect 5200 778 6000 808
rect 5073 776 6000 778
rect 5073 720 5078 776
rect 5134 720 6000 776
rect 5073 718 6000 720
rect 5073 715 5139 718
rect 5200 688 6000 718
<< via3 >>
rect 1894 22876 1958 22880
rect 1894 22820 1898 22876
rect 1898 22820 1954 22876
rect 1954 22820 1958 22876
rect 1894 22816 1958 22820
rect 1974 22876 2038 22880
rect 1974 22820 1978 22876
rect 1978 22820 2034 22876
rect 2034 22820 2038 22876
rect 1974 22816 2038 22820
rect 2054 22876 2118 22880
rect 2054 22820 2058 22876
rect 2058 22820 2114 22876
rect 2114 22820 2118 22876
rect 2054 22816 2118 22820
rect 2134 22876 2198 22880
rect 2134 22820 2138 22876
rect 2138 22820 2194 22876
rect 2194 22820 2198 22876
rect 2134 22816 2198 22820
rect 2837 22876 2901 22880
rect 2837 22820 2841 22876
rect 2841 22820 2897 22876
rect 2897 22820 2901 22876
rect 2837 22816 2901 22820
rect 2917 22876 2981 22880
rect 2917 22820 2921 22876
rect 2921 22820 2977 22876
rect 2977 22820 2981 22876
rect 2917 22816 2981 22820
rect 2997 22876 3061 22880
rect 2997 22820 3001 22876
rect 3001 22820 3057 22876
rect 3057 22820 3061 22876
rect 2997 22816 3061 22820
rect 3077 22876 3141 22880
rect 3077 22820 3081 22876
rect 3081 22820 3137 22876
rect 3137 22820 3141 22876
rect 3077 22816 3141 22820
rect 3780 22876 3844 22880
rect 3780 22820 3784 22876
rect 3784 22820 3840 22876
rect 3840 22820 3844 22876
rect 3780 22816 3844 22820
rect 3860 22876 3924 22880
rect 3860 22820 3864 22876
rect 3864 22820 3920 22876
rect 3920 22820 3924 22876
rect 3860 22816 3924 22820
rect 3940 22876 4004 22880
rect 3940 22820 3944 22876
rect 3944 22820 4000 22876
rect 4000 22820 4004 22876
rect 3940 22816 4004 22820
rect 4020 22876 4084 22880
rect 4020 22820 4024 22876
rect 4024 22820 4080 22876
rect 4080 22820 4084 22876
rect 4020 22816 4084 22820
rect 4723 22876 4787 22880
rect 4723 22820 4727 22876
rect 4727 22820 4783 22876
rect 4783 22820 4787 22876
rect 4723 22816 4787 22820
rect 4803 22876 4867 22880
rect 4803 22820 4807 22876
rect 4807 22820 4863 22876
rect 4863 22820 4867 22876
rect 4803 22816 4867 22820
rect 4883 22876 4947 22880
rect 4883 22820 4887 22876
rect 4887 22820 4943 22876
rect 4943 22820 4947 22876
rect 4883 22816 4947 22820
rect 4963 22876 5027 22880
rect 4963 22820 4967 22876
rect 4967 22820 5023 22876
rect 5023 22820 5027 22876
rect 4963 22816 5027 22820
rect 1423 22332 1487 22336
rect 1423 22276 1427 22332
rect 1427 22276 1483 22332
rect 1483 22276 1487 22332
rect 1423 22272 1487 22276
rect 1503 22332 1567 22336
rect 1503 22276 1507 22332
rect 1507 22276 1563 22332
rect 1563 22276 1567 22332
rect 1503 22272 1567 22276
rect 1583 22332 1647 22336
rect 1583 22276 1587 22332
rect 1587 22276 1643 22332
rect 1643 22276 1647 22332
rect 1583 22272 1647 22276
rect 1663 22332 1727 22336
rect 1663 22276 1667 22332
rect 1667 22276 1723 22332
rect 1723 22276 1727 22332
rect 1663 22272 1727 22276
rect 2366 22332 2430 22336
rect 2366 22276 2370 22332
rect 2370 22276 2426 22332
rect 2426 22276 2430 22332
rect 2366 22272 2430 22276
rect 2446 22332 2510 22336
rect 2446 22276 2450 22332
rect 2450 22276 2506 22332
rect 2506 22276 2510 22332
rect 2446 22272 2510 22276
rect 2526 22332 2590 22336
rect 2526 22276 2530 22332
rect 2530 22276 2586 22332
rect 2586 22276 2590 22332
rect 2526 22272 2590 22276
rect 2606 22332 2670 22336
rect 2606 22276 2610 22332
rect 2610 22276 2666 22332
rect 2666 22276 2670 22332
rect 2606 22272 2670 22276
rect 3309 22332 3373 22336
rect 3309 22276 3313 22332
rect 3313 22276 3369 22332
rect 3369 22276 3373 22332
rect 3309 22272 3373 22276
rect 3389 22332 3453 22336
rect 3389 22276 3393 22332
rect 3393 22276 3449 22332
rect 3449 22276 3453 22332
rect 3389 22272 3453 22276
rect 3469 22332 3533 22336
rect 3469 22276 3473 22332
rect 3473 22276 3529 22332
rect 3529 22276 3533 22332
rect 3469 22272 3533 22276
rect 3549 22332 3613 22336
rect 3549 22276 3553 22332
rect 3553 22276 3609 22332
rect 3609 22276 3613 22332
rect 3549 22272 3613 22276
rect 4252 22332 4316 22336
rect 4252 22276 4256 22332
rect 4256 22276 4312 22332
rect 4312 22276 4316 22332
rect 4252 22272 4316 22276
rect 4332 22332 4396 22336
rect 4332 22276 4336 22332
rect 4336 22276 4392 22332
rect 4392 22276 4396 22332
rect 4332 22272 4396 22276
rect 4412 22332 4476 22336
rect 4412 22276 4416 22332
rect 4416 22276 4472 22332
rect 4472 22276 4476 22332
rect 4412 22272 4476 22276
rect 4492 22332 4556 22336
rect 4492 22276 4496 22332
rect 4496 22276 4552 22332
rect 4552 22276 4556 22332
rect 4492 22272 4556 22276
rect 1894 21788 1958 21792
rect 1894 21732 1898 21788
rect 1898 21732 1954 21788
rect 1954 21732 1958 21788
rect 1894 21728 1958 21732
rect 1974 21788 2038 21792
rect 1974 21732 1978 21788
rect 1978 21732 2034 21788
rect 2034 21732 2038 21788
rect 1974 21728 2038 21732
rect 2054 21788 2118 21792
rect 2054 21732 2058 21788
rect 2058 21732 2114 21788
rect 2114 21732 2118 21788
rect 2054 21728 2118 21732
rect 2134 21788 2198 21792
rect 2134 21732 2138 21788
rect 2138 21732 2194 21788
rect 2194 21732 2198 21788
rect 2134 21728 2198 21732
rect 2837 21788 2901 21792
rect 2837 21732 2841 21788
rect 2841 21732 2897 21788
rect 2897 21732 2901 21788
rect 2837 21728 2901 21732
rect 2917 21788 2981 21792
rect 2917 21732 2921 21788
rect 2921 21732 2977 21788
rect 2977 21732 2981 21788
rect 2917 21728 2981 21732
rect 2997 21788 3061 21792
rect 2997 21732 3001 21788
rect 3001 21732 3057 21788
rect 3057 21732 3061 21788
rect 2997 21728 3061 21732
rect 3077 21788 3141 21792
rect 3077 21732 3081 21788
rect 3081 21732 3137 21788
rect 3137 21732 3141 21788
rect 3077 21728 3141 21732
rect 3780 21788 3844 21792
rect 3780 21732 3784 21788
rect 3784 21732 3840 21788
rect 3840 21732 3844 21788
rect 3780 21728 3844 21732
rect 3860 21788 3924 21792
rect 3860 21732 3864 21788
rect 3864 21732 3920 21788
rect 3920 21732 3924 21788
rect 3860 21728 3924 21732
rect 3940 21788 4004 21792
rect 3940 21732 3944 21788
rect 3944 21732 4000 21788
rect 4000 21732 4004 21788
rect 3940 21728 4004 21732
rect 4020 21788 4084 21792
rect 4020 21732 4024 21788
rect 4024 21732 4080 21788
rect 4080 21732 4084 21788
rect 4020 21728 4084 21732
rect 4723 21788 4787 21792
rect 4723 21732 4727 21788
rect 4727 21732 4783 21788
rect 4783 21732 4787 21788
rect 4723 21728 4787 21732
rect 4803 21788 4867 21792
rect 4803 21732 4807 21788
rect 4807 21732 4863 21788
rect 4863 21732 4867 21788
rect 4803 21728 4867 21732
rect 4883 21788 4947 21792
rect 4883 21732 4887 21788
rect 4887 21732 4943 21788
rect 4943 21732 4947 21788
rect 4883 21728 4947 21732
rect 4963 21788 5027 21792
rect 4963 21732 4967 21788
rect 4967 21732 5023 21788
rect 5023 21732 5027 21788
rect 4963 21728 5027 21732
rect 1423 21244 1487 21248
rect 1423 21188 1427 21244
rect 1427 21188 1483 21244
rect 1483 21188 1487 21244
rect 1423 21184 1487 21188
rect 1503 21244 1567 21248
rect 1503 21188 1507 21244
rect 1507 21188 1563 21244
rect 1563 21188 1567 21244
rect 1503 21184 1567 21188
rect 1583 21244 1647 21248
rect 1583 21188 1587 21244
rect 1587 21188 1643 21244
rect 1643 21188 1647 21244
rect 1583 21184 1647 21188
rect 1663 21244 1727 21248
rect 1663 21188 1667 21244
rect 1667 21188 1723 21244
rect 1723 21188 1727 21244
rect 1663 21184 1727 21188
rect 2366 21244 2430 21248
rect 2366 21188 2370 21244
rect 2370 21188 2426 21244
rect 2426 21188 2430 21244
rect 2366 21184 2430 21188
rect 2446 21244 2510 21248
rect 2446 21188 2450 21244
rect 2450 21188 2506 21244
rect 2506 21188 2510 21244
rect 2446 21184 2510 21188
rect 2526 21244 2590 21248
rect 2526 21188 2530 21244
rect 2530 21188 2586 21244
rect 2586 21188 2590 21244
rect 2526 21184 2590 21188
rect 2606 21244 2670 21248
rect 2606 21188 2610 21244
rect 2610 21188 2666 21244
rect 2666 21188 2670 21244
rect 2606 21184 2670 21188
rect 3309 21244 3373 21248
rect 3309 21188 3313 21244
rect 3313 21188 3369 21244
rect 3369 21188 3373 21244
rect 3309 21184 3373 21188
rect 3389 21244 3453 21248
rect 3389 21188 3393 21244
rect 3393 21188 3449 21244
rect 3449 21188 3453 21244
rect 3389 21184 3453 21188
rect 3469 21244 3533 21248
rect 3469 21188 3473 21244
rect 3473 21188 3529 21244
rect 3529 21188 3533 21244
rect 3469 21184 3533 21188
rect 3549 21244 3613 21248
rect 3549 21188 3553 21244
rect 3553 21188 3609 21244
rect 3609 21188 3613 21244
rect 3549 21184 3613 21188
rect 4252 21244 4316 21248
rect 4252 21188 4256 21244
rect 4256 21188 4312 21244
rect 4312 21188 4316 21244
rect 4252 21184 4316 21188
rect 4332 21244 4396 21248
rect 4332 21188 4336 21244
rect 4336 21188 4392 21244
rect 4392 21188 4396 21244
rect 4332 21184 4396 21188
rect 4412 21244 4476 21248
rect 4412 21188 4416 21244
rect 4416 21188 4472 21244
rect 4472 21188 4476 21244
rect 4412 21184 4476 21188
rect 4492 21244 4556 21248
rect 4492 21188 4496 21244
rect 4496 21188 4552 21244
rect 4552 21188 4556 21244
rect 4492 21184 4556 21188
rect 1894 20700 1958 20704
rect 1894 20644 1898 20700
rect 1898 20644 1954 20700
rect 1954 20644 1958 20700
rect 1894 20640 1958 20644
rect 1974 20700 2038 20704
rect 1974 20644 1978 20700
rect 1978 20644 2034 20700
rect 2034 20644 2038 20700
rect 1974 20640 2038 20644
rect 2054 20700 2118 20704
rect 2054 20644 2058 20700
rect 2058 20644 2114 20700
rect 2114 20644 2118 20700
rect 2054 20640 2118 20644
rect 2134 20700 2198 20704
rect 2134 20644 2138 20700
rect 2138 20644 2194 20700
rect 2194 20644 2198 20700
rect 2134 20640 2198 20644
rect 2837 20700 2901 20704
rect 2837 20644 2841 20700
rect 2841 20644 2897 20700
rect 2897 20644 2901 20700
rect 2837 20640 2901 20644
rect 2917 20700 2981 20704
rect 2917 20644 2921 20700
rect 2921 20644 2977 20700
rect 2977 20644 2981 20700
rect 2917 20640 2981 20644
rect 2997 20700 3061 20704
rect 2997 20644 3001 20700
rect 3001 20644 3057 20700
rect 3057 20644 3061 20700
rect 2997 20640 3061 20644
rect 3077 20700 3141 20704
rect 3077 20644 3081 20700
rect 3081 20644 3137 20700
rect 3137 20644 3141 20700
rect 3077 20640 3141 20644
rect 3780 20700 3844 20704
rect 3780 20644 3784 20700
rect 3784 20644 3840 20700
rect 3840 20644 3844 20700
rect 3780 20640 3844 20644
rect 3860 20700 3924 20704
rect 3860 20644 3864 20700
rect 3864 20644 3920 20700
rect 3920 20644 3924 20700
rect 3860 20640 3924 20644
rect 3940 20700 4004 20704
rect 3940 20644 3944 20700
rect 3944 20644 4000 20700
rect 4000 20644 4004 20700
rect 3940 20640 4004 20644
rect 4020 20700 4084 20704
rect 4020 20644 4024 20700
rect 4024 20644 4080 20700
rect 4080 20644 4084 20700
rect 4020 20640 4084 20644
rect 4723 20700 4787 20704
rect 4723 20644 4727 20700
rect 4727 20644 4783 20700
rect 4783 20644 4787 20700
rect 4723 20640 4787 20644
rect 4803 20700 4867 20704
rect 4803 20644 4807 20700
rect 4807 20644 4863 20700
rect 4863 20644 4867 20700
rect 4803 20640 4867 20644
rect 4883 20700 4947 20704
rect 4883 20644 4887 20700
rect 4887 20644 4943 20700
rect 4943 20644 4947 20700
rect 4883 20640 4947 20644
rect 4963 20700 5027 20704
rect 4963 20644 4967 20700
rect 4967 20644 5023 20700
rect 5023 20644 5027 20700
rect 4963 20640 5027 20644
rect 1423 20156 1487 20160
rect 1423 20100 1427 20156
rect 1427 20100 1483 20156
rect 1483 20100 1487 20156
rect 1423 20096 1487 20100
rect 1503 20156 1567 20160
rect 1503 20100 1507 20156
rect 1507 20100 1563 20156
rect 1563 20100 1567 20156
rect 1503 20096 1567 20100
rect 1583 20156 1647 20160
rect 1583 20100 1587 20156
rect 1587 20100 1643 20156
rect 1643 20100 1647 20156
rect 1583 20096 1647 20100
rect 1663 20156 1727 20160
rect 1663 20100 1667 20156
rect 1667 20100 1723 20156
rect 1723 20100 1727 20156
rect 1663 20096 1727 20100
rect 2366 20156 2430 20160
rect 2366 20100 2370 20156
rect 2370 20100 2426 20156
rect 2426 20100 2430 20156
rect 2366 20096 2430 20100
rect 2446 20156 2510 20160
rect 2446 20100 2450 20156
rect 2450 20100 2506 20156
rect 2506 20100 2510 20156
rect 2446 20096 2510 20100
rect 2526 20156 2590 20160
rect 2526 20100 2530 20156
rect 2530 20100 2586 20156
rect 2586 20100 2590 20156
rect 2526 20096 2590 20100
rect 2606 20156 2670 20160
rect 2606 20100 2610 20156
rect 2610 20100 2666 20156
rect 2666 20100 2670 20156
rect 2606 20096 2670 20100
rect 3309 20156 3373 20160
rect 3309 20100 3313 20156
rect 3313 20100 3369 20156
rect 3369 20100 3373 20156
rect 3309 20096 3373 20100
rect 3389 20156 3453 20160
rect 3389 20100 3393 20156
rect 3393 20100 3449 20156
rect 3449 20100 3453 20156
rect 3389 20096 3453 20100
rect 3469 20156 3533 20160
rect 3469 20100 3473 20156
rect 3473 20100 3529 20156
rect 3529 20100 3533 20156
rect 3469 20096 3533 20100
rect 3549 20156 3613 20160
rect 3549 20100 3553 20156
rect 3553 20100 3609 20156
rect 3609 20100 3613 20156
rect 3549 20096 3613 20100
rect 4252 20156 4316 20160
rect 4252 20100 4256 20156
rect 4256 20100 4312 20156
rect 4312 20100 4316 20156
rect 4252 20096 4316 20100
rect 4332 20156 4396 20160
rect 4332 20100 4336 20156
rect 4336 20100 4392 20156
rect 4392 20100 4396 20156
rect 4332 20096 4396 20100
rect 4412 20156 4476 20160
rect 4412 20100 4416 20156
rect 4416 20100 4472 20156
rect 4472 20100 4476 20156
rect 4412 20096 4476 20100
rect 4492 20156 4556 20160
rect 4492 20100 4496 20156
rect 4496 20100 4552 20156
rect 4552 20100 4556 20156
rect 4492 20096 4556 20100
rect 1894 19612 1958 19616
rect 1894 19556 1898 19612
rect 1898 19556 1954 19612
rect 1954 19556 1958 19612
rect 1894 19552 1958 19556
rect 1974 19612 2038 19616
rect 1974 19556 1978 19612
rect 1978 19556 2034 19612
rect 2034 19556 2038 19612
rect 1974 19552 2038 19556
rect 2054 19612 2118 19616
rect 2054 19556 2058 19612
rect 2058 19556 2114 19612
rect 2114 19556 2118 19612
rect 2054 19552 2118 19556
rect 2134 19612 2198 19616
rect 2134 19556 2138 19612
rect 2138 19556 2194 19612
rect 2194 19556 2198 19612
rect 2134 19552 2198 19556
rect 2837 19612 2901 19616
rect 2837 19556 2841 19612
rect 2841 19556 2897 19612
rect 2897 19556 2901 19612
rect 2837 19552 2901 19556
rect 2917 19612 2981 19616
rect 2917 19556 2921 19612
rect 2921 19556 2977 19612
rect 2977 19556 2981 19612
rect 2917 19552 2981 19556
rect 2997 19612 3061 19616
rect 2997 19556 3001 19612
rect 3001 19556 3057 19612
rect 3057 19556 3061 19612
rect 2997 19552 3061 19556
rect 3077 19612 3141 19616
rect 3077 19556 3081 19612
rect 3081 19556 3137 19612
rect 3137 19556 3141 19612
rect 3077 19552 3141 19556
rect 3780 19612 3844 19616
rect 3780 19556 3784 19612
rect 3784 19556 3840 19612
rect 3840 19556 3844 19612
rect 3780 19552 3844 19556
rect 3860 19612 3924 19616
rect 3860 19556 3864 19612
rect 3864 19556 3920 19612
rect 3920 19556 3924 19612
rect 3860 19552 3924 19556
rect 3940 19612 4004 19616
rect 3940 19556 3944 19612
rect 3944 19556 4000 19612
rect 4000 19556 4004 19612
rect 3940 19552 4004 19556
rect 4020 19612 4084 19616
rect 4020 19556 4024 19612
rect 4024 19556 4080 19612
rect 4080 19556 4084 19612
rect 4020 19552 4084 19556
rect 4723 19612 4787 19616
rect 4723 19556 4727 19612
rect 4727 19556 4783 19612
rect 4783 19556 4787 19612
rect 4723 19552 4787 19556
rect 4803 19612 4867 19616
rect 4803 19556 4807 19612
rect 4807 19556 4863 19612
rect 4863 19556 4867 19612
rect 4803 19552 4867 19556
rect 4883 19612 4947 19616
rect 4883 19556 4887 19612
rect 4887 19556 4943 19612
rect 4943 19556 4947 19612
rect 4883 19552 4947 19556
rect 4963 19612 5027 19616
rect 4963 19556 4967 19612
rect 4967 19556 5023 19612
rect 5023 19556 5027 19612
rect 4963 19552 5027 19556
rect 1423 19068 1487 19072
rect 1423 19012 1427 19068
rect 1427 19012 1483 19068
rect 1483 19012 1487 19068
rect 1423 19008 1487 19012
rect 1503 19068 1567 19072
rect 1503 19012 1507 19068
rect 1507 19012 1563 19068
rect 1563 19012 1567 19068
rect 1503 19008 1567 19012
rect 1583 19068 1647 19072
rect 1583 19012 1587 19068
rect 1587 19012 1643 19068
rect 1643 19012 1647 19068
rect 1583 19008 1647 19012
rect 1663 19068 1727 19072
rect 1663 19012 1667 19068
rect 1667 19012 1723 19068
rect 1723 19012 1727 19068
rect 1663 19008 1727 19012
rect 2366 19068 2430 19072
rect 2366 19012 2370 19068
rect 2370 19012 2426 19068
rect 2426 19012 2430 19068
rect 2366 19008 2430 19012
rect 2446 19068 2510 19072
rect 2446 19012 2450 19068
rect 2450 19012 2506 19068
rect 2506 19012 2510 19068
rect 2446 19008 2510 19012
rect 2526 19068 2590 19072
rect 2526 19012 2530 19068
rect 2530 19012 2586 19068
rect 2586 19012 2590 19068
rect 2526 19008 2590 19012
rect 2606 19068 2670 19072
rect 2606 19012 2610 19068
rect 2610 19012 2666 19068
rect 2666 19012 2670 19068
rect 2606 19008 2670 19012
rect 3309 19068 3373 19072
rect 3309 19012 3313 19068
rect 3313 19012 3369 19068
rect 3369 19012 3373 19068
rect 3309 19008 3373 19012
rect 3389 19068 3453 19072
rect 3389 19012 3393 19068
rect 3393 19012 3449 19068
rect 3449 19012 3453 19068
rect 3389 19008 3453 19012
rect 3469 19068 3533 19072
rect 3469 19012 3473 19068
rect 3473 19012 3529 19068
rect 3529 19012 3533 19068
rect 3469 19008 3533 19012
rect 3549 19068 3613 19072
rect 3549 19012 3553 19068
rect 3553 19012 3609 19068
rect 3609 19012 3613 19068
rect 3549 19008 3613 19012
rect 4252 19068 4316 19072
rect 4252 19012 4256 19068
rect 4256 19012 4312 19068
rect 4312 19012 4316 19068
rect 4252 19008 4316 19012
rect 4332 19068 4396 19072
rect 4332 19012 4336 19068
rect 4336 19012 4392 19068
rect 4392 19012 4396 19068
rect 4332 19008 4396 19012
rect 4412 19068 4476 19072
rect 4412 19012 4416 19068
rect 4416 19012 4472 19068
rect 4472 19012 4476 19068
rect 4412 19008 4476 19012
rect 4492 19068 4556 19072
rect 4492 19012 4496 19068
rect 4496 19012 4552 19068
rect 4552 19012 4556 19068
rect 4492 19008 4556 19012
rect 1894 18524 1958 18528
rect 1894 18468 1898 18524
rect 1898 18468 1954 18524
rect 1954 18468 1958 18524
rect 1894 18464 1958 18468
rect 1974 18524 2038 18528
rect 1974 18468 1978 18524
rect 1978 18468 2034 18524
rect 2034 18468 2038 18524
rect 1974 18464 2038 18468
rect 2054 18524 2118 18528
rect 2054 18468 2058 18524
rect 2058 18468 2114 18524
rect 2114 18468 2118 18524
rect 2054 18464 2118 18468
rect 2134 18524 2198 18528
rect 2134 18468 2138 18524
rect 2138 18468 2194 18524
rect 2194 18468 2198 18524
rect 2134 18464 2198 18468
rect 2837 18524 2901 18528
rect 2837 18468 2841 18524
rect 2841 18468 2897 18524
rect 2897 18468 2901 18524
rect 2837 18464 2901 18468
rect 2917 18524 2981 18528
rect 2917 18468 2921 18524
rect 2921 18468 2977 18524
rect 2977 18468 2981 18524
rect 2917 18464 2981 18468
rect 2997 18524 3061 18528
rect 2997 18468 3001 18524
rect 3001 18468 3057 18524
rect 3057 18468 3061 18524
rect 2997 18464 3061 18468
rect 3077 18524 3141 18528
rect 3077 18468 3081 18524
rect 3081 18468 3137 18524
rect 3137 18468 3141 18524
rect 3077 18464 3141 18468
rect 3780 18524 3844 18528
rect 3780 18468 3784 18524
rect 3784 18468 3840 18524
rect 3840 18468 3844 18524
rect 3780 18464 3844 18468
rect 3860 18524 3924 18528
rect 3860 18468 3864 18524
rect 3864 18468 3920 18524
rect 3920 18468 3924 18524
rect 3860 18464 3924 18468
rect 3940 18524 4004 18528
rect 3940 18468 3944 18524
rect 3944 18468 4000 18524
rect 4000 18468 4004 18524
rect 3940 18464 4004 18468
rect 4020 18524 4084 18528
rect 4020 18468 4024 18524
rect 4024 18468 4080 18524
rect 4080 18468 4084 18524
rect 4020 18464 4084 18468
rect 4723 18524 4787 18528
rect 4723 18468 4727 18524
rect 4727 18468 4783 18524
rect 4783 18468 4787 18524
rect 4723 18464 4787 18468
rect 4803 18524 4867 18528
rect 4803 18468 4807 18524
rect 4807 18468 4863 18524
rect 4863 18468 4867 18524
rect 4803 18464 4867 18468
rect 4883 18524 4947 18528
rect 4883 18468 4887 18524
rect 4887 18468 4943 18524
rect 4943 18468 4947 18524
rect 4883 18464 4947 18468
rect 4963 18524 5027 18528
rect 4963 18468 4967 18524
rect 4967 18468 5023 18524
rect 5023 18468 5027 18524
rect 4963 18464 5027 18468
rect 1423 17980 1487 17984
rect 1423 17924 1427 17980
rect 1427 17924 1483 17980
rect 1483 17924 1487 17980
rect 1423 17920 1487 17924
rect 1503 17980 1567 17984
rect 1503 17924 1507 17980
rect 1507 17924 1563 17980
rect 1563 17924 1567 17980
rect 1503 17920 1567 17924
rect 1583 17980 1647 17984
rect 1583 17924 1587 17980
rect 1587 17924 1643 17980
rect 1643 17924 1647 17980
rect 1583 17920 1647 17924
rect 1663 17980 1727 17984
rect 1663 17924 1667 17980
rect 1667 17924 1723 17980
rect 1723 17924 1727 17980
rect 1663 17920 1727 17924
rect 2366 17980 2430 17984
rect 2366 17924 2370 17980
rect 2370 17924 2426 17980
rect 2426 17924 2430 17980
rect 2366 17920 2430 17924
rect 2446 17980 2510 17984
rect 2446 17924 2450 17980
rect 2450 17924 2506 17980
rect 2506 17924 2510 17980
rect 2446 17920 2510 17924
rect 2526 17980 2590 17984
rect 2526 17924 2530 17980
rect 2530 17924 2586 17980
rect 2586 17924 2590 17980
rect 2526 17920 2590 17924
rect 2606 17980 2670 17984
rect 2606 17924 2610 17980
rect 2610 17924 2666 17980
rect 2666 17924 2670 17980
rect 2606 17920 2670 17924
rect 3309 17980 3373 17984
rect 3309 17924 3313 17980
rect 3313 17924 3369 17980
rect 3369 17924 3373 17980
rect 3309 17920 3373 17924
rect 3389 17980 3453 17984
rect 3389 17924 3393 17980
rect 3393 17924 3449 17980
rect 3449 17924 3453 17980
rect 3389 17920 3453 17924
rect 3469 17980 3533 17984
rect 3469 17924 3473 17980
rect 3473 17924 3529 17980
rect 3529 17924 3533 17980
rect 3469 17920 3533 17924
rect 3549 17980 3613 17984
rect 3549 17924 3553 17980
rect 3553 17924 3609 17980
rect 3609 17924 3613 17980
rect 3549 17920 3613 17924
rect 4252 17980 4316 17984
rect 4252 17924 4256 17980
rect 4256 17924 4312 17980
rect 4312 17924 4316 17980
rect 4252 17920 4316 17924
rect 4332 17980 4396 17984
rect 4332 17924 4336 17980
rect 4336 17924 4392 17980
rect 4392 17924 4396 17980
rect 4332 17920 4396 17924
rect 4412 17980 4476 17984
rect 4412 17924 4416 17980
rect 4416 17924 4472 17980
rect 4472 17924 4476 17980
rect 4412 17920 4476 17924
rect 4492 17980 4556 17984
rect 4492 17924 4496 17980
rect 4496 17924 4552 17980
rect 4552 17924 4556 17980
rect 4492 17920 4556 17924
rect 1894 17436 1958 17440
rect 1894 17380 1898 17436
rect 1898 17380 1954 17436
rect 1954 17380 1958 17436
rect 1894 17376 1958 17380
rect 1974 17436 2038 17440
rect 1974 17380 1978 17436
rect 1978 17380 2034 17436
rect 2034 17380 2038 17436
rect 1974 17376 2038 17380
rect 2054 17436 2118 17440
rect 2054 17380 2058 17436
rect 2058 17380 2114 17436
rect 2114 17380 2118 17436
rect 2054 17376 2118 17380
rect 2134 17436 2198 17440
rect 2134 17380 2138 17436
rect 2138 17380 2194 17436
rect 2194 17380 2198 17436
rect 2134 17376 2198 17380
rect 2837 17436 2901 17440
rect 2837 17380 2841 17436
rect 2841 17380 2897 17436
rect 2897 17380 2901 17436
rect 2837 17376 2901 17380
rect 2917 17436 2981 17440
rect 2917 17380 2921 17436
rect 2921 17380 2977 17436
rect 2977 17380 2981 17436
rect 2917 17376 2981 17380
rect 2997 17436 3061 17440
rect 2997 17380 3001 17436
rect 3001 17380 3057 17436
rect 3057 17380 3061 17436
rect 2997 17376 3061 17380
rect 3077 17436 3141 17440
rect 3077 17380 3081 17436
rect 3081 17380 3137 17436
rect 3137 17380 3141 17436
rect 3077 17376 3141 17380
rect 3780 17436 3844 17440
rect 3780 17380 3784 17436
rect 3784 17380 3840 17436
rect 3840 17380 3844 17436
rect 3780 17376 3844 17380
rect 3860 17436 3924 17440
rect 3860 17380 3864 17436
rect 3864 17380 3920 17436
rect 3920 17380 3924 17436
rect 3860 17376 3924 17380
rect 3940 17436 4004 17440
rect 3940 17380 3944 17436
rect 3944 17380 4000 17436
rect 4000 17380 4004 17436
rect 3940 17376 4004 17380
rect 4020 17436 4084 17440
rect 4020 17380 4024 17436
rect 4024 17380 4080 17436
rect 4080 17380 4084 17436
rect 4020 17376 4084 17380
rect 4723 17436 4787 17440
rect 4723 17380 4727 17436
rect 4727 17380 4783 17436
rect 4783 17380 4787 17436
rect 4723 17376 4787 17380
rect 4803 17436 4867 17440
rect 4803 17380 4807 17436
rect 4807 17380 4863 17436
rect 4863 17380 4867 17436
rect 4803 17376 4867 17380
rect 4883 17436 4947 17440
rect 4883 17380 4887 17436
rect 4887 17380 4943 17436
rect 4943 17380 4947 17436
rect 4883 17376 4947 17380
rect 4963 17436 5027 17440
rect 4963 17380 4967 17436
rect 4967 17380 5023 17436
rect 5023 17380 5027 17436
rect 4963 17376 5027 17380
rect 1423 16892 1487 16896
rect 1423 16836 1427 16892
rect 1427 16836 1483 16892
rect 1483 16836 1487 16892
rect 1423 16832 1487 16836
rect 1503 16892 1567 16896
rect 1503 16836 1507 16892
rect 1507 16836 1563 16892
rect 1563 16836 1567 16892
rect 1503 16832 1567 16836
rect 1583 16892 1647 16896
rect 1583 16836 1587 16892
rect 1587 16836 1643 16892
rect 1643 16836 1647 16892
rect 1583 16832 1647 16836
rect 1663 16892 1727 16896
rect 1663 16836 1667 16892
rect 1667 16836 1723 16892
rect 1723 16836 1727 16892
rect 1663 16832 1727 16836
rect 2366 16892 2430 16896
rect 2366 16836 2370 16892
rect 2370 16836 2426 16892
rect 2426 16836 2430 16892
rect 2366 16832 2430 16836
rect 2446 16892 2510 16896
rect 2446 16836 2450 16892
rect 2450 16836 2506 16892
rect 2506 16836 2510 16892
rect 2446 16832 2510 16836
rect 2526 16892 2590 16896
rect 2526 16836 2530 16892
rect 2530 16836 2586 16892
rect 2586 16836 2590 16892
rect 2526 16832 2590 16836
rect 2606 16892 2670 16896
rect 2606 16836 2610 16892
rect 2610 16836 2666 16892
rect 2666 16836 2670 16892
rect 2606 16832 2670 16836
rect 3309 16892 3373 16896
rect 3309 16836 3313 16892
rect 3313 16836 3369 16892
rect 3369 16836 3373 16892
rect 3309 16832 3373 16836
rect 3389 16892 3453 16896
rect 3389 16836 3393 16892
rect 3393 16836 3449 16892
rect 3449 16836 3453 16892
rect 3389 16832 3453 16836
rect 3469 16892 3533 16896
rect 3469 16836 3473 16892
rect 3473 16836 3529 16892
rect 3529 16836 3533 16892
rect 3469 16832 3533 16836
rect 3549 16892 3613 16896
rect 3549 16836 3553 16892
rect 3553 16836 3609 16892
rect 3609 16836 3613 16892
rect 3549 16832 3613 16836
rect 4252 16892 4316 16896
rect 4252 16836 4256 16892
rect 4256 16836 4312 16892
rect 4312 16836 4316 16892
rect 4252 16832 4316 16836
rect 4332 16892 4396 16896
rect 4332 16836 4336 16892
rect 4336 16836 4392 16892
rect 4392 16836 4396 16892
rect 4332 16832 4396 16836
rect 4412 16892 4476 16896
rect 4412 16836 4416 16892
rect 4416 16836 4472 16892
rect 4472 16836 4476 16892
rect 4412 16832 4476 16836
rect 4492 16892 4556 16896
rect 4492 16836 4496 16892
rect 4496 16836 4552 16892
rect 4552 16836 4556 16892
rect 4492 16832 4556 16836
rect 1894 16348 1958 16352
rect 1894 16292 1898 16348
rect 1898 16292 1954 16348
rect 1954 16292 1958 16348
rect 1894 16288 1958 16292
rect 1974 16348 2038 16352
rect 1974 16292 1978 16348
rect 1978 16292 2034 16348
rect 2034 16292 2038 16348
rect 1974 16288 2038 16292
rect 2054 16348 2118 16352
rect 2054 16292 2058 16348
rect 2058 16292 2114 16348
rect 2114 16292 2118 16348
rect 2054 16288 2118 16292
rect 2134 16348 2198 16352
rect 2134 16292 2138 16348
rect 2138 16292 2194 16348
rect 2194 16292 2198 16348
rect 2134 16288 2198 16292
rect 2837 16348 2901 16352
rect 2837 16292 2841 16348
rect 2841 16292 2897 16348
rect 2897 16292 2901 16348
rect 2837 16288 2901 16292
rect 2917 16348 2981 16352
rect 2917 16292 2921 16348
rect 2921 16292 2977 16348
rect 2977 16292 2981 16348
rect 2917 16288 2981 16292
rect 2997 16348 3061 16352
rect 2997 16292 3001 16348
rect 3001 16292 3057 16348
rect 3057 16292 3061 16348
rect 2997 16288 3061 16292
rect 3077 16348 3141 16352
rect 3077 16292 3081 16348
rect 3081 16292 3137 16348
rect 3137 16292 3141 16348
rect 3077 16288 3141 16292
rect 3780 16348 3844 16352
rect 3780 16292 3784 16348
rect 3784 16292 3840 16348
rect 3840 16292 3844 16348
rect 3780 16288 3844 16292
rect 3860 16348 3924 16352
rect 3860 16292 3864 16348
rect 3864 16292 3920 16348
rect 3920 16292 3924 16348
rect 3860 16288 3924 16292
rect 3940 16348 4004 16352
rect 3940 16292 3944 16348
rect 3944 16292 4000 16348
rect 4000 16292 4004 16348
rect 3940 16288 4004 16292
rect 4020 16348 4084 16352
rect 4020 16292 4024 16348
rect 4024 16292 4080 16348
rect 4080 16292 4084 16348
rect 4020 16288 4084 16292
rect 4723 16348 4787 16352
rect 4723 16292 4727 16348
rect 4727 16292 4783 16348
rect 4783 16292 4787 16348
rect 4723 16288 4787 16292
rect 4803 16348 4867 16352
rect 4803 16292 4807 16348
rect 4807 16292 4863 16348
rect 4863 16292 4867 16348
rect 4803 16288 4867 16292
rect 4883 16348 4947 16352
rect 4883 16292 4887 16348
rect 4887 16292 4943 16348
rect 4943 16292 4947 16348
rect 4883 16288 4947 16292
rect 4963 16348 5027 16352
rect 4963 16292 4967 16348
rect 4967 16292 5023 16348
rect 5023 16292 5027 16348
rect 4963 16288 5027 16292
rect 1423 15804 1487 15808
rect 1423 15748 1427 15804
rect 1427 15748 1483 15804
rect 1483 15748 1487 15804
rect 1423 15744 1487 15748
rect 1503 15804 1567 15808
rect 1503 15748 1507 15804
rect 1507 15748 1563 15804
rect 1563 15748 1567 15804
rect 1503 15744 1567 15748
rect 1583 15804 1647 15808
rect 1583 15748 1587 15804
rect 1587 15748 1643 15804
rect 1643 15748 1647 15804
rect 1583 15744 1647 15748
rect 1663 15804 1727 15808
rect 1663 15748 1667 15804
rect 1667 15748 1723 15804
rect 1723 15748 1727 15804
rect 1663 15744 1727 15748
rect 2366 15804 2430 15808
rect 2366 15748 2370 15804
rect 2370 15748 2426 15804
rect 2426 15748 2430 15804
rect 2366 15744 2430 15748
rect 2446 15804 2510 15808
rect 2446 15748 2450 15804
rect 2450 15748 2506 15804
rect 2506 15748 2510 15804
rect 2446 15744 2510 15748
rect 2526 15804 2590 15808
rect 2526 15748 2530 15804
rect 2530 15748 2586 15804
rect 2586 15748 2590 15804
rect 2526 15744 2590 15748
rect 2606 15804 2670 15808
rect 2606 15748 2610 15804
rect 2610 15748 2666 15804
rect 2666 15748 2670 15804
rect 2606 15744 2670 15748
rect 3309 15804 3373 15808
rect 3309 15748 3313 15804
rect 3313 15748 3369 15804
rect 3369 15748 3373 15804
rect 3309 15744 3373 15748
rect 3389 15804 3453 15808
rect 3389 15748 3393 15804
rect 3393 15748 3449 15804
rect 3449 15748 3453 15804
rect 3389 15744 3453 15748
rect 3469 15804 3533 15808
rect 3469 15748 3473 15804
rect 3473 15748 3529 15804
rect 3529 15748 3533 15804
rect 3469 15744 3533 15748
rect 3549 15804 3613 15808
rect 3549 15748 3553 15804
rect 3553 15748 3609 15804
rect 3609 15748 3613 15804
rect 3549 15744 3613 15748
rect 4252 15804 4316 15808
rect 4252 15748 4256 15804
rect 4256 15748 4312 15804
rect 4312 15748 4316 15804
rect 4252 15744 4316 15748
rect 4332 15804 4396 15808
rect 4332 15748 4336 15804
rect 4336 15748 4392 15804
rect 4392 15748 4396 15804
rect 4332 15744 4396 15748
rect 4412 15804 4476 15808
rect 4412 15748 4416 15804
rect 4416 15748 4472 15804
rect 4472 15748 4476 15804
rect 4412 15744 4476 15748
rect 4492 15804 4556 15808
rect 4492 15748 4496 15804
rect 4496 15748 4552 15804
rect 4552 15748 4556 15804
rect 4492 15744 4556 15748
rect 1894 15260 1958 15264
rect 1894 15204 1898 15260
rect 1898 15204 1954 15260
rect 1954 15204 1958 15260
rect 1894 15200 1958 15204
rect 1974 15260 2038 15264
rect 1974 15204 1978 15260
rect 1978 15204 2034 15260
rect 2034 15204 2038 15260
rect 1974 15200 2038 15204
rect 2054 15260 2118 15264
rect 2054 15204 2058 15260
rect 2058 15204 2114 15260
rect 2114 15204 2118 15260
rect 2054 15200 2118 15204
rect 2134 15260 2198 15264
rect 2134 15204 2138 15260
rect 2138 15204 2194 15260
rect 2194 15204 2198 15260
rect 2134 15200 2198 15204
rect 2837 15260 2901 15264
rect 2837 15204 2841 15260
rect 2841 15204 2897 15260
rect 2897 15204 2901 15260
rect 2837 15200 2901 15204
rect 2917 15260 2981 15264
rect 2917 15204 2921 15260
rect 2921 15204 2977 15260
rect 2977 15204 2981 15260
rect 2917 15200 2981 15204
rect 2997 15260 3061 15264
rect 2997 15204 3001 15260
rect 3001 15204 3057 15260
rect 3057 15204 3061 15260
rect 2997 15200 3061 15204
rect 3077 15260 3141 15264
rect 3077 15204 3081 15260
rect 3081 15204 3137 15260
rect 3137 15204 3141 15260
rect 3077 15200 3141 15204
rect 3780 15260 3844 15264
rect 3780 15204 3784 15260
rect 3784 15204 3840 15260
rect 3840 15204 3844 15260
rect 3780 15200 3844 15204
rect 3860 15260 3924 15264
rect 3860 15204 3864 15260
rect 3864 15204 3920 15260
rect 3920 15204 3924 15260
rect 3860 15200 3924 15204
rect 3940 15260 4004 15264
rect 3940 15204 3944 15260
rect 3944 15204 4000 15260
rect 4000 15204 4004 15260
rect 3940 15200 4004 15204
rect 4020 15260 4084 15264
rect 4020 15204 4024 15260
rect 4024 15204 4080 15260
rect 4080 15204 4084 15260
rect 4020 15200 4084 15204
rect 4723 15260 4787 15264
rect 4723 15204 4727 15260
rect 4727 15204 4783 15260
rect 4783 15204 4787 15260
rect 4723 15200 4787 15204
rect 4803 15260 4867 15264
rect 4803 15204 4807 15260
rect 4807 15204 4863 15260
rect 4863 15204 4867 15260
rect 4803 15200 4867 15204
rect 4883 15260 4947 15264
rect 4883 15204 4887 15260
rect 4887 15204 4943 15260
rect 4943 15204 4947 15260
rect 4883 15200 4947 15204
rect 4963 15260 5027 15264
rect 4963 15204 4967 15260
rect 4967 15204 5023 15260
rect 5023 15204 5027 15260
rect 4963 15200 5027 15204
rect 1423 14716 1487 14720
rect 1423 14660 1427 14716
rect 1427 14660 1483 14716
rect 1483 14660 1487 14716
rect 1423 14656 1487 14660
rect 1503 14716 1567 14720
rect 1503 14660 1507 14716
rect 1507 14660 1563 14716
rect 1563 14660 1567 14716
rect 1503 14656 1567 14660
rect 1583 14716 1647 14720
rect 1583 14660 1587 14716
rect 1587 14660 1643 14716
rect 1643 14660 1647 14716
rect 1583 14656 1647 14660
rect 1663 14716 1727 14720
rect 1663 14660 1667 14716
rect 1667 14660 1723 14716
rect 1723 14660 1727 14716
rect 1663 14656 1727 14660
rect 2366 14716 2430 14720
rect 2366 14660 2370 14716
rect 2370 14660 2426 14716
rect 2426 14660 2430 14716
rect 2366 14656 2430 14660
rect 2446 14716 2510 14720
rect 2446 14660 2450 14716
rect 2450 14660 2506 14716
rect 2506 14660 2510 14716
rect 2446 14656 2510 14660
rect 2526 14716 2590 14720
rect 2526 14660 2530 14716
rect 2530 14660 2586 14716
rect 2586 14660 2590 14716
rect 2526 14656 2590 14660
rect 2606 14716 2670 14720
rect 2606 14660 2610 14716
rect 2610 14660 2666 14716
rect 2666 14660 2670 14716
rect 2606 14656 2670 14660
rect 3309 14716 3373 14720
rect 3309 14660 3313 14716
rect 3313 14660 3369 14716
rect 3369 14660 3373 14716
rect 3309 14656 3373 14660
rect 3389 14716 3453 14720
rect 3389 14660 3393 14716
rect 3393 14660 3449 14716
rect 3449 14660 3453 14716
rect 3389 14656 3453 14660
rect 3469 14716 3533 14720
rect 3469 14660 3473 14716
rect 3473 14660 3529 14716
rect 3529 14660 3533 14716
rect 3469 14656 3533 14660
rect 3549 14716 3613 14720
rect 3549 14660 3553 14716
rect 3553 14660 3609 14716
rect 3609 14660 3613 14716
rect 3549 14656 3613 14660
rect 4252 14716 4316 14720
rect 4252 14660 4256 14716
rect 4256 14660 4312 14716
rect 4312 14660 4316 14716
rect 4252 14656 4316 14660
rect 4332 14716 4396 14720
rect 4332 14660 4336 14716
rect 4336 14660 4392 14716
rect 4392 14660 4396 14716
rect 4332 14656 4396 14660
rect 4412 14716 4476 14720
rect 4412 14660 4416 14716
rect 4416 14660 4472 14716
rect 4472 14660 4476 14716
rect 4412 14656 4476 14660
rect 4492 14716 4556 14720
rect 4492 14660 4496 14716
rect 4496 14660 4552 14716
rect 4552 14660 4556 14716
rect 4492 14656 4556 14660
rect 1894 14172 1958 14176
rect 1894 14116 1898 14172
rect 1898 14116 1954 14172
rect 1954 14116 1958 14172
rect 1894 14112 1958 14116
rect 1974 14172 2038 14176
rect 1974 14116 1978 14172
rect 1978 14116 2034 14172
rect 2034 14116 2038 14172
rect 1974 14112 2038 14116
rect 2054 14172 2118 14176
rect 2054 14116 2058 14172
rect 2058 14116 2114 14172
rect 2114 14116 2118 14172
rect 2054 14112 2118 14116
rect 2134 14172 2198 14176
rect 2134 14116 2138 14172
rect 2138 14116 2194 14172
rect 2194 14116 2198 14172
rect 2134 14112 2198 14116
rect 2837 14172 2901 14176
rect 2837 14116 2841 14172
rect 2841 14116 2897 14172
rect 2897 14116 2901 14172
rect 2837 14112 2901 14116
rect 2917 14172 2981 14176
rect 2917 14116 2921 14172
rect 2921 14116 2977 14172
rect 2977 14116 2981 14172
rect 2917 14112 2981 14116
rect 2997 14172 3061 14176
rect 2997 14116 3001 14172
rect 3001 14116 3057 14172
rect 3057 14116 3061 14172
rect 2997 14112 3061 14116
rect 3077 14172 3141 14176
rect 3077 14116 3081 14172
rect 3081 14116 3137 14172
rect 3137 14116 3141 14172
rect 3077 14112 3141 14116
rect 3780 14172 3844 14176
rect 3780 14116 3784 14172
rect 3784 14116 3840 14172
rect 3840 14116 3844 14172
rect 3780 14112 3844 14116
rect 3860 14172 3924 14176
rect 3860 14116 3864 14172
rect 3864 14116 3920 14172
rect 3920 14116 3924 14172
rect 3860 14112 3924 14116
rect 3940 14172 4004 14176
rect 3940 14116 3944 14172
rect 3944 14116 4000 14172
rect 4000 14116 4004 14172
rect 3940 14112 4004 14116
rect 4020 14172 4084 14176
rect 4020 14116 4024 14172
rect 4024 14116 4080 14172
rect 4080 14116 4084 14172
rect 4020 14112 4084 14116
rect 4723 14172 4787 14176
rect 4723 14116 4727 14172
rect 4727 14116 4783 14172
rect 4783 14116 4787 14172
rect 4723 14112 4787 14116
rect 4803 14172 4867 14176
rect 4803 14116 4807 14172
rect 4807 14116 4863 14172
rect 4863 14116 4867 14172
rect 4803 14112 4867 14116
rect 4883 14172 4947 14176
rect 4883 14116 4887 14172
rect 4887 14116 4943 14172
rect 4943 14116 4947 14172
rect 4883 14112 4947 14116
rect 4963 14172 5027 14176
rect 4963 14116 4967 14172
rect 4967 14116 5023 14172
rect 5023 14116 5027 14172
rect 4963 14112 5027 14116
rect 1423 13628 1487 13632
rect 1423 13572 1427 13628
rect 1427 13572 1483 13628
rect 1483 13572 1487 13628
rect 1423 13568 1487 13572
rect 1503 13628 1567 13632
rect 1503 13572 1507 13628
rect 1507 13572 1563 13628
rect 1563 13572 1567 13628
rect 1503 13568 1567 13572
rect 1583 13628 1647 13632
rect 1583 13572 1587 13628
rect 1587 13572 1643 13628
rect 1643 13572 1647 13628
rect 1583 13568 1647 13572
rect 1663 13628 1727 13632
rect 1663 13572 1667 13628
rect 1667 13572 1723 13628
rect 1723 13572 1727 13628
rect 1663 13568 1727 13572
rect 2366 13628 2430 13632
rect 2366 13572 2370 13628
rect 2370 13572 2426 13628
rect 2426 13572 2430 13628
rect 2366 13568 2430 13572
rect 2446 13628 2510 13632
rect 2446 13572 2450 13628
rect 2450 13572 2506 13628
rect 2506 13572 2510 13628
rect 2446 13568 2510 13572
rect 2526 13628 2590 13632
rect 2526 13572 2530 13628
rect 2530 13572 2586 13628
rect 2586 13572 2590 13628
rect 2526 13568 2590 13572
rect 2606 13628 2670 13632
rect 2606 13572 2610 13628
rect 2610 13572 2666 13628
rect 2666 13572 2670 13628
rect 2606 13568 2670 13572
rect 3309 13628 3373 13632
rect 3309 13572 3313 13628
rect 3313 13572 3369 13628
rect 3369 13572 3373 13628
rect 3309 13568 3373 13572
rect 3389 13628 3453 13632
rect 3389 13572 3393 13628
rect 3393 13572 3449 13628
rect 3449 13572 3453 13628
rect 3389 13568 3453 13572
rect 3469 13628 3533 13632
rect 3469 13572 3473 13628
rect 3473 13572 3529 13628
rect 3529 13572 3533 13628
rect 3469 13568 3533 13572
rect 3549 13628 3613 13632
rect 3549 13572 3553 13628
rect 3553 13572 3609 13628
rect 3609 13572 3613 13628
rect 3549 13568 3613 13572
rect 4252 13628 4316 13632
rect 4252 13572 4256 13628
rect 4256 13572 4312 13628
rect 4312 13572 4316 13628
rect 4252 13568 4316 13572
rect 4332 13628 4396 13632
rect 4332 13572 4336 13628
rect 4336 13572 4392 13628
rect 4392 13572 4396 13628
rect 4332 13568 4396 13572
rect 4412 13628 4476 13632
rect 4412 13572 4416 13628
rect 4416 13572 4472 13628
rect 4472 13572 4476 13628
rect 4412 13568 4476 13572
rect 4492 13628 4556 13632
rect 4492 13572 4496 13628
rect 4496 13572 4552 13628
rect 4552 13572 4556 13628
rect 4492 13568 4556 13572
rect 1894 13084 1958 13088
rect 1894 13028 1898 13084
rect 1898 13028 1954 13084
rect 1954 13028 1958 13084
rect 1894 13024 1958 13028
rect 1974 13084 2038 13088
rect 1974 13028 1978 13084
rect 1978 13028 2034 13084
rect 2034 13028 2038 13084
rect 1974 13024 2038 13028
rect 2054 13084 2118 13088
rect 2054 13028 2058 13084
rect 2058 13028 2114 13084
rect 2114 13028 2118 13084
rect 2054 13024 2118 13028
rect 2134 13084 2198 13088
rect 2134 13028 2138 13084
rect 2138 13028 2194 13084
rect 2194 13028 2198 13084
rect 2134 13024 2198 13028
rect 2837 13084 2901 13088
rect 2837 13028 2841 13084
rect 2841 13028 2897 13084
rect 2897 13028 2901 13084
rect 2837 13024 2901 13028
rect 2917 13084 2981 13088
rect 2917 13028 2921 13084
rect 2921 13028 2977 13084
rect 2977 13028 2981 13084
rect 2917 13024 2981 13028
rect 2997 13084 3061 13088
rect 2997 13028 3001 13084
rect 3001 13028 3057 13084
rect 3057 13028 3061 13084
rect 2997 13024 3061 13028
rect 3077 13084 3141 13088
rect 3077 13028 3081 13084
rect 3081 13028 3137 13084
rect 3137 13028 3141 13084
rect 3077 13024 3141 13028
rect 3780 13084 3844 13088
rect 3780 13028 3784 13084
rect 3784 13028 3840 13084
rect 3840 13028 3844 13084
rect 3780 13024 3844 13028
rect 3860 13084 3924 13088
rect 3860 13028 3864 13084
rect 3864 13028 3920 13084
rect 3920 13028 3924 13084
rect 3860 13024 3924 13028
rect 3940 13084 4004 13088
rect 3940 13028 3944 13084
rect 3944 13028 4000 13084
rect 4000 13028 4004 13084
rect 3940 13024 4004 13028
rect 4020 13084 4084 13088
rect 4020 13028 4024 13084
rect 4024 13028 4080 13084
rect 4080 13028 4084 13084
rect 4020 13024 4084 13028
rect 4723 13084 4787 13088
rect 4723 13028 4727 13084
rect 4727 13028 4783 13084
rect 4783 13028 4787 13084
rect 4723 13024 4787 13028
rect 4803 13084 4867 13088
rect 4803 13028 4807 13084
rect 4807 13028 4863 13084
rect 4863 13028 4867 13084
rect 4803 13024 4867 13028
rect 4883 13084 4947 13088
rect 4883 13028 4887 13084
rect 4887 13028 4943 13084
rect 4943 13028 4947 13084
rect 4883 13024 4947 13028
rect 4963 13084 5027 13088
rect 4963 13028 4967 13084
rect 4967 13028 5023 13084
rect 5023 13028 5027 13084
rect 4963 13024 5027 13028
rect 1423 12540 1487 12544
rect 1423 12484 1427 12540
rect 1427 12484 1483 12540
rect 1483 12484 1487 12540
rect 1423 12480 1487 12484
rect 1503 12540 1567 12544
rect 1503 12484 1507 12540
rect 1507 12484 1563 12540
rect 1563 12484 1567 12540
rect 1503 12480 1567 12484
rect 1583 12540 1647 12544
rect 1583 12484 1587 12540
rect 1587 12484 1643 12540
rect 1643 12484 1647 12540
rect 1583 12480 1647 12484
rect 1663 12540 1727 12544
rect 1663 12484 1667 12540
rect 1667 12484 1723 12540
rect 1723 12484 1727 12540
rect 1663 12480 1727 12484
rect 2366 12540 2430 12544
rect 2366 12484 2370 12540
rect 2370 12484 2426 12540
rect 2426 12484 2430 12540
rect 2366 12480 2430 12484
rect 2446 12540 2510 12544
rect 2446 12484 2450 12540
rect 2450 12484 2506 12540
rect 2506 12484 2510 12540
rect 2446 12480 2510 12484
rect 2526 12540 2590 12544
rect 2526 12484 2530 12540
rect 2530 12484 2586 12540
rect 2586 12484 2590 12540
rect 2526 12480 2590 12484
rect 2606 12540 2670 12544
rect 2606 12484 2610 12540
rect 2610 12484 2666 12540
rect 2666 12484 2670 12540
rect 2606 12480 2670 12484
rect 3309 12540 3373 12544
rect 3309 12484 3313 12540
rect 3313 12484 3369 12540
rect 3369 12484 3373 12540
rect 3309 12480 3373 12484
rect 3389 12540 3453 12544
rect 3389 12484 3393 12540
rect 3393 12484 3449 12540
rect 3449 12484 3453 12540
rect 3389 12480 3453 12484
rect 3469 12540 3533 12544
rect 3469 12484 3473 12540
rect 3473 12484 3529 12540
rect 3529 12484 3533 12540
rect 3469 12480 3533 12484
rect 3549 12540 3613 12544
rect 3549 12484 3553 12540
rect 3553 12484 3609 12540
rect 3609 12484 3613 12540
rect 3549 12480 3613 12484
rect 4252 12540 4316 12544
rect 4252 12484 4256 12540
rect 4256 12484 4312 12540
rect 4312 12484 4316 12540
rect 4252 12480 4316 12484
rect 4332 12540 4396 12544
rect 4332 12484 4336 12540
rect 4336 12484 4392 12540
rect 4392 12484 4396 12540
rect 4332 12480 4396 12484
rect 4412 12540 4476 12544
rect 4412 12484 4416 12540
rect 4416 12484 4472 12540
rect 4472 12484 4476 12540
rect 4412 12480 4476 12484
rect 4492 12540 4556 12544
rect 4492 12484 4496 12540
rect 4496 12484 4552 12540
rect 4552 12484 4556 12540
rect 4492 12480 4556 12484
rect 1894 11996 1958 12000
rect 1894 11940 1898 11996
rect 1898 11940 1954 11996
rect 1954 11940 1958 11996
rect 1894 11936 1958 11940
rect 1974 11996 2038 12000
rect 1974 11940 1978 11996
rect 1978 11940 2034 11996
rect 2034 11940 2038 11996
rect 1974 11936 2038 11940
rect 2054 11996 2118 12000
rect 2054 11940 2058 11996
rect 2058 11940 2114 11996
rect 2114 11940 2118 11996
rect 2054 11936 2118 11940
rect 2134 11996 2198 12000
rect 2134 11940 2138 11996
rect 2138 11940 2194 11996
rect 2194 11940 2198 11996
rect 2134 11936 2198 11940
rect 2837 11996 2901 12000
rect 2837 11940 2841 11996
rect 2841 11940 2897 11996
rect 2897 11940 2901 11996
rect 2837 11936 2901 11940
rect 2917 11996 2981 12000
rect 2917 11940 2921 11996
rect 2921 11940 2977 11996
rect 2977 11940 2981 11996
rect 2917 11936 2981 11940
rect 2997 11996 3061 12000
rect 2997 11940 3001 11996
rect 3001 11940 3057 11996
rect 3057 11940 3061 11996
rect 2997 11936 3061 11940
rect 3077 11996 3141 12000
rect 3077 11940 3081 11996
rect 3081 11940 3137 11996
rect 3137 11940 3141 11996
rect 3077 11936 3141 11940
rect 3780 11996 3844 12000
rect 3780 11940 3784 11996
rect 3784 11940 3840 11996
rect 3840 11940 3844 11996
rect 3780 11936 3844 11940
rect 3860 11996 3924 12000
rect 3860 11940 3864 11996
rect 3864 11940 3920 11996
rect 3920 11940 3924 11996
rect 3860 11936 3924 11940
rect 3940 11996 4004 12000
rect 3940 11940 3944 11996
rect 3944 11940 4000 11996
rect 4000 11940 4004 11996
rect 3940 11936 4004 11940
rect 4020 11996 4084 12000
rect 4020 11940 4024 11996
rect 4024 11940 4080 11996
rect 4080 11940 4084 11996
rect 4020 11936 4084 11940
rect 4723 11996 4787 12000
rect 4723 11940 4727 11996
rect 4727 11940 4783 11996
rect 4783 11940 4787 11996
rect 4723 11936 4787 11940
rect 4803 11996 4867 12000
rect 4803 11940 4807 11996
rect 4807 11940 4863 11996
rect 4863 11940 4867 11996
rect 4803 11936 4867 11940
rect 4883 11996 4947 12000
rect 4883 11940 4887 11996
rect 4887 11940 4943 11996
rect 4943 11940 4947 11996
rect 4883 11936 4947 11940
rect 4963 11996 5027 12000
rect 4963 11940 4967 11996
rect 4967 11940 5023 11996
rect 5023 11940 5027 11996
rect 4963 11936 5027 11940
rect 1423 11452 1487 11456
rect 1423 11396 1427 11452
rect 1427 11396 1483 11452
rect 1483 11396 1487 11452
rect 1423 11392 1487 11396
rect 1503 11452 1567 11456
rect 1503 11396 1507 11452
rect 1507 11396 1563 11452
rect 1563 11396 1567 11452
rect 1503 11392 1567 11396
rect 1583 11452 1647 11456
rect 1583 11396 1587 11452
rect 1587 11396 1643 11452
rect 1643 11396 1647 11452
rect 1583 11392 1647 11396
rect 1663 11452 1727 11456
rect 1663 11396 1667 11452
rect 1667 11396 1723 11452
rect 1723 11396 1727 11452
rect 1663 11392 1727 11396
rect 2366 11452 2430 11456
rect 2366 11396 2370 11452
rect 2370 11396 2426 11452
rect 2426 11396 2430 11452
rect 2366 11392 2430 11396
rect 2446 11452 2510 11456
rect 2446 11396 2450 11452
rect 2450 11396 2506 11452
rect 2506 11396 2510 11452
rect 2446 11392 2510 11396
rect 2526 11452 2590 11456
rect 2526 11396 2530 11452
rect 2530 11396 2586 11452
rect 2586 11396 2590 11452
rect 2526 11392 2590 11396
rect 2606 11452 2670 11456
rect 2606 11396 2610 11452
rect 2610 11396 2666 11452
rect 2666 11396 2670 11452
rect 2606 11392 2670 11396
rect 3309 11452 3373 11456
rect 3309 11396 3313 11452
rect 3313 11396 3369 11452
rect 3369 11396 3373 11452
rect 3309 11392 3373 11396
rect 3389 11452 3453 11456
rect 3389 11396 3393 11452
rect 3393 11396 3449 11452
rect 3449 11396 3453 11452
rect 3389 11392 3453 11396
rect 3469 11452 3533 11456
rect 3469 11396 3473 11452
rect 3473 11396 3529 11452
rect 3529 11396 3533 11452
rect 3469 11392 3533 11396
rect 3549 11452 3613 11456
rect 3549 11396 3553 11452
rect 3553 11396 3609 11452
rect 3609 11396 3613 11452
rect 3549 11392 3613 11396
rect 4252 11452 4316 11456
rect 4252 11396 4256 11452
rect 4256 11396 4312 11452
rect 4312 11396 4316 11452
rect 4252 11392 4316 11396
rect 4332 11452 4396 11456
rect 4332 11396 4336 11452
rect 4336 11396 4392 11452
rect 4392 11396 4396 11452
rect 4332 11392 4396 11396
rect 4412 11452 4476 11456
rect 4412 11396 4416 11452
rect 4416 11396 4472 11452
rect 4472 11396 4476 11452
rect 4412 11392 4476 11396
rect 4492 11452 4556 11456
rect 4492 11396 4496 11452
rect 4496 11396 4552 11452
rect 4552 11396 4556 11452
rect 4492 11392 4556 11396
rect 1894 10908 1958 10912
rect 1894 10852 1898 10908
rect 1898 10852 1954 10908
rect 1954 10852 1958 10908
rect 1894 10848 1958 10852
rect 1974 10908 2038 10912
rect 1974 10852 1978 10908
rect 1978 10852 2034 10908
rect 2034 10852 2038 10908
rect 1974 10848 2038 10852
rect 2054 10908 2118 10912
rect 2054 10852 2058 10908
rect 2058 10852 2114 10908
rect 2114 10852 2118 10908
rect 2054 10848 2118 10852
rect 2134 10908 2198 10912
rect 2134 10852 2138 10908
rect 2138 10852 2194 10908
rect 2194 10852 2198 10908
rect 2134 10848 2198 10852
rect 2837 10908 2901 10912
rect 2837 10852 2841 10908
rect 2841 10852 2897 10908
rect 2897 10852 2901 10908
rect 2837 10848 2901 10852
rect 2917 10908 2981 10912
rect 2917 10852 2921 10908
rect 2921 10852 2977 10908
rect 2977 10852 2981 10908
rect 2917 10848 2981 10852
rect 2997 10908 3061 10912
rect 2997 10852 3001 10908
rect 3001 10852 3057 10908
rect 3057 10852 3061 10908
rect 2997 10848 3061 10852
rect 3077 10908 3141 10912
rect 3077 10852 3081 10908
rect 3081 10852 3137 10908
rect 3137 10852 3141 10908
rect 3077 10848 3141 10852
rect 3780 10908 3844 10912
rect 3780 10852 3784 10908
rect 3784 10852 3840 10908
rect 3840 10852 3844 10908
rect 3780 10848 3844 10852
rect 3860 10908 3924 10912
rect 3860 10852 3864 10908
rect 3864 10852 3920 10908
rect 3920 10852 3924 10908
rect 3860 10848 3924 10852
rect 3940 10908 4004 10912
rect 3940 10852 3944 10908
rect 3944 10852 4000 10908
rect 4000 10852 4004 10908
rect 3940 10848 4004 10852
rect 4020 10908 4084 10912
rect 4020 10852 4024 10908
rect 4024 10852 4080 10908
rect 4080 10852 4084 10908
rect 4020 10848 4084 10852
rect 4723 10908 4787 10912
rect 4723 10852 4727 10908
rect 4727 10852 4783 10908
rect 4783 10852 4787 10908
rect 4723 10848 4787 10852
rect 4803 10908 4867 10912
rect 4803 10852 4807 10908
rect 4807 10852 4863 10908
rect 4863 10852 4867 10908
rect 4803 10848 4867 10852
rect 4883 10908 4947 10912
rect 4883 10852 4887 10908
rect 4887 10852 4943 10908
rect 4943 10852 4947 10908
rect 4883 10848 4947 10852
rect 4963 10908 5027 10912
rect 4963 10852 4967 10908
rect 4967 10852 5023 10908
rect 5023 10852 5027 10908
rect 4963 10848 5027 10852
rect 1423 10364 1487 10368
rect 1423 10308 1427 10364
rect 1427 10308 1483 10364
rect 1483 10308 1487 10364
rect 1423 10304 1487 10308
rect 1503 10364 1567 10368
rect 1503 10308 1507 10364
rect 1507 10308 1563 10364
rect 1563 10308 1567 10364
rect 1503 10304 1567 10308
rect 1583 10364 1647 10368
rect 1583 10308 1587 10364
rect 1587 10308 1643 10364
rect 1643 10308 1647 10364
rect 1583 10304 1647 10308
rect 1663 10364 1727 10368
rect 1663 10308 1667 10364
rect 1667 10308 1723 10364
rect 1723 10308 1727 10364
rect 1663 10304 1727 10308
rect 2366 10364 2430 10368
rect 2366 10308 2370 10364
rect 2370 10308 2426 10364
rect 2426 10308 2430 10364
rect 2366 10304 2430 10308
rect 2446 10364 2510 10368
rect 2446 10308 2450 10364
rect 2450 10308 2506 10364
rect 2506 10308 2510 10364
rect 2446 10304 2510 10308
rect 2526 10364 2590 10368
rect 2526 10308 2530 10364
rect 2530 10308 2586 10364
rect 2586 10308 2590 10364
rect 2526 10304 2590 10308
rect 2606 10364 2670 10368
rect 2606 10308 2610 10364
rect 2610 10308 2666 10364
rect 2666 10308 2670 10364
rect 2606 10304 2670 10308
rect 3309 10364 3373 10368
rect 3309 10308 3313 10364
rect 3313 10308 3369 10364
rect 3369 10308 3373 10364
rect 3309 10304 3373 10308
rect 3389 10364 3453 10368
rect 3389 10308 3393 10364
rect 3393 10308 3449 10364
rect 3449 10308 3453 10364
rect 3389 10304 3453 10308
rect 3469 10364 3533 10368
rect 3469 10308 3473 10364
rect 3473 10308 3529 10364
rect 3529 10308 3533 10364
rect 3469 10304 3533 10308
rect 3549 10364 3613 10368
rect 3549 10308 3553 10364
rect 3553 10308 3609 10364
rect 3609 10308 3613 10364
rect 3549 10304 3613 10308
rect 4252 10364 4316 10368
rect 4252 10308 4256 10364
rect 4256 10308 4312 10364
rect 4312 10308 4316 10364
rect 4252 10304 4316 10308
rect 4332 10364 4396 10368
rect 4332 10308 4336 10364
rect 4336 10308 4392 10364
rect 4392 10308 4396 10364
rect 4332 10304 4396 10308
rect 4412 10364 4476 10368
rect 4412 10308 4416 10364
rect 4416 10308 4472 10364
rect 4472 10308 4476 10364
rect 4412 10304 4476 10308
rect 4492 10364 4556 10368
rect 4492 10308 4496 10364
rect 4496 10308 4552 10364
rect 4552 10308 4556 10364
rect 4492 10304 4556 10308
rect 1894 9820 1958 9824
rect 1894 9764 1898 9820
rect 1898 9764 1954 9820
rect 1954 9764 1958 9820
rect 1894 9760 1958 9764
rect 1974 9820 2038 9824
rect 1974 9764 1978 9820
rect 1978 9764 2034 9820
rect 2034 9764 2038 9820
rect 1974 9760 2038 9764
rect 2054 9820 2118 9824
rect 2054 9764 2058 9820
rect 2058 9764 2114 9820
rect 2114 9764 2118 9820
rect 2054 9760 2118 9764
rect 2134 9820 2198 9824
rect 2134 9764 2138 9820
rect 2138 9764 2194 9820
rect 2194 9764 2198 9820
rect 2134 9760 2198 9764
rect 2837 9820 2901 9824
rect 2837 9764 2841 9820
rect 2841 9764 2897 9820
rect 2897 9764 2901 9820
rect 2837 9760 2901 9764
rect 2917 9820 2981 9824
rect 2917 9764 2921 9820
rect 2921 9764 2977 9820
rect 2977 9764 2981 9820
rect 2917 9760 2981 9764
rect 2997 9820 3061 9824
rect 2997 9764 3001 9820
rect 3001 9764 3057 9820
rect 3057 9764 3061 9820
rect 2997 9760 3061 9764
rect 3077 9820 3141 9824
rect 3077 9764 3081 9820
rect 3081 9764 3137 9820
rect 3137 9764 3141 9820
rect 3077 9760 3141 9764
rect 3780 9820 3844 9824
rect 3780 9764 3784 9820
rect 3784 9764 3840 9820
rect 3840 9764 3844 9820
rect 3780 9760 3844 9764
rect 3860 9820 3924 9824
rect 3860 9764 3864 9820
rect 3864 9764 3920 9820
rect 3920 9764 3924 9820
rect 3860 9760 3924 9764
rect 3940 9820 4004 9824
rect 3940 9764 3944 9820
rect 3944 9764 4000 9820
rect 4000 9764 4004 9820
rect 3940 9760 4004 9764
rect 4020 9820 4084 9824
rect 4020 9764 4024 9820
rect 4024 9764 4080 9820
rect 4080 9764 4084 9820
rect 4020 9760 4084 9764
rect 4723 9820 4787 9824
rect 4723 9764 4727 9820
rect 4727 9764 4783 9820
rect 4783 9764 4787 9820
rect 4723 9760 4787 9764
rect 4803 9820 4867 9824
rect 4803 9764 4807 9820
rect 4807 9764 4863 9820
rect 4863 9764 4867 9820
rect 4803 9760 4867 9764
rect 4883 9820 4947 9824
rect 4883 9764 4887 9820
rect 4887 9764 4943 9820
rect 4943 9764 4947 9820
rect 4883 9760 4947 9764
rect 4963 9820 5027 9824
rect 4963 9764 4967 9820
rect 4967 9764 5023 9820
rect 5023 9764 5027 9820
rect 4963 9760 5027 9764
rect 1423 9276 1487 9280
rect 1423 9220 1427 9276
rect 1427 9220 1483 9276
rect 1483 9220 1487 9276
rect 1423 9216 1487 9220
rect 1503 9276 1567 9280
rect 1503 9220 1507 9276
rect 1507 9220 1563 9276
rect 1563 9220 1567 9276
rect 1503 9216 1567 9220
rect 1583 9276 1647 9280
rect 1583 9220 1587 9276
rect 1587 9220 1643 9276
rect 1643 9220 1647 9276
rect 1583 9216 1647 9220
rect 1663 9276 1727 9280
rect 1663 9220 1667 9276
rect 1667 9220 1723 9276
rect 1723 9220 1727 9276
rect 1663 9216 1727 9220
rect 2366 9276 2430 9280
rect 2366 9220 2370 9276
rect 2370 9220 2426 9276
rect 2426 9220 2430 9276
rect 2366 9216 2430 9220
rect 2446 9276 2510 9280
rect 2446 9220 2450 9276
rect 2450 9220 2506 9276
rect 2506 9220 2510 9276
rect 2446 9216 2510 9220
rect 2526 9276 2590 9280
rect 2526 9220 2530 9276
rect 2530 9220 2586 9276
rect 2586 9220 2590 9276
rect 2526 9216 2590 9220
rect 2606 9276 2670 9280
rect 2606 9220 2610 9276
rect 2610 9220 2666 9276
rect 2666 9220 2670 9276
rect 2606 9216 2670 9220
rect 3309 9276 3373 9280
rect 3309 9220 3313 9276
rect 3313 9220 3369 9276
rect 3369 9220 3373 9276
rect 3309 9216 3373 9220
rect 3389 9276 3453 9280
rect 3389 9220 3393 9276
rect 3393 9220 3449 9276
rect 3449 9220 3453 9276
rect 3389 9216 3453 9220
rect 3469 9276 3533 9280
rect 3469 9220 3473 9276
rect 3473 9220 3529 9276
rect 3529 9220 3533 9276
rect 3469 9216 3533 9220
rect 3549 9276 3613 9280
rect 3549 9220 3553 9276
rect 3553 9220 3609 9276
rect 3609 9220 3613 9276
rect 3549 9216 3613 9220
rect 4252 9276 4316 9280
rect 4252 9220 4256 9276
rect 4256 9220 4312 9276
rect 4312 9220 4316 9276
rect 4252 9216 4316 9220
rect 4332 9276 4396 9280
rect 4332 9220 4336 9276
rect 4336 9220 4392 9276
rect 4392 9220 4396 9276
rect 4332 9216 4396 9220
rect 4412 9276 4476 9280
rect 4412 9220 4416 9276
rect 4416 9220 4472 9276
rect 4472 9220 4476 9276
rect 4412 9216 4476 9220
rect 4492 9276 4556 9280
rect 4492 9220 4496 9276
rect 4496 9220 4552 9276
rect 4552 9220 4556 9276
rect 4492 9216 4556 9220
rect 1894 8732 1958 8736
rect 1894 8676 1898 8732
rect 1898 8676 1954 8732
rect 1954 8676 1958 8732
rect 1894 8672 1958 8676
rect 1974 8732 2038 8736
rect 1974 8676 1978 8732
rect 1978 8676 2034 8732
rect 2034 8676 2038 8732
rect 1974 8672 2038 8676
rect 2054 8732 2118 8736
rect 2054 8676 2058 8732
rect 2058 8676 2114 8732
rect 2114 8676 2118 8732
rect 2054 8672 2118 8676
rect 2134 8732 2198 8736
rect 2134 8676 2138 8732
rect 2138 8676 2194 8732
rect 2194 8676 2198 8732
rect 2134 8672 2198 8676
rect 2837 8732 2901 8736
rect 2837 8676 2841 8732
rect 2841 8676 2897 8732
rect 2897 8676 2901 8732
rect 2837 8672 2901 8676
rect 2917 8732 2981 8736
rect 2917 8676 2921 8732
rect 2921 8676 2977 8732
rect 2977 8676 2981 8732
rect 2917 8672 2981 8676
rect 2997 8732 3061 8736
rect 2997 8676 3001 8732
rect 3001 8676 3057 8732
rect 3057 8676 3061 8732
rect 2997 8672 3061 8676
rect 3077 8732 3141 8736
rect 3077 8676 3081 8732
rect 3081 8676 3137 8732
rect 3137 8676 3141 8732
rect 3077 8672 3141 8676
rect 3780 8732 3844 8736
rect 3780 8676 3784 8732
rect 3784 8676 3840 8732
rect 3840 8676 3844 8732
rect 3780 8672 3844 8676
rect 3860 8732 3924 8736
rect 3860 8676 3864 8732
rect 3864 8676 3920 8732
rect 3920 8676 3924 8732
rect 3860 8672 3924 8676
rect 3940 8732 4004 8736
rect 3940 8676 3944 8732
rect 3944 8676 4000 8732
rect 4000 8676 4004 8732
rect 3940 8672 4004 8676
rect 4020 8732 4084 8736
rect 4020 8676 4024 8732
rect 4024 8676 4080 8732
rect 4080 8676 4084 8732
rect 4020 8672 4084 8676
rect 4723 8732 4787 8736
rect 4723 8676 4727 8732
rect 4727 8676 4783 8732
rect 4783 8676 4787 8732
rect 4723 8672 4787 8676
rect 4803 8732 4867 8736
rect 4803 8676 4807 8732
rect 4807 8676 4863 8732
rect 4863 8676 4867 8732
rect 4803 8672 4867 8676
rect 4883 8732 4947 8736
rect 4883 8676 4887 8732
rect 4887 8676 4943 8732
rect 4943 8676 4947 8732
rect 4883 8672 4947 8676
rect 4963 8732 5027 8736
rect 4963 8676 4967 8732
rect 4967 8676 5023 8732
rect 5023 8676 5027 8732
rect 4963 8672 5027 8676
rect 1423 8188 1487 8192
rect 1423 8132 1427 8188
rect 1427 8132 1483 8188
rect 1483 8132 1487 8188
rect 1423 8128 1487 8132
rect 1503 8188 1567 8192
rect 1503 8132 1507 8188
rect 1507 8132 1563 8188
rect 1563 8132 1567 8188
rect 1503 8128 1567 8132
rect 1583 8188 1647 8192
rect 1583 8132 1587 8188
rect 1587 8132 1643 8188
rect 1643 8132 1647 8188
rect 1583 8128 1647 8132
rect 1663 8188 1727 8192
rect 1663 8132 1667 8188
rect 1667 8132 1723 8188
rect 1723 8132 1727 8188
rect 1663 8128 1727 8132
rect 2366 8188 2430 8192
rect 2366 8132 2370 8188
rect 2370 8132 2426 8188
rect 2426 8132 2430 8188
rect 2366 8128 2430 8132
rect 2446 8188 2510 8192
rect 2446 8132 2450 8188
rect 2450 8132 2506 8188
rect 2506 8132 2510 8188
rect 2446 8128 2510 8132
rect 2526 8188 2590 8192
rect 2526 8132 2530 8188
rect 2530 8132 2586 8188
rect 2586 8132 2590 8188
rect 2526 8128 2590 8132
rect 2606 8188 2670 8192
rect 2606 8132 2610 8188
rect 2610 8132 2666 8188
rect 2666 8132 2670 8188
rect 2606 8128 2670 8132
rect 3309 8188 3373 8192
rect 3309 8132 3313 8188
rect 3313 8132 3369 8188
rect 3369 8132 3373 8188
rect 3309 8128 3373 8132
rect 3389 8188 3453 8192
rect 3389 8132 3393 8188
rect 3393 8132 3449 8188
rect 3449 8132 3453 8188
rect 3389 8128 3453 8132
rect 3469 8188 3533 8192
rect 3469 8132 3473 8188
rect 3473 8132 3529 8188
rect 3529 8132 3533 8188
rect 3469 8128 3533 8132
rect 3549 8188 3613 8192
rect 3549 8132 3553 8188
rect 3553 8132 3609 8188
rect 3609 8132 3613 8188
rect 3549 8128 3613 8132
rect 4252 8188 4316 8192
rect 4252 8132 4256 8188
rect 4256 8132 4312 8188
rect 4312 8132 4316 8188
rect 4252 8128 4316 8132
rect 4332 8188 4396 8192
rect 4332 8132 4336 8188
rect 4336 8132 4392 8188
rect 4392 8132 4396 8188
rect 4332 8128 4396 8132
rect 4412 8188 4476 8192
rect 4412 8132 4416 8188
rect 4416 8132 4472 8188
rect 4472 8132 4476 8188
rect 4412 8128 4476 8132
rect 4492 8188 4556 8192
rect 4492 8132 4496 8188
rect 4496 8132 4552 8188
rect 4552 8132 4556 8188
rect 4492 8128 4556 8132
rect 1894 7644 1958 7648
rect 1894 7588 1898 7644
rect 1898 7588 1954 7644
rect 1954 7588 1958 7644
rect 1894 7584 1958 7588
rect 1974 7644 2038 7648
rect 1974 7588 1978 7644
rect 1978 7588 2034 7644
rect 2034 7588 2038 7644
rect 1974 7584 2038 7588
rect 2054 7644 2118 7648
rect 2054 7588 2058 7644
rect 2058 7588 2114 7644
rect 2114 7588 2118 7644
rect 2054 7584 2118 7588
rect 2134 7644 2198 7648
rect 2134 7588 2138 7644
rect 2138 7588 2194 7644
rect 2194 7588 2198 7644
rect 2134 7584 2198 7588
rect 2837 7644 2901 7648
rect 2837 7588 2841 7644
rect 2841 7588 2897 7644
rect 2897 7588 2901 7644
rect 2837 7584 2901 7588
rect 2917 7644 2981 7648
rect 2917 7588 2921 7644
rect 2921 7588 2977 7644
rect 2977 7588 2981 7644
rect 2917 7584 2981 7588
rect 2997 7644 3061 7648
rect 2997 7588 3001 7644
rect 3001 7588 3057 7644
rect 3057 7588 3061 7644
rect 2997 7584 3061 7588
rect 3077 7644 3141 7648
rect 3077 7588 3081 7644
rect 3081 7588 3137 7644
rect 3137 7588 3141 7644
rect 3077 7584 3141 7588
rect 3780 7644 3844 7648
rect 3780 7588 3784 7644
rect 3784 7588 3840 7644
rect 3840 7588 3844 7644
rect 3780 7584 3844 7588
rect 3860 7644 3924 7648
rect 3860 7588 3864 7644
rect 3864 7588 3920 7644
rect 3920 7588 3924 7644
rect 3860 7584 3924 7588
rect 3940 7644 4004 7648
rect 3940 7588 3944 7644
rect 3944 7588 4000 7644
rect 4000 7588 4004 7644
rect 3940 7584 4004 7588
rect 4020 7644 4084 7648
rect 4020 7588 4024 7644
rect 4024 7588 4080 7644
rect 4080 7588 4084 7644
rect 4020 7584 4084 7588
rect 4723 7644 4787 7648
rect 4723 7588 4727 7644
rect 4727 7588 4783 7644
rect 4783 7588 4787 7644
rect 4723 7584 4787 7588
rect 4803 7644 4867 7648
rect 4803 7588 4807 7644
rect 4807 7588 4863 7644
rect 4863 7588 4867 7644
rect 4803 7584 4867 7588
rect 4883 7644 4947 7648
rect 4883 7588 4887 7644
rect 4887 7588 4943 7644
rect 4943 7588 4947 7644
rect 4883 7584 4947 7588
rect 4963 7644 5027 7648
rect 4963 7588 4967 7644
rect 4967 7588 5023 7644
rect 5023 7588 5027 7644
rect 4963 7584 5027 7588
rect 1423 7100 1487 7104
rect 1423 7044 1427 7100
rect 1427 7044 1483 7100
rect 1483 7044 1487 7100
rect 1423 7040 1487 7044
rect 1503 7100 1567 7104
rect 1503 7044 1507 7100
rect 1507 7044 1563 7100
rect 1563 7044 1567 7100
rect 1503 7040 1567 7044
rect 1583 7100 1647 7104
rect 1583 7044 1587 7100
rect 1587 7044 1643 7100
rect 1643 7044 1647 7100
rect 1583 7040 1647 7044
rect 1663 7100 1727 7104
rect 1663 7044 1667 7100
rect 1667 7044 1723 7100
rect 1723 7044 1727 7100
rect 1663 7040 1727 7044
rect 2366 7100 2430 7104
rect 2366 7044 2370 7100
rect 2370 7044 2426 7100
rect 2426 7044 2430 7100
rect 2366 7040 2430 7044
rect 2446 7100 2510 7104
rect 2446 7044 2450 7100
rect 2450 7044 2506 7100
rect 2506 7044 2510 7100
rect 2446 7040 2510 7044
rect 2526 7100 2590 7104
rect 2526 7044 2530 7100
rect 2530 7044 2586 7100
rect 2586 7044 2590 7100
rect 2526 7040 2590 7044
rect 2606 7100 2670 7104
rect 2606 7044 2610 7100
rect 2610 7044 2666 7100
rect 2666 7044 2670 7100
rect 2606 7040 2670 7044
rect 3309 7100 3373 7104
rect 3309 7044 3313 7100
rect 3313 7044 3369 7100
rect 3369 7044 3373 7100
rect 3309 7040 3373 7044
rect 3389 7100 3453 7104
rect 3389 7044 3393 7100
rect 3393 7044 3449 7100
rect 3449 7044 3453 7100
rect 3389 7040 3453 7044
rect 3469 7100 3533 7104
rect 3469 7044 3473 7100
rect 3473 7044 3529 7100
rect 3529 7044 3533 7100
rect 3469 7040 3533 7044
rect 3549 7100 3613 7104
rect 3549 7044 3553 7100
rect 3553 7044 3609 7100
rect 3609 7044 3613 7100
rect 3549 7040 3613 7044
rect 4252 7100 4316 7104
rect 4252 7044 4256 7100
rect 4256 7044 4312 7100
rect 4312 7044 4316 7100
rect 4252 7040 4316 7044
rect 4332 7100 4396 7104
rect 4332 7044 4336 7100
rect 4336 7044 4392 7100
rect 4392 7044 4396 7100
rect 4332 7040 4396 7044
rect 4412 7100 4476 7104
rect 4412 7044 4416 7100
rect 4416 7044 4472 7100
rect 4472 7044 4476 7100
rect 4412 7040 4476 7044
rect 4492 7100 4556 7104
rect 4492 7044 4496 7100
rect 4496 7044 4552 7100
rect 4552 7044 4556 7100
rect 4492 7040 4556 7044
rect 1894 6556 1958 6560
rect 1894 6500 1898 6556
rect 1898 6500 1954 6556
rect 1954 6500 1958 6556
rect 1894 6496 1958 6500
rect 1974 6556 2038 6560
rect 1974 6500 1978 6556
rect 1978 6500 2034 6556
rect 2034 6500 2038 6556
rect 1974 6496 2038 6500
rect 2054 6556 2118 6560
rect 2054 6500 2058 6556
rect 2058 6500 2114 6556
rect 2114 6500 2118 6556
rect 2054 6496 2118 6500
rect 2134 6556 2198 6560
rect 2134 6500 2138 6556
rect 2138 6500 2194 6556
rect 2194 6500 2198 6556
rect 2134 6496 2198 6500
rect 2837 6556 2901 6560
rect 2837 6500 2841 6556
rect 2841 6500 2897 6556
rect 2897 6500 2901 6556
rect 2837 6496 2901 6500
rect 2917 6556 2981 6560
rect 2917 6500 2921 6556
rect 2921 6500 2977 6556
rect 2977 6500 2981 6556
rect 2917 6496 2981 6500
rect 2997 6556 3061 6560
rect 2997 6500 3001 6556
rect 3001 6500 3057 6556
rect 3057 6500 3061 6556
rect 2997 6496 3061 6500
rect 3077 6556 3141 6560
rect 3077 6500 3081 6556
rect 3081 6500 3137 6556
rect 3137 6500 3141 6556
rect 3077 6496 3141 6500
rect 3780 6556 3844 6560
rect 3780 6500 3784 6556
rect 3784 6500 3840 6556
rect 3840 6500 3844 6556
rect 3780 6496 3844 6500
rect 3860 6556 3924 6560
rect 3860 6500 3864 6556
rect 3864 6500 3920 6556
rect 3920 6500 3924 6556
rect 3860 6496 3924 6500
rect 3940 6556 4004 6560
rect 3940 6500 3944 6556
rect 3944 6500 4000 6556
rect 4000 6500 4004 6556
rect 3940 6496 4004 6500
rect 4020 6556 4084 6560
rect 4020 6500 4024 6556
rect 4024 6500 4080 6556
rect 4080 6500 4084 6556
rect 4020 6496 4084 6500
rect 4723 6556 4787 6560
rect 4723 6500 4727 6556
rect 4727 6500 4783 6556
rect 4783 6500 4787 6556
rect 4723 6496 4787 6500
rect 4803 6556 4867 6560
rect 4803 6500 4807 6556
rect 4807 6500 4863 6556
rect 4863 6500 4867 6556
rect 4803 6496 4867 6500
rect 4883 6556 4947 6560
rect 4883 6500 4887 6556
rect 4887 6500 4943 6556
rect 4943 6500 4947 6556
rect 4883 6496 4947 6500
rect 4963 6556 5027 6560
rect 4963 6500 4967 6556
rect 4967 6500 5023 6556
rect 5023 6500 5027 6556
rect 4963 6496 5027 6500
rect 1423 6012 1487 6016
rect 1423 5956 1427 6012
rect 1427 5956 1483 6012
rect 1483 5956 1487 6012
rect 1423 5952 1487 5956
rect 1503 6012 1567 6016
rect 1503 5956 1507 6012
rect 1507 5956 1563 6012
rect 1563 5956 1567 6012
rect 1503 5952 1567 5956
rect 1583 6012 1647 6016
rect 1583 5956 1587 6012
rect 1587 5956 1643 6012
rect 1643 5956 1647 6012
rect 1583 5952 1647 5956
rect 1663 6012 1727 6016
rect 1663 5956 1667 6012
rect 1667 5956 1723 6012
rect 1723 5956 1727 6012
rect 1663 5952 1727 5956
rect 2366 6012 2430 6016
rect 2366 5956 2370 6012
rect 2370 5956 2426 6012
rect 2426 5956 2430 6012
rect 2366 5952 2430 5956
rect 2446 6012 2510 6016
rect 2446 5956 2450 6012
rect 2450 5956 2506 6012
rect 2506 5956 2510 6012
rect 2446 5952 2510 5956
rect 2526 6012 2590 6016
rect 2526 5956 2530 6012
rect 2530 5956 2586 6012
rect 2586 5956 2590 6012
rect 2526 5952 2590 5956
rect 2606 6012 2670 6016
rect 2606 5956 2610 6012
rect 2610 5956 2666 6012
rect 2666 5956 2670 6012
rect 2606 5952 2670 5956
rect 3309 6012 3373 6016
rect 3309 5956 3313 6012
rect 3313 5956 3369 6012
rect 3369 5956 3373 6012
rect 3309 5952 3373 5956
rect 3389 6012 3453 6016
rect 3389 5956 3393 6012
rect 3393 5956 3449 6012
rect 3449 5956 3453 6012
rect 3389 5952 3453 5956
rect 3469 6012 3533 6016
rect 3469 5956 3473 6012
rect 3473 5956 3529 6012
rect 3529 5956 3533 6012
rect 3469 5952 3533 5956
rect 3549 6012 3613 6016
rect 3549 5956 3553 6012
rect 3553 5956 3609 6012
rect 3609 5956 3613 6012
rect 3549 5952 3613 5956
rect 4252 6012 4316 6016
rect 4252 5956 4256 6012
rect 4256 5956 4312 6012
rect 4312 5956 4316 6012
rect 4252 5952 4316 5956
rect 4332 6012 4396 6016
rect 4332 5956 4336 6012
rect 4336 5956 4392 6012
rect 4392 5956 4396 6012
rect 4332 5952 4396 5956
rect 4412 6012 4476 6016
rect 4412 5956 4416 6012
rect 4416 5956 4472 6012
rect 4472 5956 4476 6012
rect 4412 5952 4476 5956
rect 4492 6012 4556 6016
rect 4492 5956 4496 6012
rect 4496 5956 4552 6012
rect 4552 5956 4556 6012
rect 4492 5952 4556 5956
rect 1894 5468 1958 5472
rect 1894 5412 1898 5468
rect 1898 5412 1954 5468
rect 1954 5412 1958 5468
rect 1894 5408 1958 5412
rect 1974 5468 2038 5472
rect 1974 5412 1978 5468
rect 1978 5412 2034 5468
rect 2034 5412 2038 5468
rect 1974 5408 2038 5412
rect 2054 5468 2118 5472
rect 2054 5412 2058 5468
rect 2058 5412 2114 5468
rect 2114 5412 2118 5468
rect 2054 5408 2118 5412
rect 2134 5468 2198 5472
rect 2134 5412 2138 5468
rect 2138 5412 2194 5468
rect 2194 5412 2198 5468
rect 2134 5408 2198 5412
rect 2837 5468 2901 5472
rect 2837 5412 2841 5468
rect 2841 5412 2897 5468
rect 2897 5412 2901 5468
rect 2837 5408 2901 5412
rect 2917 5468 2981 5472
rect 2917 5412 2921 5468
rect 2921 5412 2977 5468
rect 2977 5412 2981 5468
rect 2917 5408 2981 5412
rect 2997 5468 3061 5472
rect 2997 5412 3001 5468
rect 3001 5412 3057 5468
rect 3057 5412 3061 5468
rect 2997 5408 3061 5412
rect 3077 5468 3141 5472
rect 3077 5412 3081 5468
rect 3081 5412 3137 5468
rect 3137 5412 3141 5468
rect 3077 5408 3141 5412
rect 3780 5468 3844 5472
rect 3780 5412 3784 5468
rect 3784 5412 3840 5468
rect 3840 5412 3844 5468
rect 3780 5408 3844 5412
rect 3860 5468 3924 5472
rect 3860 5412 3864 5468
rect 3864 5412 3920 5468
rect 3920 5412 3924 5468
rect 3860 5408 3924 5412
rect 3940 5468 4004 5472
rect 3940 5412 3944 5468
rect 3944 5412 4000 5468
rect 4000 5412 4004 5468
rect 3940 5408 4004 5412
rect 4020 5468 4084 5472
rect 4020 5412 4024 5468
rect 4024 5412 4080 5468
rect 4080 5412 4084 5468
rect 4020 5408 4084 5412
rect 4723 5468 4787 5472
rect 4723 5412 4727 5468
rect 4727 5412 4783 5468
rect 4783 5412 4787 5468
rect 4723 5408 4787 5412
rect 4803 5468 4867 5472
rect 4803 5412 4807 5468
rect 4807 5412 4863 5468
rect 4863 5412 4867 5468
rect 4803 5408 4867 5412
rect 4883 5468 4947 5472
rect 4883 5412 4887 5468
rect 4887 5412 4943 5468
rect 4943 5412 4947 5468
rect 4883 5408 4947 5412
rect 4963 5468 5027 5472
rect 4963 5412 4967 5468
rect 4967 5412 5023 5468
rect 5023 5412 5027 5468
rect 4963 5408 5027 5412
rect 1423 4924 1487 4928
rect 1423 4868 1427 4924
rect 1427 4868 1483 4924
rect 1483 4868 1487 4924
rect 1423 4864 1487 4868
rect 1503 4924 1567 4928
rect 1503 4868 1507 4924
rect 1507 4868 1563 4924
rect 1563 4868 1567 4924
rect 1503 4864 1567 4868
rect 1583 4924 1647 4928
rect 1583 4868 1587 4924
rect 1587 4868 1643 4924
rect 1643 4868 1647 4924
rect 1583 4864 1647 4868
rect 1663 4924 1727 4928
rect 1663 4868 1667 4924
rect 1667 4868 1723 4924
rect 1723 4868 1727 4924
rect 1663 4864 1727 4868
rect 2366 4924 2430 4928
rect 2366 4868 2370 4924
rect 2370 4868 2426 4924
rect 2426 4868 2430 4924
rect 2366 4864 2430 4868
rect 2446 4924 2510 4928
rect 2446 4868 2450 4924
rect 2450 4868 2506 4924
rect 2506 4868 2510 4924
rect 2446 4864 2510 4868
rect 2526 4924 2590 4928
rect 2526 4868 2530 4924
rect 2530 4868 2586 4924
rect 2586 4868 2590 4924
rect 2526 4864 2590 4868
rect 2606 4924 2670 4928
rect 2606 4868 2610 4924
rect 2610 4868 2666 4924
rect 2666 4868 2670 4924
rect 2606 4864 2670 4868
rect 3309 4924 3373 4928
rect 3309 4868 3313 4924
rect 3313 4868 3369 4924
rect 3369 4868 3373 4924
rect 3309 4864 3373 4868
rect 3389 4924 3453 4928
rect 3389 4868 3393 4924
rect 3393 4868 3449 4924
rect 3449 4868 3453 4924
rect 3389 4864 3453 4868
rect 3469 4924 3533 4928
rect 3469 4868 3473 4924
rect 3473 4868 3529 4924
rect 3529 4868 3533 4924
rect 3469 4864 3533 4868
rect 3549 4924 3613 4928
rect 3549 4868 3553 4924
rect 3553 4868 3609 4924
rect 3609 4868 3613 4924
rect 3549 4864 3613 4868
rect 4252 4924 4316 4928
rect 4252 4868 4256 4924
rect 4256 4868 4312 4924
rect 4312 4868 4316 4924
rect 4252 4864 4316 4868
rect 4332 4924 4396 4928
rect 4332 4868 4336 4924
rect 4336 4868 4392 4924
rect 4392 4868 4396 4924
rect 4332 4864 4396 4868
rect 4412 4924 4476 4928
rect 4412 4868 4416 4924
rect 4416 4868 4472 4924
rect 4472 4868 4476 4924
rect 4412 4864 4476 4868
rect 4492 4924 4556 4928
rect 4492 4868 4496 4924
rect 4496 4868 4552 4924
rect 4552 4868 4556 4924
rect 4492 4864 4556 4868
rect 1894 4380 1958 4384
rect 1894 4324 1898 4380
rect 1898 4324 1954 4380
rect 1954 4324 1958 4380
rect 1894 4320 1958 4324
rect 1974 4380 2038 4384
rect 1974 4324 1978 4380
rect 1978 4324 2034 4380
rect 2034 4324 2038 4380
rect 1974 4320 2038 4324
rect 2054 4380 2118 4384
rect 2054 4324 2058 4380
rect 2058 4324 2114 4380
rect 2114 4324 2118 4380
rect 2054 4320 2118 4324
rect 2134 4380 2198 4384
rect 2134 4324 2138 4380
rect 2138 4324 2194 4380
rect 2194 4324 2198 4380
rect 2134 4320 2198 4324
rect 2837 4380 2901 4384
rect 2837 4324 2841 4380
rect 2841 4324 2897 4380
rect 2897 4324 2901 4380
rect 2837 4320 2901 4324
rect 2917 4380 2981 4384
rect 2917 4324 2921 4380
rect 2921 4324 2977 4380
rect 2977 4324 2981 4380
rect 2917 4320 2981 4324
rect 2997 4380 3061 4384
rect 2997 4324 3001 4380
rect 3001 4324 3057 4380
rect 3057 4324 3061 4380
rect 2997 4320 3061 4324
rect 3077 4380 3141 4384
rect 3077 4324 3081 4380
rect 3081 4324 3137 4380
rect 3137 4324 3141 4380
rect 3077 4320 3141 4324
rect 3780 4380 3844 4384
rect 3780 4324 3784 4380
rect 3784 4324 3840 4380
rect 3840 4324 3844 4380
rect 3780 4320 3844 4324
rect 3860 4380 3924 4384
rect 3860 4324 3864 4380
rect 3864 4324 3920 4380
rect 3920 4324 3924 4380
rect 3860 4320 3924 4324
rect 3940 4380 4004 4384
rect 3940 4324 3944 4380
rect 3944 4324 4000 4380
rect 4000 4324 4004 4380
rect 3940 4320 4004 4324
rect 4020 4380 4084 4384
rect 4020 4324 4024 4380
rect 4024 4324 4080 4380
rect 4080 4324 4084 4380
rect 4020 4320 4084 4324
rect 4723 4380 4787 4384
rect 4723 4324 4727 4380
rect 4727 4324 4783 4380
rect 4783 4324 4787 4380
rect 4723 4320 4787 4324
rect 4803 4380 4867 4384
rect 4803 4324 4807 4380
rect 4807 4324 4863 4380
rect 4863 4324 4867 4380
rect 4803 4320 4867 4324
rect 4883 4380 4947 4384
rect 4883 4324 4887 4380
rect 4887 4324 4943 4380
rect 4943 4324 4947 4380
rect 4883 4320 4947 4324
rect 4963 4380 5027 4384
rect 4963 4324 4967 4380
rect 4967 4324 5023 4380
rect 5023 4324 5027 4380
rect 4963 4320 5027 4324
rect 1423 3836 1487 3840
rect 1423 3780 1427 3836
rect 1427 3780 1483 3836
rect 1483 3780 1487 3836
rect 1423 3776 1487 3780
rect 1503 3836 1567 3840
rect 1503 3780 1507 3836
rect 1507 3780 1563 3836
rect 1563 3780 1567 3836
rect 1503 3776 1567 3780
rect 1583 3836 1647 3840
rect 1583 3780 1587 3836
rect 1587 3780 1643 3836
rect 1643 3780 1647 3836
rect 1583 3776 1647 3780
rect 1663 3836 1727 3840
rect 1663 3780 1667 3836
rect 1667 3780 1723 3836
rect 1723 3780 1727 3836
rect 1663 3776 1727 3780
rect 2366 3836 2430 3840
rect 2366 3780 2370 3836
rect 2370 3780 2426 3836
rect 2426 3780 2430 3836
rect 2366 3776 2430 3780
rect 2446 3836 2510 3840
rect 2446 3780 2450 3836
rect 2450 3780 2506 3836
rect 2506 3780 2510 3836
rect 2446 3776 2510 3780
rect 2526 3836 2590 3840
rect 2526 3780 2530 3836
rect 2530 3780 2586 3836
rect 2586 3780 2590 3836
rect 2526 3776 2590 3780
rect 2606 3836 2670 3840
rect 2606 3780 2610 3836
rect 2610 3780 2666 3836
rect 2666 3780 2670 3836
rect 2606 3776 2670 3780
rect 3309 3836 3373 3840
rect 3309 3780 3313 3836
rect 3313 3780 3369 3836
rect 3369 3780 3373 3836
rect 3309 3776 3373 3780
rect 3389 3836 3453 3840
rect 3389 3780 3393 3836
rect 3393 3780 3449 3836
rect 3449 3780 3453 3836
rect 3389 3776 3453 3780
rect 3469 3836 3533 3840
rect 3469 3780 3473 3836
rect 3473 3780 3529 3836
rect 3529 3780 3533 3836
rect 3469 3776 3533 3780
rect 3549 3836 3613 3840
rect 3549 3780 3553 3836
rect 3553 3780 3609 3836
rect 3609 3780 3613 3836
rect 3549 3776 3613 3780
rect 4252 3836 4316 3840
rect 4252 3780 4256 3836
rect 4256 3780 4312 3836
rect 4312 3780 4316 3836
rect 4252 3776 4316 3780
rect 4332 3836 4396 3840
rect 4332 3780 4336 3836
rect 4336 3780 4392 3836
rect 4392 3780 4396 3836
rect 4332 3776 4396 3780
rect 4412 3836 4476 3840
rect 4412 3780 4416 3836
rect 4416 3780 4472 3836
rect 4472 3780 4476 3836
rect 4412 3776 4476 3780
rect 4492 3836 4556 3840
rect 4492 3780 4496 3836
rect 4496 3780 4552 3836
rect 4552 3780 4556 3836
rect 4492 3776 4556 3780
rect 1894 3292 1958 3296
rect 1894 3236 1898 3292
rect 1898 3236 1954 3292
rect 1954 3236 1958 3292
rect 1894 3232 1958 3236
rect 1974 3292 2038 3296
rect 1974 3236 1978 3292
rect 1978 3236 2034 3292
rect 2034 3236 2038 3292
rect 1974 3232 2038 3236
rect 2054 3292 2118 3296
rect 2054 3236 2058 3292
rect 2058 3236 2114 3292
rect 2114 3236 2118 3292
rect 2054 3232 2118 3236
rect 2134 3292 2198 3296
rect 2134 3236 2138 3292
rect 2138 3236 2194 3292
rect 2194 3236 2198 3292
rect 2134 3232 2198 3236
rect 2837 3292 2901 3296
rect 2837 3236 2841 3292
rect 2841 3236 2897 3292
rect 2897 3236 2901 3292
rect 2837 3232 2901 3236
rect 2917 3292 2981 3296
rect 2917 3236 2921 3292
rect 2921 3236 2977 3292
rect 2977 3236 2981 3292
rect 2917 3232 2981 3236
rect 2997 3292 3061 3296
rect 2997 3236 3001 3292
rect 3001 3236 3057 3292
rect 3057 3236 3061 3292
rect 2997 3232 3061 3236
rect 3077 3292 3141 3296
rect 3077 3236 3081 3292
rect 3081 3236 3137 3292
rect 3137 3236 3141 3292
rect 3077 3232 3141 3236
rect 3780 3292 3844 3296
rect 3780 3236 3784 3292
rect 3784 3236 3840 3292
rect 3840 3236 3844 3292
rect 3780 3232 3844 3236
rect 3860 3292 3924 3296
rect 3860 3236 3864 3292
rect 3864 3236 3920 3292
rect 3920 3236 3924 3292
rect 3860 3232 3924 3236
rect 3940 3292 4004 3296
rect 3940 3236 3944 3292
rect 3944 3236 4000 3292
rect 4000 3236 4004 3292
rect 3940 3232 4004 3236
rect 4020 3292 4084 3296
rect 4020 3236 4024 3292
rect 4024 3236 4080 3292
rect 4080 3236 4084 3292
rect 4020 3232 4084 3236
rect 4723 3292 4787 3296
rect 4723 3236 4727 3292
rect 4727 3236 4783 3292
rect 4783 3236 4787 3292
rect 4723 3232 4787 3236
rect 4803 3292 4867 3296
rect 4803 3236 4807 3292
rect 4807 3236 4863 3292
rect 4863 3236 4867 3292
rect 4803 3232 4867 3236
rect 4883 3292 4947 3296
rect 4883 3236 4887 3292
rect 4887 3236 4943 3292
rect 4943 3236 4947 3292
rect 4883 3232 4947 3236
rect 4963 3292 5027 3296
rect 4963 3236 4967 3292
rect 4967 3236 5023 3292
rect 5023 3236 5027 3292
rect 4963 3232 5027 3236
rect 1423 2748 1487 2752
rect 1423 2692 1427 2748
rect 1427 2692 1483 2748
rect 1483 2692 1487 2748
rect 1423 2688 1487 2692
rect 1503 2748 1567 2752
rect 1503 2692 1507 2748
rect 1507 2692 1563 2748
rect 1563 2692 1567 2748
rect 1503 2688 1567 2692
rect 1583 2748 1647 2752
rect 1583 2692 1587 2748
rect 1587 2692 1643 2748
rect 1643 2692 1647 2748
rect 1583 2688 1647 2692
rect 1663 2748 1727 2752
rect 1663 2692 1667 2748
rect 1667 2692 1723 2748
rect 1723 2692 1727 2748
rect 1663 2688 1727 2692
rect 2366 2748 2430 2752
rect 2366 2692 2370 2748
rect 2370 2692 2426 2748
rect 2426 2692 2430 2748
rect 2366 2688 2430 2692
rect 2446 2748 2510 2752
rect 2446 2692 2450 2748
rect 2450 2692 2506 2748
rect 2506 2692 2510 2748
rect 2446 2688 2510 2692
rect 2526 2748 2590 2752
rect 2526 2692 2530 2748
rect 2530 2692 2586 2748
rect 2586 2692 2590 2748
rect 2526 2688 2590 2692
rect 2606 2748 2670 2752
rect 2606 2692 2610 2748
rect 2610 2692 2666 2748
rect 2666 2692 2670 2748
rect 2606 2688 2670 2692
rect 3309 2748 3373 2752
rect 3309 2692 3313 2748
rect 3313 2692 3369 2748
rect 3369 2692 3373 2748
rect 3309 2688 3373 2692
rect 3389 2748 3453 2752
rect 3389 2692 3393 2748
rect 3393 2692 3449 2748
rect 3449 2692 3453 2748
rect 3389 2688 3453 2692
rect 3469 2748 3533 2752
rect 3469 2692 3473 2748
rect 3473 2692 3529 2748
rect 3529 2692 3533 2748
rect 3469 2688 3533 2692
rect 3549 2748 3613 2752
rect 3549 2692 3553 2748
rect 3553 2692 3609 2748
rect 3609 2692 3613 2748
rect 3549 2688 3613 2692
rect 4252 2748 4316 2752
rect 4252 2692 4256 2748
rect 4256 2692 4312 2748
rect 4312 2692 4316 2748
rect 4252 2688 4316 2692
rect 4332 2748 4396 2752
rect 4332 2692 4336 2748
rect 4336 2692 4392 2748
rect 4392 2692 4396 2748
rect 4332 2688 4396 2692
rect 4412 2748 4476 2752
rect 4412 2692 4416 2748
rect 4416 2692 4472 2748
rect 4472 2692 4476 2748
rect 4412 2688 4476 2692
rect 4492 2748 4556 2752
rect 4492 2692 4496 2748
rect 4496 2692 4552 2748
rect 4552 2692 4556 2748
rect 4492 2688 4556 2692
rect 1894 2204 1958 2208
rect 1894 2148 1898 2204
rect 1898 2148 1954 2204
rect 1954 2148 1958 2204
rect 1894 2144 1958 2148
rect 1974 2204 2038 2208
rect 1974 2148 1978 2204
rect 1978 2148 2034 2204
rect 2034 2148 2038 2204
rect 1974 2144 2038 2148
rect 2054 2204 2118 2208
rect 2054 2148 2058 2204
rect 2058 2148 2114 2204
rect 2114 2148 2118 2204
rect 2054 2144 2118 2148
rect 2134 2204 2198 2208
rect 2134 2148 2138 2204
rect 2138 2148 2194 2204
rect 2194 2148 2198 2204
rect 2134 2144 2198 2148
rect 2837 2204 2901 2208
rect 2837 2148 2841 2204
rect 2841 2148 2897 2204
rect 2897 2148 2901 2204
rect 2837 2144 2901 2148
rect 2917 2204 2981 2208
rect 2917 2148 2921 2204
rect 2921 2148 2977 2204
rect 2977 2148 2981 2204
rect 2917 2144 2981 2148
rect 2997 2204 3061 2208
rect 2997 2148 3001 2204
rect 3001 2148 3057 2204
rect 3057 2148 3061 2204
rect 2997 2144 3061 2148
rect 3077 2204 3141 2208
rect 3077 2148 3081 2204
rect 3081 2148 3137 2204
rect 3137 2148 3141 2204
rect 3077 2144 3141 2148
rect 3780 2204 3844 2208
rect 3780 2148 3784 2204
rect 3784 2148 3840 2204
rect 3840 2148 3844 2204
rect 3780 2144 3844 2148
rect 3860 2204 3924 2208
rect 3860 2148 3864 2204
rect 3864 2148 3920 2204
rect 3920 2148 3924 2204
rect 3860 2144 3924 2148
rect 3940 2204 4004 2208
rect 3940 2148 3944 2204
rect 3944 2148 4000 2204
rect 4000 2148 4004 2204
rect 3940 2144 4004 2148
rect 4020 2204 4084 2208
rect 4020 2148 4024 2204
rect 4024 2148 4080 2204
rect 4080 2148 4084 2204
rect 4020 2144 4084 2148
rect 4723 2204 4787 2208
rect 4723 2148 4727 2204
rect 4727 2148 4783 2204
rect 4783 2148 4787 2204
rect 4723 2144 4787 2148
rect 4803 2204 4867 2208
rect 4803 2148 4807 2204
rect 4807 2148 4863 2204
rect 4863 2148 4867 2204
rect 4803 2144 4867 2148
rect 4883 2204 4947 2208
rect 4883 2148 4887 2204
rect 4887 2148 4943 2204
rect 4943 2148 4947 2204
rect 4883 2144 4947 2148
rect 4963 2204 5027 2208
rect 4963 2148 4967 2204
rect 4967 2148 5023 2204
rect 5023 2148 5027 2204
rect 4963 2144 5027 2148
rect 1423 1660 1487 1664
rect 1423 1604 1427 1660
rect 1427 1604 1483 1660
rect 1483 1604 1487 1660
rect 1423 1600 1487 1604
rect 1503 1660 1567 1664
rect 1503 1604 1507 1660
rect 1507 1604 1563 1660
rect 1563 1604 1567 1660
rect 1503 1600 1567 1604
rect 1583 1660 1647 1664
rect 1583 1604 1587 1660
rect 1587 1604 1643 1660
rect 1643 1604 1647 1660
rect 1583 1600 1647 1604
rect 1663 1660 1727 1664
rect 1663 1604 1667 1660
rect 1667 1604 1723 1660
rect 1723 1604 1727 1660
rect 1663 1600 1727 1604
rect 2366 1660 2430 1664
rect 2366 1604 2370 1660
rect 2370 1604 2426 1660
rect 2426 1604 2430 1660
rect 2366 1600 2430 1604
rect 2446 1660 2510 1664
rect 2446 1604 2450 1660
rect 2450 1604 2506 1660
rect 2506 1604 2510 1660
rect 2446 1600 2510 1604
rect 2526 1660 2590 1664
rect 2526 1604 2530 1660
rect 2530 1604 2586 1660
rect 2586 1604 2590 1660
rect 2526 1600 2590 1604
rect 2606 1660 2670 1664
rect 2606 1604 2610 1660
rect 2610 1604 2666 1660
rect 2666 1604 2670 1660
rect 2606 1600 2670 1604
rect 3309 1660 3373 1664
rect 3309 1604 3313 1660
rect 3313 1604 3369 1660
rect 3369 1604 3373 1660
rect 3309 1600 3373 1604
rect 3389 1660 3453 1664
rect 3389 1604 3393 1660
rect 3393 1604 3449 1660
rect 3449 1604 3453 1660
rect 3389 1600 3453 1604
rect 3469 1660 3533 1664
rect 3469 1604 3473 1660
rect 3473 1604 3529 1660
rect 3529 1604 3533 1660
rect 3469 1600 3533 1604
rect 3549 1660 3613 1664
rect 3549 1604 3553 1660
rect 3553 1604 3609 1660
rect 3609 1604 3613 1660
rect 3549 1600 3613 1604
rect 4252 1660 4316 1664
rect 4252 1604 4256 1660
rect 4256 1604 4312 1660
rect 4312 1604 4316 1660
rect 4252 1600 4316 1604
rect 4332 1660 4396 1664
rect 4332 1604 4336 1660
rect 4336 1604 4392 1660
rect 4392 1604 4396 1660
rect 4332 1600 4396 1604
rect 4412 1660 4476 1664
rect 4412 1604 4416 1660
rect 4416 1604 4472 1660
rect 4472 1604 4476 1660
rect 4412 1600 4476 1604
rect 4492 1660 4556 1664
rect 4492 1604 4496 1660
rect 4496 1604 4552 1660
rect 4552 1604 4556 1660
rect 4492 1600 4556 1604
rect 1894 1116 1958 1120
rect 1894 1060 1898 1116
rect 1898 1060 1954 1116
rect 1954 1060 1958 1116
rect 1894 1056 1958 1060
rect 1974 1116 2038 1120
rect 1974 1060 1978 1116
rect 1978 1060 2034 1116
rect 2034 1060 2038 1116
rect 1974 1056 2038 1060
rect 2054 1116 2118 1120
rect 2054 1060 2058 1116
rect 2058 1060 2114 1116
rect 2114 1060 2118 1116
rect 2054 1056 2118 1060
rect 2134 1116 2198 1120
rect 2134 1060 2138 1116
rect 2138 1060 2194 1116
rect 2194 1060 2198 1116
rect 2134 1056 2198 1060
rect 2837 1116 2901 1120
rect 2837 1060 2841 1116
rect 2841 1060 2897 1116
rect 2897 1060 2901 1116
rect 2837 1056 2901 1060
rect 2917 1116 2981 1120
rect 2917 1060 2921 1116
rect 2921 1060 2977 1116
rect 2977 1060 2981 1116
rect 2917 1056 2981 1060
rect 2997 1116 3061 1120
rect 2997 1060 3001 1116
rect 3001 1060 3057 1116
rect 3057 1060 3061 1116
rect 2997 1056 3061 1060
rect 3077 1116 3141 1120
rect 3077 1060 3081 1116
rect 3081 1060 3137 1116
rect 3137 1060 3141 1116
rect 3077 1056 3141 1060
rect 3780 1116 3844 1120
rect 3780 1060 3784 1116
rect 3784 1060 3840 1116
rect 3840 1060 3844 1116
rect 3780 1056 3844 1060
rect 3860 1116 3924 1120
rect 3860 1060 3864 1116
rect 3864 1060 3920 1116
rect 3920 1060 3924 1116
rect 3860 1056 3924 1060
rect 3940 1116 4004 1120
rect 3940 1060 3944 1116
rect 3944 1060 4000 1116
rect 4000 1060 4004 1116
rect 3940 1056 4004 1060
rect 4020 1116 4084 1120
rect 4020 1060 4024 1116
rect 4024 1060 4080 1116
rect 4080 1060 4084 1116
rect 4020 1056 4084 1060
rect 4723 1116 4787 1120
rect 4723 1060 4727 1116
rect 4727 1060 4783 1116
rect 4783 1060 4787 1116
rect 4723 1056 4787 1060
rect 4803 1116 4867 1120
rect 4803 1060 4807 1116
rect 4807 1060 4863 1116
rect 4863 1060 4867 1116
rect 4803 1056 4867 1060
rect 4883 1116 4947 1120
rect 4883 1060 4887 1116
rect 4887 1060 4943 1116
rect 4943 1060 4947 1116
rect 4883 1056 4947 1060
rect 4963 1116 5027 1120
rect 4963 1060 4967 1116
rect 4967 1060 5023 1116
rect 5023 1060 5027 1116
rect 4963 1056 5027 1060
<< metal4 >>
rect 1415 22336 1735 22896
rect 1415 22272 1423 22336
rect 1487 22272 1503 22336
rect 1567 22272 1583 22336
rect 1647 22272 1663 22336
rect 1727 22272 1735 22336
rect 1415 21248 1735 22272
rect 1415 21184 1423 21248
rect 1487 21184 1503 21248
rect 1567 21184 1583 21248
rect 1647 21184 1663 21248
rect 1727 21184 1735 21248
rect 1415 20160 1735 21184
rect 1415 20096 1423 20160
rect 1487 20096 1503 20160
rect 1567 20096 1583 20160
rect 1647 20096 1663 20160
rect 1727 20096 1735 20160
rect 1415 19072 1735 20096
rect 1415 19008 1423 19072
rect 1487 19008 1503 19072
rect 1567 19008 1583 19072
rect 1647 19008 1663 19072
rect 1727 19008 1735 19072
rect 1415 17984 1735 19008
rect 1415 17920 1423 17984
rect 1487 17920 1503 17984
rect 1567 17920 1583 17984
rect 1647 17920 1663 17984
rect 1727 17920 1735 17984
rect 1415 16896 1735 17920
rect 1415 16832 1423 16896
rect 1487 16832 1503 16896
rect 1567 16832 1583 16896
rect 1647 16832 1663 16896
rect 1727 16832 1735 16896
rect 1415 15808 1735 16832
rect 1415 15744 1423 15808
rect 1487 15744 1503 15808
rect 1567 15744 1583 15808
rect 1647 15744 1663 15808
rect 1727 15744 1735 15808
rect 1415 14720 1735 15744
rect 1415 14656 1423 14720
rect 1487 14656 1503 14720
rect 1567 14656 1583 14720
rect 1647 14656 1663 14720
rect 1727 14656 1735 14720
rect 1415 13632 1735 14656
rect 1415 13568 1423 13632
rect 1487 13568 1503 13632
rect 1567 13568 1583 13632
rect 1647 13568 1663 13632
rect 1727 13568 1735 13632
rect 1415 12544 1735 13568
rect 1415 12480 1423 12544
rect 1487 12480 1503 12544
rect 1567 12480 1583 12544
rect 1647 12480 1663 12544
rect 1727 12480 1735 12544
rect 1415 11456 1735 12480
rect 1415 11392 1423 11456
rect 1487 11392 1503 11456
rect 1567 11392 1583 11456
rect 1647 11392 1663 11456
rect 1727 11392 1735 11456
rect 1415 10368 1735 11392
rect 1415 10304 1423 10368
rect 1487 10304 1503 10368
rect 1567 10304 1583 10368
rect 1647 10304 1663 10368
rect 1727 10304 1735 10368
rect 1415 9280 1735 10304
rect 1415 9216 1423 9280
rect 1487 9216 1503 9280
rect 1567 9216 1583 9280
rect 1647 9216 1663 9280
rect 1727 9216 1735 9280
rect 1415 8192 1735 9216
rect 1415 8128 1423 8192
rect 1487 8128 1503 8192
rect 1567 8128 1583 8192
rect 1647 8128 1663 8192
rect 1727 8128 1735 8192
rect 1415 7104 1735 8128
rect 1415 7040 1423 7104
rect 1487 7040 1503 7104
rect 1567 7040 1583 7104
rect 1647 7040 1663 7104
rect 1727 7040 1735 7104
rect 1415 6016 1735 7040
rect 1415 5952 1423 6016
rect 1487 5952 1503 6016
rect 1567 5952 1583 6016
rect 1647 5952 1663 6016
rect 1727 5952 1735 6016
rect 1415 4928 1735 5952
rect 1415 4864 1423 4928
rect 1487 4864 1503 4928
rect 1567 4864 1583 4928
rect 1647 4864 1663 4928
rect 1727 4864 1735 4928
rect 1415 3840 1735 4864
rect 1415 3776 1423 3840
rect 1487 3776 1503 3840
rect 1567 3776 1583 3840
rect 1647 3776 1663 3840
rect 1727 3776 1735 3840
rect 1415 2752 1735 3776
rect 1415 2688 1423 2752
rect 1487 2688 1503 2752
rect 1567 2688 1583 2752
rect 1647 2688 1663 2752
rect 1727 2688 1735 2752
rect 1415 1664 1735 2688
rect 1415 1600 1423 1664
rect 1487 1600 1503 1664
rect 1567 1600 1583 1664
rect 1647 1600 1663 1664
rect 1727 1600 1735 1664
rect 1415 1040 1735 1600
rect 1886 22880 2206 22896
rect 1886 22816 1894 22880
rect 1958 22816 1974 22880
rect 2038 22816 2054 22880
rect 2118 22816 2134 22880
rect 2198 22816 2206 22880
rect 1886 21792 2206 22816
rect 1886 21728 1894 21792
rect 1958 21728 1974 21792
rect 2038 21728 2054 21792
rect 2118 21728 2134 21792
rect 2198 21728 2206 21792
rect 1886 20704 2206 21728
rect 1886 20640 1894 20704
rect 1958 20640 1974 20704
rect 2038 20640 2054 20704
rect 2118 20640 2134 20704
rect 2198 20640 2206 20704
rect 1886 19616 2206 20640
rect 1886 19552 1894 19616
rect 1958 19552 1974 19616
rect 2038 19552 2054 19616
rect 2118 19552 2134 19616
rect 2198 19552 2206 19616
rect 1886 18528 2206 19552
rect 1886 18464 1894 18528
rect 1958 18464 1974 18528
rect 2038 18464 2054 18528
rect 2118 18464 2134 18528
rect 2198 18464 2206 18528
rect 1886 17440 2206 18464
rect 1886 17376 1894 17440
rect 1958 17376 1974 17440
rect 2038 17376 2054 17440
rect 2118 17376 2134 17440
rect 2198 17376 2206 17440
rect 1886 16352 2206 17376
rect 1886 16288 1894 16352
rect 1958 16288 1974 16352
rect 2038 16288 2054 16352
rect 2118 16288 2134 16352
rect 2198 16288 2206 16352
rect 1886 15264 2206 16288
rect 1886 15200 1894 15264
rect 1958 15200 1974 15264
rect 2038 15200 2054 15264
rect 2118 15200 2134 15264
rect 2198 15200 2206 15264
rect 1886 14176 2206 15200
rect 1886 14112 1894 14176
rect 1958 14112 1974 14176
rect 2038 14112 2054 14176
rect 2118 14112 2134 14176
rect 2198 14112 2206 14176
rect 1886 13088 2206 14112
rect 1886 13024 1894 13088
rect 1958 13024 1974 13088
rect 2038 13024 2054 13088
rect 2118 13024 2134 13088
rect 2198 13024 2206 13088
rect 1886 12000 2206 13024
rect 1886 11936 1894 12000
rect 1958 11936 1974 12000
rect 2038 11936 2054 12000
rect 2118 11936 2134 12000
rect 2198 11936 2206 12000
rect 1886 10912 2206 11936
rect 1886 10848 1894 10912
rect 1958 10848 1974 10912
rect 2038 10848 2054 10912
rect 2118 10848 2134 10912
rect 2198 10848 2206 10912
rect 1886 9824 2206 10848
rect 1886 9760 1894 9824
rect 1958 9760 1974 9824
rect 2038 9760 2054 9824
rect 2118 9760 2134 9824
rect 2198 9760 2206 9824
rect 1886 8736 2206 9760
rect 1886 8672 1894 8736
rect 1958 8672 1974 8736
rect 2038 8672 2054 8736
rect 2118 8672 2134 8736
rect 2198 8672 2206 8736
rect 1886 7648 2206 8672
rect 1886 7584 1894 7648
rect 1958 7584 1974 7648
rect 2038 7584 2054 7648
rect 2118 7584 2134 7648
rect 2198 7584 2206 7648
rect 1886 6560 2206 7584
rect 1886 6496 1894 6560
rect 1958 6496 1974 6560
rect 2038 6496 2054 6560
rect 2118 6496 2134 6560
rect 2198 6496 2206 6560
rect 1886 5472 2206 6496
rect 1886 5408 1894 5472
rect 1958 5408 1974 5472
rect 2038 5408 2054 5472
rect 2118 5408 2134 5472
rect 2198 5408 2206 5472
rect 1886 4384 2206 5408
rect 1886 4320 1894 4384
rect 1958 4320 1974 4384
rect 2038 4320 2054 4384
rect 2118 4320 2134 4384
rect 2198 4320 2206 4384
rect 1886 3296 2206 4320
rect 1886 3232 1894 3296
rect 1958 3232 1974 3296
rect 2038 3232 2054 3296
rect 2118 3232 2134 3296
rect 2198 3232 2206 3296
rect 1886 2208 2206 3232
rect 1886 2144 1894 2208
rect 1958 2144 1974 2208
rect 2038 2144 2054 2208
rect 2118 2144 2134 2208
rect 2198 2144 2206 2208
rect 1886 1120 2206 2144
rect 1886 1056 1894 1120
rect 1958 1056 1974 1120
rect 2038 1056 2054 1120
rect 2118 1056 2134 1120
rect 2198 1056 2206 1120
rect 1886 1040 2206 1056
rect 2358 22336 2678 22896
rect 2358 22272 2366 22336
rect 2430 22272 2446 22336
rect 2510 22272 2526 22336
rect 2590 22272 2606 22336
rect 2670 22272 2678 22336
rect 2358 21248 2678 22272
rect 2358 21184 2366 21248
rect 2430 21184 2446 21248
rect 2510 21184 2526 21248
rect 2590 21184 2606 21248
rect 2670 21184 2678 21248
rect 2358 20160 2678 21184
rect 2358 20096 2366 20160
rect 2430 20096 2446 20160
rect 2510 20096 2526 20160
rect 2590 20096 2606 20160
rect 2670 20096 2678 20160
rect 2358 19072 2678 20096
rect 2358 19008 2366 19072
rect 2430 19008 2446 19072
rect 2510 19008 2526 19072
rect 2590 19008 2606 19072
rect 2670 19008 2678 19072
rect 2358 17984 2678 19008
rect 2358 17920 2366 17984
rect 2430 17920 2446 17984
rect 2510 17920 2526 17984
rect 2590 17920 2606 17984
rect 2670 17920 2678 17984
rect 2358 16896 2678 17920
rect 2358 16832 2366 16896
rect 2430 16832 2446 16896
rect 2510 16832 2526 16896
rect 2590 16832 2606 16896
rect 2670 16832 2678 16896
rect 2358 15808 2678 16832
rect 2358 15744 2366 15808
rect 2430 15744 2446 15808
rect 2510 15744 2526 15808
rect 2590 15744 2606 15808
rect 2670 15744 2678 15808
rect 2358 14720 2678 15744
rect 2358 14656 2366 14720
rect 2430 14656 2446 14720
rect 2510 14656 2526 14720
rect 2590 14656 2606 14720
rect 2670 14656 2678 14720
rect 2358 13632 2678 14656
rect 2358 13568 2366 13632
rect 2430 13568 2446 13632
rect 2510 13568 2526 13632
rect 2590 13568 2606 13632
rect 2670 13568 2678 13632
rect 2358 12544 2678 13568
rect 2358 12480 2366 12544
rect 2430 12480 2446 12544
rect 2510 12480 2526 12544
rect 2590 12480 2606 12544
rect 2670 12480 2678 12544
rect 2358 11456 2678 12480
rect 2358 11392 2366 11456
rect 2430 11392 2446 11456
rect 2510 11392 2526 11456
rect 2590 11392 2606 11456
rect 2670 11392 2678 11456
rect 2358 10368 2678 11392
rect 2358 10304 2366 10368
rect 2430 10304 2446 10368
rect 2510 10304 2526 10368
rect 2590 10304 2606 10368
rect 2670 10304 2678 10368
rect 2358 9280 2678 10304
rect 2358 9216 2366 9280
rect 2430 9216 2446 9280
rect 2510 9216 2526 9280
rect 2590 9216 2606 9280
rect 2670 9216 2678 9280
rect 2358 8192 2678 9216
rect 2358 8128 2366 8192
rect 2430 8128 2446 8192
rect 2510 8128 2526 8192
rect 2590 8128 2606 8192
rect 2670 8128 2678 8192
rect 2358 7104 2678 8128
rect 2358 7040 2366 7104
rect 2430 7040 2446 7104
rect 2510 7040 2526 7104
rect 2590 7040 2606 7104
rect 2670 7040 2678 7104
rect 2358 6016 2678 7040
rect 2358 5952 2366 6016
rect 2430 5952 2446 6016
rect 2510 5952 2526 6016
rect 2590 5952 2606 6016
rect 2670 5952 2678 6016
rect 2358 4928 2678 5952
rect 2358 4864 2366 4928
rect 2430 4864 2446 4928
rect 2510 4864 2526 4928
rect 2590 4864 2606 4928
rect 2670 4864 2678 4928
rect 2358 3840 2678 4864
rect 2358 3776 2366 3840
rect 2430 3776 2446 3840
rect 2510 3776 2526 3840
rect 2590 3776 2606 3840
rect 2670 3776 2678 3840
rect 2358 2752 2678 3776
rect 2358 2688 2366 2752
rect 2430 2688 2446 2752
rect 2510 2688 2526 2752
rect 2590 2688 2606 2752
rect 2670 2688 2678 2752
rect 2358 1664 2678 2688
rect 2358 1600 2366 1664
rect 2430 1600 2446 1664
rect 2510 1600 2526 1664
rect 2590 1600 2606 1664
rect 2670 1600 2678 1664
rect 2358 1040 2678 1600
rect 2829 22880 3149 22896
rect 2829 22816 2837 22880
rect 2901 22816 2917 22880
rect 2981 22816 2997 22880
rect 3061 22816 3077 22880
rect 3141 22816 3149 22880
rect 2829 21792 3149 22816
rect 2829 21728 2837 21792
rect 2901 21728 2917 21792
rect 2981 21728 2997 21792
rect 3061 21728 3077 21792
rect 3141 21728 3149 21792
rect 2829 20704 3149 21728
rect 2829 20640 2837 20704
rect 2901 20640 2917 20704
rect 2981 20640 2997 20704
rect 3061 20640 3077 20704
rect 3141 20640 3149 20704
rect 2829 19616 3149 20640
rect 2829 19552 2837 19616
rect 2901 19552 2917 19616
rect 2981 19552 2997 19616
rect 3061 19552 3077 19616
rect 3141 19552 3149 19616
rect 2829 18528 3149 19552
rect 2829 18464 2837 18528
rect 2901 18464 2917 18528
rect 2981 18464 2997 18528
rect 3061 18464 3077 18528
rect 3141 18464 3149 18528
rect 2829 17440 3149 18464
rect 2829 17376 2837 17440
rect 2901 17376 2917 17440
rect 2981 17376 2997 17440
rect 3061 17376 3077 17440
rect 3141 17376 3149 17440
rect 2829 16352 3149 17376
rect 2829 16288 2837 16352
rect 2901 16288 2917 16352
rect 2981 16288 2997 16352
rect 3061 16288 3077 16352
rect 3141 16288 3149 16352
rect 2829 15264 3149 16288
rect 2829 15200 2837 15264
rect 2901 15200 2917 15264
rect 2981 15200 2997 15264
rect 3061 15200 3077 15264
rect 3141 15200 3149 15264
rect 2829 14176 3149 15200
rect 2829 14112 2837 14176
rect 2901 14112 2917 14176
rect 2981 14112 2997 14176
rect 3061 14112 3077 14176
rect 3141 14112 3149 14176
rect 2829 13088 3149 14112
rect 2829 13024 2837 13088
rect 2901 13024 2917 13088
rect 2981 13024 2997 13088
rect 3061 13024 3077 13088
rect 3141 13024 3149 13088
rect 2829 12000 3149 13024
rect 2829 11936 2837 12000
rect 2901 11936 2917 12000
rect 2981 11936 2997 12000
rect 3061 11936 3077 12000
rect 3141 11936 3149 12000
rect 2829 10912 3149 11936
rect 2829 10848 2837 10912
rect 2901 10848 2917 10912
rect 2981 10848 2997 10912
rect 3061 10848 3077 10912
rect 3141 10848 3149 10912
rect 2829 9824 3149 10848
rect 2829 9760 2837 9824
rect 2901 9760 2917 9824
rect 2981 9760 2997 9824
rect 3061 9760 3077 9824
rect 3141 9760 3149 9824
rect 2829 8736 3149 9760
rect 2829 8672 2837 8736
rect 2901 8672 2917 8736
rect 2981 8672 2997 8736
rect 3061 8672 3077 8736
rect 3141 8672 3149 8736
rect 2829 7648 3149 8672
rect 2829 7584 2837 7648
rect 2901 7584 2917 7648
rect 2981 7584 2997 7648
rect 3061 7584 3077 7648
rect 3141 7584 3149 7648
rect 2829 6560 3149 7584
rect 2829 6496 2837 6560
rect 2901 6496 2917 6560
rect 2981 6496 2997 6560
rect 3061 6496 3077 6560
rect 3141 6496 3149 6560
rect 2829 5472 3149 6496
rect 2829 5408 2837 5472
rect 2901 5408 2917 5472
rect 2981 5408 2997 5472
rect 3061 5408 3077 5472
rect 3141 5408 3149 5472
rect 2829 4384 3149 5408
rect 2829 4320 2837 4384
rect 2901 4320 2917 4384
rect 2981 4320 2997 4384
rect 3061 4320 3077 4384
rect 3141 4320 3149 4384
rect 2829 3296 3149 4320
rect 2829 3232 2837 3296
rect 2901 3232 2917 3296
rect 2981 3232 2997 3296
rect 3061 3232 3077 3296
rect 3141 3232 3149 3296
rect 2829 2208 3149 3232
rect 2829 2144 2837 2208
rect 2901 2144 2917 2208
rect 2981 2144 2997 2208
rect 3061 2144 3077 2208
rect 3141 2144 3149 2208
rect 2829 1120 3149 2144
rect 2829 1056 2837 1120
rect 2901 1056 2917 1120
rect 2981 1056 2997 1120
rect 3061 1056 3077 1120
rect 3141 1056 3149 1120
rect 2829 1040 3149 1056
rect 3301 22336 3621 22896
rect 3301 22272 3309 22336
rect 3373 22272 3389 22336
rect 3453 22272 3469 22336
rect 3533 22272 3549 22336
rect 3613 22272 3621 22336
rect 3301 21248 3621 22272
rect 3301 21184 3309 21248
rect 3373 21184 3389 21248
rect 3453 21184 3469 21248
rect 3533 21184 3549 21248
rect 3613 21184 3621 21248
rect 3301 20160 3621 21184
rect 3301 20096 3309 20160
rect 3373 20096 3389 20160
rect 3453 20096 3469 20160
rect 3533 20096 3549 20160
rect 3613 20096 3621 20160
rect 3301 19072 3621 20096
rect 3301 19008 3309 19072
rect 3373 19008 3389 19072
rect 3453 19008 3469 19072
rect 3533 19008 3549 19072
rect 3613 19008 3621 19072
rect 3301 17984 3621 19008
rect 3301 17920 3309 17984
rect 3373 17920 3389 17984
rect 3453 17920 3469 17984
rect 3533 17920 3549 17984
rect 3613 17920 3621 17984
rect 3301 16896 3621 17920
rect 3301 16832 3309 16896
rect 3373 16832 3389 16896
rect 3453 16832 3469 16896
rect 3533 16832 3549 16896
rect 3613 16832 3621 16896
rect 3301 15808 3621 16832
rect 3301 15744 3309 15808
rect 3373 15744 3389 15808
rect 3453 15744 3469 15808
rect 3533 15744 3549 15808
rect 3613 15744 3621 15808
rect 3301 14720 3621 15744
rect 3301 14656 3309 14720
rect 3373 14656 3389 14720
rect 3453 14656 3469 14720
rect 3533 14656 3549 14720
rect 3613 14656 3621 14720
rect 3301 13632 3621 14656
rect 3301 13568 3309 13632
rect 3373 13568 3389 13632
rect 3453 13568 3469 13632
rect 3533 13568 3549 13632
rect 3613 13568 3621 13632
rect 3301 12544 3621 13568
rect 3301 12480 3309 12544
rect 3373 12480 3389 12544
rect 3453 12480 3469 12544
rect 3533 12480 3549 12544
rect 3613 12480 3621 12544
rect 3301 11456 3621 12480
rect 3301 11392 3309 11456
rect 3373 11392 3389 11456
rect 3453 11392 3469 11456
rect 3533 11392 3549 11456
rect 3613 11392 3621 11456
rect 3301 10368 3621 11392
rect 3301 10304 3309 10368
rect 3373 10304 3389 10368
rect 3453 10304 3469 10368
rect 3533 10304 3549 10368
rect 3613 10304 3621 10368
rect 3301 9280 3621 10304
rect 3301 9216 3309 9280
rect 3373 9216 3389 9280
rect 3453 9216 3469 9280
rect 3533 9216 3549 9280
rect 3613 9216 3621 9280
rect 3301 8192 3621 9216
rect 3301 8128 3309 8192
rect 3373 8128 3389 8192
rect 3453 8128 3469 8192
rect 3533 8128 3549 8192
rect 3613 8128 3621 8192
rect 3301 7104 3621 8128
rect 3301 7040 3309 7104
rect 3373 7040 3389 7104
rect 3453 7040 3469 7104
rect 3533 7040 3549 7104
rect 3613 7040 3621 7104
rect 3301 6016 3621 7040
rect 3301 5952 3309 6016
rect 3373 5952 3389 6016
rect 3453 5952 3469 6016
rect 3533 5952 3549 6016
rect 3613 5952 3621 6016
rect 3301 4928 3621 5952
rect 3301 4864 3309 4928
rect 3373 4864 3389 4928
rect 3453 4864 3469 4928
rect 3533 4864 3549 4928
rect 3613 4864 3621 4928
rect 3301 3840 3621 4864
rect 3301 3776 3309 3840
rect 3373 3776 3389 3840
rect 3453 3776 3469 3840
rect 3533 3776 3549 3840
rect 3613 3776 3621 3840
rect 3301 2752 3621 3776
rect 3301 2688 3309 2752
rect 3373 2688 3389 2752
rect 3453 2688 3469 2752
rect 3533 2688 3549 2752
rect 3613 2688 3621 2752
rect 3301 1664 3621 2688
rect 3301 1600 3309 1664
rect 3373 1600 3389 1664
rect 3453 1600 3469 1664
rect 3533 1600 3549 1664
rect 3613 1600 3621 1664
rect 3301 1040 3621 1600
rect 3772 22880 4092 22896
rect 3772 22816 3780 22880
rect 3844 22816 3860 22880
rect 3924 22816 3940 22880
rect 4004 22816 4020 22880
rect 4084 22816 4092 22880
rect 3772 21792 4092 22816
rect 3772 21728 3780 21792
rect 3844 21728 3860 21792
rect 3924 21728 3940 21792
rect 4004 21728 4020 21792
rect 4084 21728 4092 21792
rect 3772 20704 4092 21728
rect 3772 20640 3780 20704
rect 3844 20640 3860 20704
rect 3924 20640 3940 20704
rect 4004 20640 4020 20704
rect 4084 20640 4092 20704
rect 3772 19616 4092 20640
rect 3772 19552 3780 19616
rect 3844 19552 3860 19616
rect 3924 19552 3940 19616
rect 4004 19552 4020 19616
rect 4084 19552 4092 19616
rect 3772 18528 4092 19552
rect 3772 18464 3780 18528
rect 3844 18464 3860 18528
rect 3924 18464 3940 18528
rect 4004 18464 4020 18528
rect 4084 18464 4092 18528
rect 3772 17440 4092 18464
rect 3772 17376 3780 17440
rect 3844 17376 3860 17440
rect 3924 17376 3940 17440
rect 4004 17376 4020 17440
rect 4084 17376 4092 17440
rect 3772 16352 4092 17376
rect 3772 16288 3780 16352
rect 3844 16288 3860 16352
rect 3924 16288 3940 16352
rect 4004 16288 4020 16352
rect 4084 16288 4092 16352
rect 3772 15264 4092 16288
rect 3772 15200 3780 15264
rect 3844 15200 3860 15264
rect 3924 15200 3940 15264
rect 4004 15200 4020 15264
rect 4084 15200 4092 15264
rect 3772 14176 4092 15200
rect 3772 14112 3780 14176
rect 3844 14112 3860 14176
rect 3924 14112 3940 14176
rect 4004 14112 4020 14176
rect 4084 14112 4092 14176
rect 3772 13088 4092 14112
rect 3772 13024 3780 13088
rect 3844 13024 3860 13088
rect 3924 13024 3940 13088
rect 4004 13024 4020 13088
rect 4084 13024 4092 13088
rect 3772 12000 4092 13024
rect 3772 11936 3780 12000
rect 3844 11936 3860 12000
rect 3924 11936 3940 12000
rect 4004 11936 4020 12000
rect 4084 11936 4092 12000
rect 3772 10912 4092 11936
rect 3772 10848 3780 10912
rect 3844 10848 3860 10912
rect 3924 10848 3940 10912
rect 4004 10848 4020 10912
rect 4084 10848 4092 10912
rect 3772 9824 4092 10848
rect 3772 9760 3780 9824
rect 3844 9760 3860 9824
rect 3924 9760 3940 9824
rect 4004 9760 4020 9824
rect 4084 9760 4092 9824
rect 3772 8736 4092 9760
rect 3772 8672 3780 8736
rect 3844 8672 3860 8736
rect 3924 8672 3940 8736
rect 4004 8672 4020 8736
rect 4084 8672 4092 8736
rect 3772 7648 4092 8672
rect 3772 7584 3780 7648
rect 3844 7584 3860 7648
rect 3924 7584 3940 7648
rect 4004 7584 4020 7648
rect 4084 7584 4092 7648
rect 3772 6560 4092 7584
rect 3772 6496 3780 6560
rect 3844 6496 3860 6560
rect 3924 6496 3940 6560
rect 4004 6496 4020 6560
rect 4084 6496 4092 6560
rect 3772 5472 4092 6496
rect 3772 5408 3780 5472
rect 3844 5408 3860 5472
rect 3924 5408 3940 5472
rect 4004 5408 4020 5472
rect 4084 5408 4092 5472
rect 3772 4384 4092 5408
rect 3772 4320 3780 4384
rect 3844 4320 3860 4384
rect 3924 4320 3940 4384
rect 4004 4320 4020 4384
rect 4084 4320 4092 4384
rect 3772 3296 4092 4320
rect 3772 3232 3780 3296
rect 3844 3232 3860 3296
rect 3924 3232 3940 3296
rect 4004 3232 4020 3296
rect 4084 3232 4092 3296
rect 3772 2208 4092 3232
rect 3772 2144 3780 2208
rect 3844 2144 3860 2208
rect 3924 2144 3940 2208
rect 4004 2144 4020 2208
rect 4084 2144 4092 2208
rect 3772 1120 4092 2144
rect 3772 1056 3780 1120
rect 3844 1056 3860 1120
rect 3924 1056 3940 1120
rect 4004 1056 4020 1120
rect 4084 1056 4092 1120
rect 3772 1040 4092 1056
rect 4244 22336 4564 22896
rect 4244 22272 4252 22336
rect 4316 22272 4332 22336
rect 4396 22272 4412 22336
rect 4476 22272 4492 22336
rect 4556 22272 4564 22336
rect 4244 21248 4564 22272
rect 4244 21184 4252 21248
rect 4316 21184 4332 21248
rect 4396 21184 4412 21248
rect 4476 21184 4492 21248
rect 4556 21184 4564 21248
rect 4244 20160 4564 21184
rect 4244 20096 4252 20160
rect 4316 20096 4332 20160
rect 4396 20096 4412 20160
rect 4476 20096 4492 20160
rect 4556 20096 4564 20160
rect 4244 19072 4564 20096
rect 4244 19008 4252 19072
rect 4316 19008 4332 19072
rect 4396 19008 4412 19072
rect 4476 19008 4492 19072
rect 4556 19008 4564 19072
rect 4244 17984 4564 19008
rect 4244 17920 4252 17984
rect 4316 17920 4332 17984
rect 4396 17920 4412 17984
rect 4476 17920 4492 17984
rect 4556 17920 4564 17984
rect 4244 16896 4564 17920
rect 4244 16832 4252 16896
rect 4316 16832 4332 16896
rect 4396 16832 4412 16896
rect 4476 16832 4492 16896
rect 4556 16832 4564 16896
rect 4244 15808 4564 16832
rect 4244 15744 4252 15808
rect 4316 15744 4332 15808
rect 4396 15744 4412 15808
rect 4476 15744 4492 15808
rect 4556 15744 4564 15808
rect 4244 14720 4564 15744
rect 4244 14656 4252 14720
rect 4316 14656 4332 14720
rect 4396 14656 4412 14720
rect 4476 14656 4492 14720
rect 4556 14656 4564 14720
rect 4244 13632 4564 14656
rect 4244 13568 4252 13632
rect 4316 13568 4332 13632
rect 4396 13568 4412 13632
rect 4476 13568 4492 13632
rect 4556 13568 4564 13632
rect 4244 12544 4564 13568
rect 4244 12480 4252 12544
rect 4316 12480 4332 12544
rect 4396 12480 4412 12544
rect 4476 12480 4492 12544
rect 4556 12480 4564 12544
rect 4244 11456 4564 12480
rect 4244 11392 4252 11456
rect 4316 11392 4332 11456
rect 4396 11392 4412 11456
rect 4476 11392 4492 11456
rect 4556 11392 4564 11456
rect 4244 10368 4564 11392
rect 4244 10304 4252 10368
rect 4316 10304 4332 10368
rect 4396 10304 4412 10368
rect 4476 10304 4492 10368
rect 4556 10304 4564 10368
rect 4244 9280 4564 10304
rect 4244 9216 4252 9280
rect 4316 9216 4332 9280
rect 4396 9216 4412 9280
rect 4476 9216 4492 9280
rect 4556 9216 4564 9280
rect 4244 8192 4564 9216
rect 4244 8128 4252 8192
rect 4316 8128 4332 8192
rect 4396 8128 4412 8192
rect 4476 8128 4492 8192
rect 4556 8128 4564 8192
rect 4244 7104 4564 8128
rect 4244 7040 4252 7104
rect 4316 7040 4332 7104
rect 4396 7040 4412 7104
rect 4476 7040 4492 7104
rect 4556 7040 4564 7104
rect 4244 6016 4564 7040
rect 4244 5952 4252 6016
rect 4316 5952 4332 6016
rect 4396 5952 4412 6016
rect 4476 5952 4492 6016
rect 4556 5952 4564 6016
rect 4244 4928 4564 5952
rect 4244 4864 4252 4928
rect 4316 4864 4332 4928
rect 4396 4864 4412 4928
rect 4476 4864 4492 4928
rect 4556 4864 4564 4928
rect 4244 3840 4564 4864
rect 4244 3776 4252 3840
rect 4316 3776 4332 3840
rect 4396 3776 4412 3840
rect 4476 3776 4492 3840
rect 4556 3776 4564 3840
rect 4244 2752 4564 3776
rect 4244 2688 4252 2752
rect 4316 2688 4332 2752
rect 4396 2688 4412 2752
rect 4476 2688 4492 2752
rect 4556 2688 4564 2752
rect 4244 1664 4564 2688
rect 4244 1600 4252 1664
rect 4316 1600 4332 1664
rect 4396 1600 4412 1664
rect 4476 1600 4492 1664
rect 4556 1600 4564 1664
rect 4244 1040 4564 1600
rect 4715 22880 5035 22896
rect 4715 22816 4723 22880
rect 4787 22816 4803 22880
rect 4867 22816 4883 22880
rect 4947 22816 4963 22880
rect 5027 22816 5035 22880
rect 4715 21792 5035 22816
rect 4715 21728 4723 21792
rect 4787 21728 4803 21792
rect 4867 21728 4883 21792
rect 4947 21728 4963 21792
rect 5027 21728 5035 21792
rect 4715 20704 5035 21728
rect 4715 20640 4723 20704
rect 4787 20640 4803 20704
rect 4867 20640 4883 20704
rect 4947 20640 4963 20704
rect 5027 20640 5035 20704
rect 4715 19616 5035 20640
rect 4715 19552 4723 19616
rect 4787 19552 4803 19616
rect 4867 19552 4883 19616
rect 4947 19552 4963 19616
rect 5027 19552 5035 19616
rect 4715 18528 5035 19552
rect 4715 18464 4723 18528
rect 4787 18464 4803 18528
rect 4867 18464 4883 18528
rect 4947 18464 4963 18528
rect 5027 18464 5035 18528
rect 4715 17440 5035 18464
rect 4715 17376 4723 17440
rect 4787 17376 4803 17440
rect 4867 17376 4883 17440
rect 4947 17376 4963 17440
rect 5027 17376 5035 17440
rect 4715 16352 5035 17376
rect 4715 16288 4723 16352
rect 4787 16288 4803 16352
rect 4867 16288 4883 16352
rect 4947 16288 4963 16352
rect 5027 16288 5035 16352
rect 4715 15264 5035 16288
rect 4715 15200 4723 15264
rect 4787 15200 4803 15264
rect 4867 15200 4883 15264
rect 4947 15200 4963 15264
rect 5027 15200 5035 15264
rect 4715 14176 5035 15200
rect 4715 14112 4723 14176
rect 4787 14112 4803 14176
rect 4867 14112 4883 14176
rect 4947 14112 4963 14176
rect 5027 14112 5035 14176
rect 4715 13088 5035 14112
rect 4715 13024 4723 13088
rect 4787 13024 4803 13088
rect 4867 13024 4883 13088
rect 4947 13024 4963 13088
rect 5027 13024 5035 13088
rect 4715 12000 5035 13024
rect 4715 11936 4723 12000
rect 4787 11936 4803 12000
rect 4867 11936 4883 12000
rect 4947 11936 4963 12000
rect 5027 11936 5035 12000
rect 4715 10912 5035 11936
rect 4715 10848 4723 10912
rect 4787 10848 4803 10912
rect 4867 10848 4883 10912
rect 4947 10848 4963 10912
rect 5027 10848 5035 10912
rect 4715 9824 5035 10848
rect 4715 9760 4723 9824
rect 4787 9760 4803 9824
rect 4867 9760 4883 9824
rect 4947 9760 4963 9824
rect 5027 9760 5035 9824
rect 4715 8736 5035 9760
rect 4715 8672 4723 8736
rect 4787 8672 4803 8736
rect 4867 8672 4883 8736
rect 4947 8672 4963 8736
rect 5027 8672 5035 8736
rect 4715 7648 5035 8672
rect 4715 7584 4723 7648
rect 4787 7584 4803 7648
rect 4867 7584 4883 7648
rect 4947 7584 4963 7648
rect 5027 7584 5035 7648
rect 4715 6560 5035 7584
rect 4715 6496 4723 6560
rect 4787 6496 4803 6560
rect 4867 6496 4883 6560
rect 4947 6496 4963 6560
rect 5027 6496 5035 6560
rect 4715 5472 5035 6496
rect 4715 5408 4723 5472
rect 4787 5408 4803 5472
rect 4867 5408 4883 5472
rect 4947 5408 4963 5472
rect 5027 5408 5035 5472
rect 4715 4384 5035 5408
rect 4715 4320 4723 4384
rect 4787 4320 4803 4384
rect 4867 4320 4883 4384
rect 4947 4320 4963 4384
rect 5027 4320 5035 4384
rect 4715 3296 5035 4320
rect 4715 3232 4723 3296
rect 4787 3232 4803 3296
rect 4867 3232 4883 3296
rect 4947 3232 4963 3296
rect 5027 3232 5035 3296
rect 4715 2208 5035 3232
rect 4715 2144 4723 2208
rect 4787 2144 4803 2208
rect 4867 2144 4883 2208
rect 4947 2144 4963 2208
rect 5027 2144 5035 2208
rect 4715 1120 5035 2144
rect 4715 1056 4723 1120
rect 4787 1056 4803 1120
rect 4867 1056 4883 1120
rect 4947 1056 4963 1120
rect 5027 1056 5035 1120
rect 4715 1040 5035 1056
use sky130_ef_sc_hd__decap_12  FILLER_0_3 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 1380 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 2484 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 2852 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3496 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3772 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37
timestamp 1676037725
transform 1 0 4508 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_1_3 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 1380 0 -1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_1_16
timestamp 1676037725
transform 1 0 2576 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_34
timestamp 1676037725
transform 1 0 4232 0 -1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3
timestamp 1676037725
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_15
timestamp 1676037725
transform 1 0 2484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 1676037725
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_29
timestamp 1676037725
transform 1 0 3772 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_37
timestamp 1676037725
transform 1 0 4508 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3
timestamp 1676037725
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_15
timestamp 1676037725
transform 1 0 2484 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_23
timestamp 1676037725
transform 1 0 3220 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_36
timestamp 1676037725
transform 1 0 4416 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3
timestamp 1676037725
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_15
timestamp 1676037725
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1676037725
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_29
timestamp 1676037725
transform 1 0 3772 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_37
timestamp 1676037725
transform 1 0 4508 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3
timestamp 1676037725
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_15
timestamp 1676037725
transform 1 0 2484 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_23
timestamp 1676037725
transform 1 0 3220 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_36
timestamp 1676037725
transform 1 0 4416 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_6_3
timestamp 1676037725
transform 1 0 1380 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_6_11 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 2116 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_26
timestamp 1676037725
transform 1 0 3496 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_29
timestamp 1676037725
transform 1 0 3772 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_35
timestamp 1676037725
transform 1 0 4324 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_7_3
timestamp 1676037725
transform 1 0 1380 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_7
timestamp 1676037725
transform 1 0 1748 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_20
timestamp 1676037725
transform 1 0 2944 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_36
timestamp 1676037725
transform 1 0 4416 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_8_3
timestamp 1676037725
transform 1 0 1380 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_8_11
timestamp 1676037725
transform 1 0 2116 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_26
timestamp 1676037725
transform 1 0 3496 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_8_29
timestamp 1676037725
transform 1 0 3772 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_37
timestamp 1676037725
transform 1 0 4508 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_3
timestamp 1676037725
transform 1 0 1380 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_11
timestamp 1676037725
transform 1 0 2116 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_36
timestamp 1676037725
transform 1 0 4416 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_10_3
timestamp 1676037725
transform 1 0 1380 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_10_11
timestamp 1676037725
transform 1 0 2116 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_26
timestamp 1676037725
transform 1 0 3496 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_29
timestamp 1676037725
transform 1 0 3772 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_34
timestamp 1676037725
transform 1 0 4232 0 1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3
timestamp 1676037725
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_36
timestamp 1676037725
transform 1 0 4416 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_3
timestamp 1676037725
transform 1 0 1380 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_26
timestamp 1676037725
transform 1 0 3496 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_29
timestamp 1676037725
transform 1 0 3772 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_37
timestamp 1676037725
transform 1 0 4508 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3
timestamp 1676037725
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_36
timestamp 1676037725
transform 1 0 4416 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_3
timestamp 1676037725
transform 1 0 1380 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_26
timestamp 1676037725
transform 1 0 3496 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_14_29
timestamp 1676037725
transform 1 0 3772 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_37
timestamp 1676037725
transform 1 0 4508 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_3
timestamp 1676037725
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_15_36
timestamp 1676037725
transform 1 0 4416 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_3
timestamp 1676037725
transform 1 0 1380 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_26
timestamp 1676037725
transform 1 0 3496 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_16_29
timestamp 1676037725
transform 1 0 3772 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_37
timestamp 1676037725
transform 1 0 4508 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_3
timestamp 1676037725
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_36
timestamp 1676037725
transform 1 0 4416 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_3
timestamp 1676037725
transform 1 0 1380 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_18_11
timestamp 1676037725
transform 1 0 2116 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_26
timestamp 1676037725
transform 1 0 3496 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_29
timestamp 1676037725
transform 1 0 3772 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_37
timestamp 1676037725
transform 1 0 4508 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_3
timestamp 1676037725
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_19_36
timestamp 1676037725
transform 1 0 4416 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_3
timestamp 1676037725
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_15
timestamp 1676037725
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1676037725
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_29
timestamp 1676037725
transform 1 0 3772 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_37
timestamp 1676037725
transform 1 0 4508 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_3
timestamp 1676037725
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_15
timestamp 1676037725
transform 1 0 2484 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_27
timestamp 1676037725
transform 1 0 3588 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_35
timestamp 1676037725
transform 1 0 4324 0 -1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_22_3
timestamp 1676037725
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_15
timestamp 1676037725
transform 1 0 2484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 1676037725
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_29
timestamp 1676037725
transform 1 0 3772 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_37
timestamp 1676037725
transform 1 0 4508 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_3
timestamp 1676037725
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_15
timestamp 1676037725
transform 1 0 2484 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_27
timestamp 1676037725
transform 1 0 3588 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_23_35
timestamp 1676037725
transform 1 0 4324 0 -1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_24_3
timestamp 1676037725
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_15
timestamp 1676037725
transform 1 0 2484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1676037725
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_29
timestamp 1676037725
transform 1 0 3772 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_37
timestamp 1676037725
transform 1 0 4508 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_3
timestamp 1676037725
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_15
timestamp 1676037725
transform 1 0 2484 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_27
timestamp 1676037725
transform 1 0 3588 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_25_35
timestamp 1676037725
transform 1 0 4324 0 -1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_26_3
timestamp 1676037725
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_15
timestamp 1676037725
transform 1 0 2484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 1676037725
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_29
timestamp 1676037725
transform 1 0 3772 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_37
timestamp 1676037725
transform 1 0 4508 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_3
timestamp 1676037725
transform 1 0 1380 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_15
timestamp 1676037725
transform 1 0 2484 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_27
timestamp 1676037725
transform 1 0 3588 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_35
timestamp 1676037725
transform 1 0 4324 0 -1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_28_3
timestamp 1676037725
transform 1 0 1380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_15
timestamp 1676037725
transform 1 0 2484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_27
timestamp 1676037725
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_29
timestamp 1676037725
transform 1 0 3772 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_37
timestamp 1676037725
transform 1 0 4508 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_3
timestamp 1676037725
transform 1 0 1380 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_15
timestamp 1676037725
transform 1 0 2484 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_27
timestamp 1676037725
transform 1 0 3588 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_29_35
timestamp 1676037725
transform 1 0 4324 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_30_3
timestamp 1676037725
transform 1 0 1380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_15
timestamp 1676037725
transform 1 0 2484 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_27
timestamp 1676037725
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_29
timestamp 1676037725
transform 1 0 3772 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_37
timestamp 1676037725
transform 1 0 4508 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_3
timestamp 1676037725
transform 1 0 1380 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_15
timestamp 1676037725
transform 1 0 2484 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_27
timestamp 1676037725
transform 1 0 3588 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_31_35
timestamp 1676037725
transform 1 0 4324 0 -1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_32_3
timestamp 1676037725
transform 1 0 1380 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_15
timestamp 1676037725
transform 1 0 2484 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_27
timestamp 1676037725
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_29
timestamp 1676037725
transform 1 0 3772 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_37
timestamp 1676037725
transform 1 0 4508 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_3
timestamp 1676037725
transform 1 0 1380 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_15
timestamp 1676037725
transform 1 0 2484 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_27
timestamp 1676037725
transform 1 0 3588 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_33_35
timestamp 1676037725
transform 1 0 4324 0 -1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_34_3
timestamp 1676037725
transform 1 0 1380 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_15
timestamp 1676037725
transform 1 0 2484 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_27
timestamp 1676037725
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_34_29
timestamp 1676037725
transform 1 0 3772 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_37
timestamp 1676037725
transform 1 0 4508 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_3
timestamp 1676037725
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_15
timestamp 1676037725
transform 1 0 2484 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_27
timestamp 1676037725
transform 1 0 3588 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_35_35
timestamp 1676037725
transform 1 0 4324 0 -1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_36_3
timestamp 1676037725
transform 1 0 1380 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_15
timestamp 1676037725
transform 1 0 2484 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_27
timestamp 1676037725
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_29
timestamp 1676037725
transform 1 0 3772 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_37
timestamp 1676037725
transform 1 0 4508 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_3
timestamp 1676037725
transform 1 0 1380 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_15
timestamp 1676037725
transform 1 0 2484 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_27
timestamp 1676037725
transform 1 0 3588 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_37_35
timestamp 1676037725
transform 1 0 4324 0 -1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_38_3
timestamp 1676037725
transform 1 0 1380 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_15
timestamp 1676037725
transform 1 0 2484 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_27
timestamp 1676037725
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_38_29
timestamp 1676037725
transform 1 0 3772 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_38_37
timestamp 1676037725
transform 1 0 4508 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_3
timestamp 1676037725
transform 1 0 1380 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_15
timestamp 1676037725
transform 1 0 2484 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_39_27
timestamp 1676037725
transform 1 0 3588 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_39_29
timestamp 1676037725
transform 1 0 3772 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_37
timestamp 1676037725
transform 1 0 4508 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1676037725
transform 1 0 1104 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1676037725
transform -1 0 4876 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1676037725
transform 1 0 1104 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1676037725
transform -1 0 4876 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1676037725
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1676037725
transform -1 0 4876 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1676037725
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1676037725
transform -1 0 4876 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1676037725
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1676037725
transform -1 0 4876 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1676037725
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1676037725
transform -1 0 4876 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1676037725
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1676037725
transform -1 0 4876 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1676037725
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1676037725
transform -1 0 4876 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1676037725
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1676037725
transform -1 0 4876 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1676037725
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1676037725
transform -1 0 4876 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1676037725
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1676037725
transform -1 0 4876 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1676037725
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1676037725
transform -1 0 4876 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1676037725
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1676037725
transform -1 0 4876 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1676037725
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1676037725
transform -1 0 4876 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1676037725
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1676037725
transform -1 0 4876 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1676037725
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1676037725
transform -1 0 4876 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1676037725
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1676037725
transform -1 0 4876 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1676037725
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1676037725
transform -1 0 4876 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1676037725
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1676037725
transform -1 0 4876 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1676037725
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1676037725
transform -1 0 4876 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1676037725
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1676037725
transform -1 0 4876 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1676037725
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1676037725
transform -1 0 4876 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1676037725
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1676037725
transform -1 0 4876 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1676037725
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1676037725
transform -1 0 4876 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1676037725
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1676037725
transform -1 0 4876 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1676037725
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1676037725
transform -1 0 4876 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1676037725
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1676037725
transform -1 0 4876 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1676037725
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1676037725
transform -1 0 4876 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1676037725
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1676037725
transform -1 0 4876 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1676037725
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1676037725
transform -1 0 4876 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1676037725
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1676037725
transform -1 0 4876 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1676037725
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1676037725
transform -1 0 4876 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1676037725
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1676037725
transform -1 0 4876 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1676037725
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1676037725
transform -1 0 4876 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1676037725
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1676037725
transform -1 0 4876 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1676037725
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1676037725
transform -1 0 4876 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1676037725
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1676037725
transform -1 0 4876 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1676037725
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1676037725
transform -1 0 4876 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1676037725
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1676037725
transform -1 0 4876 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1676037725
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1676037725
transform -1 0 4876 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_80 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3680 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_81
timestamp 1676037725
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_82
timestamp 1676037725
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_83
timestamp 1676037725
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_84
timestamp 1676037725
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_85
timestamp 1676037725
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_86
timestamp 1676037725
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_87
timestamp 1676037725
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_88
timestamp 1676037725
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_89
timestamp 1676037725
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_90
timestamp 1676037725
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_91
timestamp 1676037725
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_92
timestamp 1676037725
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_93
timestamp 1676037725
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94
timestamp 1676037725
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1676037725
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 1676037725
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 1676037725
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 1676037725
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 1676037725
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 1676037725
transform 1 0 3680 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__clkinv_2  buf_clk_int pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 4324 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_4  buf_clk pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 1932 0 -1 2176
box -38 -48 682 592
use sky130_fd_sc_hd__dlxtp_1  latch\[0\] pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3312 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  latch\[1\]
timestamp 1676037725
transform 1 0 1840 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  latch\[2\]
timestamp 1676037725
transform 1 0 2392 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  latch\[3\]
timestamp 1676037725
transform 1 0 3312 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  latch\[4\]
timestamp 1676037725
transform 1 0 2392 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  latch\[5\]
timestamp 1676037725
transform 1 0 3312 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  latch\[6\]
timestamp 1676037725
transform 1 0 2392 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  latch\[7\]
timestamp 1676037725
transform 1 0 2392 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  out_flop_1 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3956 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_4  out_flop pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 2300 0 -1 6528
box -38 -48 2154 592
use sky130_fd_sc_hd__sdfxtp_1  scan_flop\[0\] pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 1564 0 1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__sdfxtp_1  scan_flop\[1\]
timestamp 1676037725
transform -1 0 4416 0 -1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__sdfxtp_1  scan_flop\[2\]
timestamp 1676037725
transform 1 0 1564 0 1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__sdfxtp_1  scan_flop\[3\]
timestamp 1676037725
transform -1 0 4416 0 -1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__sdfxtp_1  scan_flop\[4\]
timestamp 1676037725
transform -1 0 4416 0 -1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__sdfxtp_1  scan_flop\[5\]
timestamp 1676037725
transform 1 0 1564 0 1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__sdfxtp_1  scan_flop\[6\]
timestamp 1676037725
transform -1 0 4416 0 -1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__sdfxtp_1  scan_flop\[7\]
timestamp 1676037725
transform -1 0 4416 0 -1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__buf_4  through_buffers\[0\] pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 2944 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  through_buffers\[1\]
timestamp 1676037725
transform 1 0 3680 0 -1 2176
box -38 -48 590 592
<< labels >>
flabel metal2 s 386 0 442 800 0 FreeSans 224 90 0 0 clk_in
port 0 nsew signal input
flabel metal2 s 5538 0 5594 800 0 FreeSans 224 90 0 0 clk_out
port 1 nsew signal tristate
flabel metal2 s 1122 0 1178 800 0 FreeSans 224 90 0 0 data_in
port 2 nsew signal input
flabel metal2 s 4802 0 4858 800 0 FreeSans 224 90 0 0 data_out
port 3 nsew signal tristate
flabel metal2 s 2594 0 2650 800 0 FreeSans 224 90 0 0 latch_enable_in
port 4 nsew signal input
flabel metal2 s 3330 0 3386 800 0 FreeSans 224 90 0 0 latch_enable_out
port 5 nsew signal tristate
flabel metal3 s 5200 688 6000 808 0 FreeSans 480 0 0 0 module_data_in[0]
port 6 nsew signal tristate
flabel metal3 s 5200 2184 6000 2304 0 FreeSans 480 0 0 0 module_data_in[1]
port 7 nsew signal tristate
flabel metal3 s 5200 3680 6000 3800 0 FreeSans 480 0 0 0 module_data_in[2]
port 8 nsew signal tristate
flabel metal3 s 5200 5176 6000 5296 0 FreeSans 480 0 0 0 module_data_in[3]
port 9 nsew signal tristate
flabel metal3 s 5200 6672 6000 6792 0 FreeSans 480 0 0 0 module_data_in[4]
port 10 nsew signal tristate
flabel metal3 s 5200 8168 6000 8288 0 FreeSans 480 0 0 0 module_data_in[5]
port 11 nsew signal tristate
flabel metal3 s 5200 9664 6000 9784 0 FreeSans 480 0 0 0 module_data_in[6]
port 12 nsew signal tristate
flabel metal3 s 5200 11160 6000 11280 0 FreeSans 480 0 0 0 module_data_in[7]
port 13 nsew signal tristate
flabel metal3 s 5200 12656 6000 12776 0 FreeSans 480 0 0 0 module_data_out[0]
port 14 nsew signal input
flabel metal3 s 5200 14152 6000 14272 0 FreeSans 480 0 0 0 module_data_out[1]
port 15 nsew signal input
flabel metal3 s 5200 15648 6000 15768 0 FreeSans 480 0 0 0 module_data_out[2]
port 16 nsew signal input
flabel metal3 s 5200 17144 6000 17264 0 FreeSans 480 0 0 0 module_data_out[3]
port 17 nsew signal input
flabel metal3 s 5200 18640 6000 18760 0 FreeSans 480 0 0 0 module_data_out[4]
port 18 nsew signal input
flabel metal3 s 5200 20136 6000 20256 0 FreeSans 480 0 0 0 module_data_out[5]
port 19 nsew signal input
flabel metal3 s 5200 21632 6000 21752 0 FreeSans 480 0 0 0 module_data_out[6]
port 20 nsew signal input
flabel metal3 s 5200 23128 6000 23248 0 FreeSans 480 0 0 0 module_data_out[7]
port 21 nsew signal input
flabel metal2 s 1858 0 1914 800 0 FreeSans 224 90 0 0 scan_select_in
port 22 nsew signal input
flabel metal2 s 4066 0 4122 800 0 FreeSans 224 90 0 0 scan_select_out
port 23 nsew signal tristate
flabel metal4 s 1415 1040 1735 22896 0 FreeSans 1920 90 0 0 vccd1
port 24 nsew power bidirectional
flabel metal4 s 2358 1040 2678 22896 0 FreeSans 1920 90 0 0 vccd1
port 24 nsew power bidirectional
flabel metal4 s 3301 1040 3621 22896 0 FreeSans 1920 90 0 0 vccd1
port 24 nsew power bidirectional
flabel metal4 s 4244 1040 4564 22896 0 FreeSans 1920 90 0 0 vccd1
port 24 nsew power bidirectional
flabel metal4 s 1886 1040 2206 22896 0 FreeSans 1920 90 0 0 vssd1
port 25 nsew ground bidirectional
flabel metal4 s 2829 1040 3149 22896 0 FreeSans 1920 90 0 0 vssd1
port 25 nsew ground bidirectional
flabel metal4 s 3772 1040 4092 22896 0 FreeSans 1920 90 0 0 vssd1
port 25 nsew ground bidirectional
flabel metal4 s 4715 1040 5035 22896 0 FreeSans 1920 90 0 0 vssd1
port 25 nsew ground bidirectional
rlabel metal1 2990 22304 2990 22304 0 vccd1
rlabel via1 3069 22848 3069 22848 0 vssd1
rlabel metal1 4232 4794 4232 4794 0 clk
rlabel metal2 414 1350 414 1350 0 clk_in
rlabel metal1 4048 2006 4048 2006 0 clk_out
rlabel metal1 1979 7904 1979 7904 0 data_in
rlabel metal2 4830 823 4830 823 0 data_out
rlabel metal1 2806 1326 2806 1326 0 latch_enable_in
rlabel metal2 3358 1010 3358 1010 0 latch_enable_out
rlabel metal1 4738 2822 4738 2822 0 module_data_in[0]
rlabel metal1 2806 4998 2806 4998 0 module_data_in[1]
rlabel metal1 4324 4454 4324 4454 0 module_data_in[2]
rlabel metal1 4738 4250 4738 4250 0 module_data_in[3]
rlabel metal1 3588 5882 3588 5882 0 module_data_in[4]
rlabel metal1 4784 5338 4784 5338 0 module_data_in[5]
rlabel metal1 4324 6970 4324 6970 0 module_data_in[6]
rlabel via2 3450 11237 3450 11237 0 module_data_in[7]
rlabel metal1 3910 7922 3910 7922 0 module_data_out[0]
rlabel metal1 4508 7378 4508 7378 0 module_data_out[1]
rlabel metal3 4209 15572 4209 15572 0 module_data_out[2]
rlabel metal3 5160 17204 5160 17204 0 module_data_out[3]
rlabel metal3 4930 18700 4930 18700 0 module_data_out[4]
rlabel metal3 5313 19924 5313 19924 0 module_data_out[5]
rlabel metal1 4416 10642 4416 10642 0 module_data_out[6]
rlabel metal2 5198 23188 5198 23188 0 module_data_out[7]
rlabel metal1 3864 6630 3864 6630 0 net1
rlabel metal1 3680 3026 3680 3026 0 scan_data_in\[1\]
rlabel metal1 2208 5202 2208 5202 0 scan_data_in\[2\]
rlabel metal1 4646 4658 4646 4658 0 scan_data_in\[3\]
rlabel metal1 4554 4114 4554 4114 0 scan_data_in\[4\]
rlabel metal1 1932 8262 1932 8262 0 scan_data_in\[5\]
rlabel metal1 3450 5202 3450 5202 0 scan_data_in\[6\]
rlabel metal1 2852 10438 2852 10438 0 scan_data_in\[7\]
rlabel metal1 2622 9350 2622 9350 0 scan_data_out\[7\]
rlabel metal1 3726 1904 3726 1904 0 scan_select_in
rlabel metal2 4094 823 4094 823 0 scan_select_out
<< properties >>
string FIXED_BBOX 0 0 6000 24000
<< end >>
