module MichaelBell_6bit_fifo (vccd1,
    vssd1,
    io_in,
    io_out);
 input vccd1;
 input vssd1;
 input [7:0] io_in;
 output [7:0] io_out;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire _203_;
 wire _204_;
 wire _205_;
 wire _206_;
 wire _207_;
 wire _208_;
 wire _209_;
 wire _210_;
 wire _211_;
 wire _212_;
 wire _213_;
 wire _214_;
 wire _215_;
 wire _216_;
 wire _217_;
 wire _218_;
 wire _219_;
 wire _220_;
 wire _221_;
 wire _222_;
 wire _223_;
 wire _224_;
 wire _225_;
 wire _226_;
 wire _227_;
 wire _228_;
 wire _229_;
 wire _230_;
 wire _231_;
 wire _232_;
 wire _233_;
 wire _234_;
 wire _235_;
 wire _236_;
 wire _237_;
 wire _238_;
 wire _239_;
 wire _240_;
 wire _241_;
 wire _242_;
 wire _243_;
 wire _244_;
 wire _245_;
 wire _246_;
 wire _247_;
 wire _248_;
 wire _249_;
 wire _250_;
 wire _251_;
 wire \data_in_buffer[0].A ;
 wire \data_in_buffer[0].X ;
 wire \data_in_buffer[0].b[0] ;
 wire \data_in_buffer[0].genblk1[0].mid ;
 wire \data_in_buffer[0].genblk1[1].mid ;
 wire \data_in_buffer[1].A ;
 wire \data_in_buffer[1].X ;
 wire \data_in_buffer[1].b[0] ;
 wire \data_in_buffer[1].genblk1[0].mid ;
 wire \data_in_buffer[1].genblk1[1].mid ;
 wire \data_in_buffer[2].A ;
 wire \data_in_buffer[2].X ;
 wire \data_in_buffer[2].b[0] ;
 wire \data_in_buffer[2].genblk1[0].mid ;
 wire \data_in_buffer[2].genblk1[1].mid ;
 wire \data_in_buffer[3].A ;
 wire \data_in_buffer[3].X ;
 wire \data_in_buffer[3].b[0] ;
 wire \data_in_buffer[3].genblk1[0].mid ;
 wire \data_in_buffer[3].genblk1[1].mid ;
 wire \data_in_buffer[4].A ;
 wire \data_in_buffer[4].X ;
 wire \data_in_buffer[4].b[0] ;
 wire \data_in_buffer[4].genblk1[0].mid ;
 wire \data_in_buffer[4].genblk1[1].mid ;
 wire \data_in_buffer[5].A ;
 wire \data_in_buffer[5].X ;
 wire \data_in_buffer[5].b[0] ;
 wire \data_in_buffer[5].genblk1[0].mid ;
 wire \data_in_buffer[5].genblk1[1].mid ;
 wire \f_fifo.data_in[0] ;
 wire \f_fifo.data_in[1] ;
 wire \f_fifo.data_in[2] ;
 wire \f_fifo.data_in[3] ;
 wire \f_fifo.data_in[4] ;
 wire \f_fifo.data_in[5] ;
 wire \f_fifo.empty_n ;
 wire \f_fifo.fifo_data[0][0] ;
 wire \f_fifo.fifo_data[0][1] ;
 wire \f_fifo.fifo_data[0][2] ;
 wire \f_fifo.fifo_data[0][3] ;
 wire \f_fifo.fifo_data[0][4] ;
 wire \f_fifo.fifo_data[0][5] ;
 wire \f_fifo.fifo_data[1][0] ;
 wire \f_fifo.fifo_data[1][1] ;
 wire \f_fifo.fifo_data[1][2] ;
 wire \f_fifo.fifo_data[1][3] ;
 wire \f_fifo.fifo_data[1][4] ;
 wire \f_fifo.fifo_data[1][5] ;
 wire \f_fifo.fifo_data[2][0] ;
 wire \f_fifo.fifo_data[2][1] ;
 wire \f_fifo.fifo_data[2][2] ;
 wire \f_fifo.fifo_data[2][3] ;
 wire \f_fifo.fifo_data[2][4] ;
 wire \f_fifo.fifo_data[2][5] ;
 wire \f_fifo.fifo_data[3][0] ;
 wire \f_fifo.fifo_data[3][1] ;
 wire \f_fifo.fifo_data[3][2] ;
 wire \f_fifo.fifo_data[3][3] ;
 wire \f_fifo.fifo_data[3][4] ;
 wire \f_fifo.fifo_data[3][5] ;
 wire \f_fifo.read_addr[0] ;
 wire \f_fifo.read_addr[1] ;
 wire \f_fifo.reset_n ;
 wire \f_fifo.write_addr[0] ;
 wire \f_fifo.write_addr[1] ;
 wire \l_fifo.genblk1[0].entry.empty ;
 wire \l_fifo.genblk1[0].entry.input_buf[0].A ;
 wire \l_fifo.genblk1[0].entry.input_buf[0].X ;
 wire \l_fifo.genblk1[0].entry.input_buf[0].genblk1[0].mid ;
 wire \l_fifo.genblk1[0].entry.input_buf[1].A ;
 wire \l_fifo.genblk1[0].entry.input_buf[1].X ;
 wire \l_fifo.genblk1[0].entry.input_buf[1].genblk1[0].mid ;
 wire \l_fifo.genblk1[0].entry.input_buf[2].A ;
 wire \l_fifo.genblk1[0].entry.input_buf[2].X ;
 wire \l_fifo.genblk1[0].entry.input_buf[2].genblk1[0].mid ;
 wire \l_fifo.genblk1[0].entry.input_buf[3].A ;
 wire \l_fifo.genblk1[0].entry.input_buf[3].X ;
 wire \l_fifo.genblk1[0].entry.input_buf[3].genblk1[0].mid ;
 wire \l_fifo.genblk1[0].entry.input_buf[4].A ;
 wire \l_fifo.genblk1[0].entry.input_buf[4].X ;
 wire \l_fifo.genblk1[0].entry.input_buf[4].genblk1[0].mid ;
 wire \l_fifo.genblk1[0].entry.input_buf[5].A ;
 wire \l_fifo.genblk1[0].entry.input_buf[5].X ;
 wire \l_fifo.genblk1[0].entry.input_buf[5].genblk1[0].mid ;
 wire \l_fifo.genblk1[10].entry.empty ;
 wire \l_fifo.genblk1[10].entry.input_buf[0].A ;
 wire \l_fifo.genblk1[10].entry.input_buf[0].X ;
 wire \l_fifo.genblk1[10].entry.input_buf[0].genblk1[0].mid ;
 wire \l_fifo.genblk1[10].entry.input_buf[1].A ;
 wire \l_fifo.genblk1[10].entry.input_buf[1].X ;
 wire \l_fifo.genblk1[10].entry.input_buf[1].genblk1[0].mid ;
 wire \l_fifo.genblk1[10].entry.input_buf[2].A ;
 wire \l_fifo.genblk1[10].entry.input_buf[2].X ;
 wire \l_fifo.genblk1[10].entry.input_buf[2].genblk1[0].mid ;
 wire \l_fifo.genblk1[10].entry.input_buf[3].A ;
 wire \l_fifo.genblk1[10].entry.input_buf[3].X ;
 wire \l_fifo.genblk1[10].entry.input_buf[3].genblk1[0].mid ;
 wire \l_fifo.genblk1[10].entry.input_buf[4].A ;
 wire \l_fifo.genblk1[10].entry.input_buf[4].X ;
 wire \l_fifo.genblk1[10].entry.input_buf[4].genblk1[0].mid ;
 wire \l_fifo.genblk1[10].entry.input_buf[5].A ;
 wire \l_fifo.genblk1[10].entry.input_buf[5].X ;
 wire \l_fifo.genblk1[10].entry.input_buf[5].genblk1[0].mid ;
 wire \l_fifo.genblk1[10].entry.next_is_empty ;
 wire \l_fifo.genblk1[11].entry.empty ;
 wire \l_fifo.genblk1[11].entry.input_buf[0].A ;
 wire \l_fifo.genblk1[11].entry.input_buf[0].X ;
 wire \l_fifo.genblk1[11].entry.input_buf[0].genblk1[0].mid ;
 wire \l_fifo.genblk1[11].entry.input_buf[1].A ;
 wire \l_fifo.genblk1[11].entry.input_buf[1].X ;
 wire \l_fifo.genblk1[11].entry.input_buf[1].genblk1[0].mid ;
 wire \l_fifo.genblk1[11].entry.input_buf[2].A ;
 wire \l_fifo.genblk1[11].entry.input_buf[2].X ;
 wire \l_fifo.genblk1[11].entry.input_buf[2].genblk1[0].mid ;
 wire \l_fifo.genblk1[11].entry.input_buf[3].A ;
 wire \l_fifo.genblk1[11].entry.input_buf[3].X ;
 wire \l_fifo.genblk1[11].entry.input_buf[3].genblk1[0].mid ;
 wire \l_fifo.genblk1[11].entry.input_buf[4].A ;
 wire \l_fifo.genblk1[11].entry.input_buf[4].X ;
 wire \l_fifo.genblk1[11].entry.input_buf[4].genblk1[0].mid ;
 wire \l_fifo.genblk1[11].entry.input_buf[5].A ;
 wire \l_fifo.genblk1[11].entry.input_buf[5].X ;
 wire \l_fifo.genblk1[11].entry.input_buf[5].genblk1[0].mid ;
 wire \l_fifo.genblk1[12].entry.empty ;
 wire \l_fifo.genblk1[12].entry.input_buf[0].A ;
 wire \l_fifo.genblk1[12].entry.input_buf[0].X ;
 wire \l_fifo.genblk1[12].entry.input_buf[0].genblk1[0].mid ;
 wire \l_fifo.genblk1[12].entry.input_buf[1].A ;
 wire \l_fifo.genblk1[12].entry.input_buf[1].X ;
 wire \l_fifo.genblk1[12].entry.input_buf[1].genblk1[0].mid ;
 wire \l_fifo.genblk1[12].entry.input_buf[2].A ;
 wire \l_fifo.genblk1[12].entry.input_buf[2].X ;
 wire \l_fifo.genblk1[12].entry.input_buf[2].genblk1[0].mid ;
 wire \l_fifo.genblk1[12].entry.input_buf[3].A ;
 wire \l_fifo.genblk1[12].entry.input_buf[3].X ;
 wire \l_fifo.genblk1[12].entry.input_buf[3].genblk1[0].mid ;
 wire \l_fifo.genblk1[12].entry.input_buf[4].A ;
 wire \l_fifo.genblk1[12].entry.input_buf[4].X ;
 wire \l_fifo.genblk1[12].entry.input_buf[4].genblk1[0].mid ;
 wire \l_fifo.genblk1[12].entry.input_buf[5].A ;
 wire \l_fifo.genblk1[12].entry.input_buf[5].X ;
 wire \l_fifo.genblk1[12].entry.input_buf[5].genblk1[0].mid ;
 wire \l_fifo.genblk1[13].entry.empty ;
 wire \l_fifo.genblk1[13].entry.input_buf[0].A ;
 wire \l_fifo.genblk1[13].entry.input_buf[0].X ;
 wire \l_fifo.genblk1[13].entry.input_buf[0].genblk1[0].mid ;
 wire \l_fifo.genblk1[13].entry.input_buf[1].A ;
 wire \l_fifo.genblk1[13].entry.input_buf[1].X ;
 wire \l_fifo.genblk1[13].entry.input_buf[1].genblk1[0].mid ;
 wire \l_fifo.genblk1[13].entry.input_buf[2].A ;
 wire \l_fifo.genblk1[13].entry.input_buf[2].X ;
 wire \l_fifo.genblk1[13].entry.input_buf[2].genblk1[0].mid ;
 wire \l_fifo.genblk1[13].entry.input_buf[3].A ;
 wire \l_fifo.genblk1[13].entry.input_buf[3].X ;
 wire \l_fifo.genblk1[13].entry.input_buf[3].genblk1[0].mid ;
 wire \l_fifo.genblk1[13].entry.input_buf[4].A ;
 wire \l_fifo.genblk1[13].entry.input_buf[4].X ;
 wire \l_fifo.genblk1[13].entry.input_buf[4].genblk1[0].mid ;
 wire \l_fifo.genblk1[13].entry.input_buf[5].A ;
 wire \l_fifo.genblk1[13].entry.input_buf[5].X ;
 wire \l_fifo.genblk1[13].entry.input_buf[5].genblk1[0].mid ;
 wire \l_fifo.genblk1[14].entry.empty ;
 wire \l_fifo.genblk1[14].entry.input_buf[0].A ;
 wire \l_fifo.genblk1[14].entry.input_buf[0].X ;
 wire \l_fifo.genblk1[14].entry.input_buf[0].genblk1[0].mid ;
 wire \l_fifo.genblk1[14].entry.input_buf[1].A ;
 wire \l_fifo.genblk1[14].entry.input_buf[1].X ;
 wire \l_fifo.genblk1[14].entry.input_buf[1].genblk1[0].mid ;
 wire \l_fifo.genblk1[14].entry.input_buf[2].A ;
 wire \l_fifo.genblk1[14].entry.input_buf[2].X ;
 wire \l_fifo.genblk1[14].entry.input_buf[2].genblk1[0].mid ;
 wire \l_fifo.genblk1[14].entry.input_buf[3].A ;
 wire \l_fifo.genblk1[14].entry.input_buf[3].X ;
 wire \l_fifo.genblk1[14].entry.input_buf[3].genblk1[0].mid ;
 wire \l_fifo.genblk1[14].entry.input_buf[4].A ;
 wire \l_fifo.genblk1[14].entry.input_buf[4].X ;
 wire \l_fifo.genblk1[14].entry.input_buf[4].genblk1[0].mid ;
 wire \l_fifo.genblk1[14].entry.input_buf[5].A ;
 wire \l_fifo.genblk1[14].entry.input_buf[5].X ;
 wire \l_fifo.genblk1[14].entry.input_buf[5].genblk1[0].mid ;
 wire \l_fifo.genblk1[15].entry.empty ;
 wire \l_fifo.genblk1[15].entry.input_buf[0].A ;
 wire \l_fifo.genblk1[15].entry.input_buf[0].X ;
 wire \l_fifo.genblk1[15].entry.input_buf[0].genblk1[0].mid ;
 wire \l_fifo.genblk1[15].entry.input_buf[1].A ;
 wire \l_fifo.genblk1[15].entry.input_buf[1].X ;
 wire \l_fifo.genblk1[15].entry.input_buf[1].genblk1[0].mid ;
 wire \l_fifo.genblk1[15].entry.input_buf[2].A ;
 wire \l_fifo.genblk1[15].entry.input_buf[2].X ;
 wire \l_fifo.genblk1[15].entry.input_buf[2].genblk1[0].mid ;
 wire \l_fifo.genblk1[15].entry.input_buf[3].A ;
 wire \l_fifo.genblk1[15].entry.input_buf[3].X ;
 wire \l_fifo.genblk1[15].entry.input_buf[3].genblk1[0].mid ;
 wire \l_fifo.genblk1[15].entry.input_buf[4].A ;
 wire \l_fifo.genblk1[15].entry.input_buf[4].X ;
 wire \l_fifo.genblk1[15].entry.input_buf[4].genblk1[0].mid ;
 wire \l_fifo.genblk1[15].entry.input_buf[5].A ;
 wire \l_fifo.genblk1[15].entry.input_buf[5].X ;
 wire \l_fifo.genblk1[15].entry.input_buf[5].genblk1[0].mid ;
 wire \l_fifo.genblk1[16].entry.empty ;
 wire \l_fifo.genblk1[16].entry.input_buf[0].A ;
 wire \l_fifo.genblk1[16].entry.input_buf[0].X ;
 wire \l_fifo.genblk1[16].entry.input_buf[0].genblk1[0].mid ;
 wire \l_fifo.genblk1[16].entry.input_buf[1].A ;
 wire \l_fifo.genblk1[16].entry.input_buf[1].X ;
 wire \l_fifo.genblk1[16].entry.input_buf[1].genblk1[0].mid ;
 wire \l_fifo.genblk1[16].entry.input_buf[2].A ;
 wire \l_fifo.genblk1[16].entry.input_buf[2].X ;
 wire \l_fifo.genblk1[16].entry.input_buf[2].genblk1[0].mid ;
 wire \l_fifo.genblk1[16].entry.input_buf[3].A ;
 wire \l_fifo.genblk1[16].entry.input_buf[3].X ;
 wire \l_fifo.genblk1[16].entry.input_buf[3].genblk1[0].mid ;
 wire \l_fifo.genblk1[16].entry.input_buf[4].A ;
 wire \l_fifo.genblk1[16].entry.input_buf[4].X ;
 wire \l_fifo.genblk1[16].entry.input_buf[4].genblk1[0].mid ;
 wire \l_fifo.genblk1[16].entry.input_buf[5].A ;
 wire \l_fifo.genblk1[16].entry.input_buf[5].X ;
 wire \l_fifo.genblk1[16].entry.input_buf[5].genblk1[0].mid ;
 wire \l_fifo.genblk1[17].entry.empty ;
 wire \l_fifo.genblk1[17].entry.input_buf[0].A ;
 wire \l_fifo.genblk1[17].entry.input_buf[0].X ;
 wire \l_fifo.genblk1[17].entry.input_buf[0].genblk1[0].mid ;
 wire \l_fifo.genblk1[17].entry.input_buf[1].A ;
 wire \l_fifo.genblk1[17].entry.input_buf[1].X ;
 wire \l_fifo.genblk1[17].entry.input_buf[1].genblk1[0].mid ;
 wire \l_fifo.genblk1[17].entry.input_buf[2].A ;
 wire \l_fifo.genblk1[17].entry.input_buf[2].X ;
 wire \l_fifo.genblk1[17].entry.input_buf[2].genblk1[0].mid ;
 wire \l_fifo.genblk1[17].entry.input_buf[3].A ;
 wire \l_fifo.genblk1[17].entry.input_buf[3].X ;
 wire \l_fifo.genblk1[17].entry.input_buf[3].genblk1[0].mid ;
 wire \l_fifo.genblk1[17].entry.input_buf[4].A ;
 wire \l_fifo.genblk1[17].entry.input_buf[4].X ;
 wire \l_fifo.genblk1[17].entry.input_buf[4].genblk1[0].mid ;
 wire \l_fifo.genblk1[17].entry.input_buf[5].A ;
 wire \l_fifo.genblk1[17].entry.input_buf[5].X ;
 wire \l_fifo.genblk1[17].entry.input_buf[5].genblk1[0].mid ;
 wire \l_fifo.genblk1[18].entry.empty ;
 wire \l_fifo.genblk1[18].entry.input_buf[0].A ;
 wire \l_fifo.genblk1[18].entry.input_buf[0].X ;
 wire \l_fifo.genblk1[18].entry.input_buf[0].genblk1[0].mid ;
 wire \l_fifo.genblk1[18].entry.input_buf[1].A ;
 wire \l_fifo.genblk1[18].entry.input_buf[1].X ;
 wire \l_fifo.genblk1[18].entry.input_buf[1].genblk1[0].mid ;
 wire \l_fifo.genblk1[18].entry.input_buf[2].A ;
 wire \l_fifo.genblk1[18].entry.input_buf[2].X ;
 wire \l_fifo.genblk1[18].entry.input_buf[2].genblk1[0].mid ;
 wire \l_fifo.genblk1[18].entry.input_buf[3].A ;
 wire \l_fifo.genblk1[18].entry.input_buf[3].X ;
 wire \l_fifo.genblk1[18].entry.input_buf[3].genblk1[0].mid ;
 wire \l_fifo.genblk1[18].entry.input_buf[4].A ;
 wire \l_fifo.genblk1[18].entry.input_buf[4].X ;
 wire \l_fifo.genblk1[18].entry.input_buf[4].genblk1[0].mid ;
 wire \l_fifo.genblk1[18].entry.input_buf[5].A ;
 wire \l_fifo.genblk1[18].entry.input_buf[5].X ;
 wire \l_fifo.genblk1[18].entry.input_buf[5].genblk1[0].mid ;
 wire \l_fifo.genblk1[19].entry.empty ;
 wire \l_fifo.genblk1[19].entry.input_buf[0].A ;
 wire \l_fifo.genblk1[19].entry.input_buf[0].X ;
 wire \l_fifo.genblk1[19].entry.input_buf[0].genblk1[0].mid ;
 wire \l_fifo.genblk1[19].entry.input_buf[1].A ;
 wire \l_fifo.genblk1[19].entry.input_buf[1].X ;
 wire \l_fifo.genblk1[19].entry.input_buf[1].genblk1[0].mid ;
 wire \l_fifo.genblk1[19].entry.input_buf[2].A ;
 wire \l_fifo.genblk1[19].entry.input_buf[2].X ;
 wire \l_fifo.genblk1[19].entry.input_buf[2].genblk1[0].mid ;
 wire \l_fifo.genblk1[19].entry.input_buf[3].A ;
 wire \l_fifo.genblk1[19].entry.input_buf[3].X ;
 wire \l_fifo.genblk1[19].entry.input_buf[3].genblk1[0].mid ;
 wire \l_fifo.genblk1[19].entry.input_buf[4].A ;
 wire \l_fifo.genblk1[19].entry.input_buf[4].X ;
 wire \l_fifo.genblk1[19].entry.input_buf[4].genblk1[0].mid ;
 wire \l_fifo.genblk1[19].entry.input_buf[5].A ;
 wire \l_fifo.genblk1[19].entry.input_buf[5].X ;
 wire \l_fifo.genblk1[19].entry.input_buf[5].genblk1[0].mid ;
 wire \l_fifo.genblk1[1].entry.empty ;
 wire \l_fifo.genblk1[1].entry.input_buf[0].A ;
 wire \l_fifo.genblk1[1].entry.input_buf[0].X ;
 wire \l_fifo.genblk1[1].entry.input_buf[0].genblk1[0].mid ;
 wire \l_fifo.genblk1[1].entry.input_buf[1].A ;
 wire \l_fifo.genblk1[1].entry.input_buf[1].X ;
 wire \l_fifo.genblk1[1].entry.input_buf[1].genblk1[0].mid ;
 wire \l_fifo.genblk1[1].entry.input_buf[2].A ;
 wire \l_fifo.genblk1[1].entry.input_buf[2].X ;
 wire \l_fifo.genblk1[1].entry.input_buf[2].genblk1[0].mid ;
 wire \l_fifo.genblk1[1].entry.input_buf[3].A ;
 wire \l_fifo.genblk1[1].entry.input_buf[3].X ;
 wire \l_fifo.genblk1[1].entry.input_buf[3].genblk1[0].mid ;
 wire \l_fifo.genblk1[1].entry.input_buf[4].A ;
 wire \l_fifo.genblk1[1].entry.input_buf[4].X ;
 wire \l_fifo.genblk1[1].entry.input_buf[4].genblk1[0].mid ;
 wire \l_fifo.genblk1[1].entry.input_buf[5].A ;
 wire \l_fifo.genblk1[1].entry.input_buf[5].X ;
 wire \l_fifo.genblk1[1].entry.input_buf[5].genblk1[0].mid ;
 wire \l_fifo.genblk1[20].entry.empty ;
 wire \l_fifo.genblk1[20].entry.input_buf[0].A ;
 wire \l_fifo.genblk1[20].entry.input_buf[0].X ;
 wire \l_fifo.genblk1[20].entry.input_buf[0].genblk1[0].mid ;
 wire \l_fifo.genblk1[20].entry.input_buf[1].A ;
 wire \l_fifo.genblk1[20].entry.input_buf[1].X ;
 wire \l_fifo.genblk1[20].entry.input_buf[1].genblk1[0].mid ;
 wire \l_fifo.genblk1[20].entry.input_buf[2].A ;
 wire \l_fifo.genblk1[20].entry.input_buf[2].X ;
 wire \l_fifo.genblk1[20].entry.input_buf[2].genblk1[0].mid ;
 wire \l_fifo.genblk1[20].entry.input_buf[3].A ;
 wire \l_fifo.genblk1[20].entry.input_buf[3].X ;
 wire \l_fifo.genblk1[20].entry.input_buf[3].genblk1[0].mid ;
 wire \l_fifo.genblk1[20].entry.input_buf[4].A ;
 wire \l_fifo.genblk1[20].entry.input_buf[4].X ;
 wire \l_fifo.genblk1[20].entry.input_buf[4].genblk1[0].mid ;
 wire \l_fifo.genblk1[20].entry.input_buf[5].A ;
 wire \l_fifo.genblk1[20].entry.input_buf[5].X ;
 wire \l_fifo.genblk1[20].entry.input_buf[5].genblk1[0].mid ;
 wire \l_fifo.genblk1[21].entry.empty ;
 wire \l_fifo.genblk1[21].entry.input_buf[0].A ;
 wire \l_fifo.genblk1[21].entry.input_buf[0].X ;
 wire \l_fifo.genblk1[21].entry.input_buf[0].genblk1[0].mid ;
 wire \l_fifo.genblk1[21].entry.input_buf[1].A ;
 wire \l_fifo.genblk1[21].entry.input_buf[1].X ;
 wire \l_fifo.genblk1[21].entry.input_buf[1].genblk1[0].mid ;
 wire \l_fifo.genblk1[21].entry.input_buf[2].A ;
 wire \l_fifo.genblk1[21].entry.input_buf[2].X ;
 wire \l_fifo.genblk1[21].entry.input_buf[2].genblk1[0].mid ;
 wire \l_fifo.genblk1[21].entry.input_buf[3].A ;
 wire \l_fifo.genblk1[21].entry.input_buf[3].X ;
 wire \l_fifo.genblk1[21].entry.input_buf[3].genblk1[0].mid ;
 wire \l_fifo.genblk1[21].entry.input_buf[4].A ;
 wire \l_fifo.genblk1[21].entry.input_buf[4].X ;
 wire \l_fifo.genblk1[21].entry.input_buf[4].genblk1[0].mid ;
 wire \l_fifo.genblk1[21].entry.input_buf[5].A ;
 wire \l_fifo.genblk1[21].entry.input_buf[5].X ;
 wire \l_fifo.genblk1[21].entry.input_buf[5].genblk1[0].mid ;
 wire \l_fifo.genblk1[22].entry.empty ;
 wire \l_fifo.genblk1[22].entry.input_buf[0].A ;
 wire \l_fifo.genblk1[22].entry.input_buf[0].X ;
 wire \l_fifo.genblk1[22].entry.input_buf[0].genblk1[0].mid ;
 wire \l_fifo.genblk1[22].entry.input_buf[1].A ;
 wire \l_fifo.genblk1[22].entry.input_buf[1].X ;
 wire \l_fifo.genblk1[22].entry.input_buf[1].genblk1[0].mid ;
 wire \l_fifo.genblk1[22].entry.input_buf[2].A ;
 wire \l_fifo.genblk1[22].entry.input_buf[2].X ;
 wire \l_fifo.genblk1[22].entry.input_buf[2].genblk1[0].mid ;
 wire \l_fifo.genblk1[22].entry.input_buf[3].A ;
 wire \l_fifo.genblk1[22].entry.input_buf[3].X ;
 wire \l_fifo.genblk1[22].entry.input_buf[3].genblk1[0].mid ;
 wire \l_fifo.genblk1[22].entry.input_buf[4].A ;
 wire \l_fifo.genblk1[22].entry.input_buf[4].X ;
 wire \l_fifo.genblk1[22].entry.input_buf[4].genblk1[0].mid ;
 wire \l_fifo.genblk1[22].entry.input_buf[5].A ;
 wire \l_fifo.genblk1[22].entry.input_buf[5].X ;
 wire \l_fifo.genblk1[22].entry.input_buf[5].genblk1[0].mid ;
 wire \l_fifo.genblk1[23].entry.empty ;
 wire \l_fifo.genblk1[23].entry.input_buf[0].A ;
 wire \l_fifo.genblk1[23].entry.input_buf[0].X ;
 wire \l_fifo.genblk1[23].entry.input_buf[0].genblk1[0].mid ;
 wire \l_fifo.genblk1[23].entry.input_buf[1].A ;
 wire \l_fifo.genblk1[23].entry.input_buf[1].X ;
 wire \l_fifo.genblk1[23].entry.input_buf[1].genblk1[0].mid ;
 wire \l_fifo.genblk1[23].entry.input_buf[2].A ;
 wire \l_fifo.genblk1[23].entry.input_buf[2].X ;
 wire \l_fifo.genblk1[23].entry.input_buf[2].genblk1[0].mid ;
 wire \l_fifo.genblk1[23].entry.input_buf[3].A ;
 wire \l_fifo.genblk1[23].entry.input_buf[3].X ;
 wire \l_fifo.genblk1[23].entry.input_buf[3].genblk1[0].mid ;
 wire \l_fifo.genblk1[23].entry.input_buf[4].A ;
 wire \l_fifo.genblk1[23].entry.input_buf[4].X ;
 wire \l_fifo.genblk1[23].entry.input_buf[4].genblk1[0].mid ;
 wire \l_fifo.genblk1[23].entry.input_buf[5].A ;
 wire \l_fifo.genblk1[23].entry.input_buf[5].X ;
 wire \l_fifo.genblk1[23].entry.input_buf[5].genblk1[0].mid ;
 wire \l_fifo.genblk1[24].entry.empty ;
 wire \l_fifo.genblk1[24].entry.input_buf[0].A ;
 wire \l_fifo.genblk1[24].entry.input_buf[0].X ;
 wire \l_fifo.genblk1[24].entry.input_buf[0].genblk1[0].mid ;
 wire \l_fifo.genblk1[24].entry.input_buf[1].A ;
 wire \l_fifo.genblk1[24].entry.input_buf[1].X ;
 wire \l_fifo.genblk1[24].entry.input_buf[1].genblk1[0].mid ;
 wire \l_fifo.genblk1[24].entry.input_buf[2].A ;
 wire \l_fifo.genblk1[24].entry.input_buf[2].X ;
 wire \l_fifo.genblk1[24].entry.input_buf[2].genblk1[0].mid ;
 wire \l_fifo.genblk1[24].entry.input_buf[3].A ;
 wire \l_fifo.genblk1[24].entry.input_buf[3].X ;
 wire \l_fifo.genblk1[24].entry.input_buf[3].genblk1[0].mid ;
 wire \l_fifo.genblk1[24].entry.input_buf[4].A ;
 wire \l_fifo.genblk1[24].entry.input_buf[4].X ;
 wire \l_fifo.genblk1[24].entry.input_buf[4].genblk1[0].mid ;
 wire \l_fifo.genblk1[24].entry.input_buf[5].A ;
 wire \l_fifo.genblk1[24].entry.input_buf[5].X ;
 wire \l_fifo.genblk1[24].entry.input_buf[5].genblk1[0].mid ;
 wire \l_fifo.genblk1[25].entry.empty ;
 wire \l_fifo.genblk1[25].entry.input_buf[0].A ;
 wire \l_fifo.genblk1[25].entry.input_buf[0].X ;
 wire \l_fifo.genblk1[25].entry.input_buf[0].genblk1[0].mid ;
 wire \l_fifo.genblk1[25].entry.input_buf[1].A ;
 wire \l_fifo.genblk1[25].entry.input_buf[1].X ;
 wire \l_fifo.genblk1[25].entry.input_buf[1].genblk1[0].mid ;
 wire \l_fifo.genblk1[25].entry.input_buf[2].A ;
 wire \l_fifo.genblk1[25].entry.input_buf[2].X ;
 wire \l_fifo.genblk1[25].entry.input_buf[2].genblk1[0].mid ;
 wire \l_fifo.genblk1[25].entry.input_buf[3].A ;
 wire \l_fifo.genblk1[25].entry.input_buf[3].X ;
 wire \l_fifo.genblk1[25].entry.input_buf[3].genblk1[0].mid ;
 wire \l_fifo.genblk1[25].entry.input_buf[4].A ;
 wire \l_fifo.genblk1[25].entry.input_buf[4].X ;
 wire \l_fifo.genblk1[25].entry.input_buf[4].genblk1[0].mid ;
 wire \l_fifo.genblk1[25].entry.input_buf[5].A ;
 wire \l_fifo.genblk1[25].entry.input_buf[5].X ;
 wire \l_fifo.genblk1[25].entry.input_buf[5].genblk1[0].mid ;
 wire \l_fifo.genblk1[26].entry.empty ;
 wire \l_fifo.genblk1[26].entry.input_buf[0].A ;
 wire \l_fifo.genblk1[26].entry.input_buf[0].X ;
 wire \l_fifo.genblk1[26].entry.input_buf[0].genblk1[0].mid ;
 wire \l_fifo.genblk1[26].entry.input_buf[1].A ;
 wire \l_fifo.genblk1[26].entry.input_buf[1].X ;
 wire \l_fifo.genblk1[26].entry.input_buf[1].genblk1[0].mid ;
 wire \l_fifo.genblk1[26].entry.input_buf[2].A ;
 wire \l_fifo.genblk1[26].entry.input_buf[2].X ;
 wire \l_fifo.genblk1[26].entry.input_buf[2].genblk1[0].mid ;
 wire \l_fifo.genblk1[26].entry.input_buf[3].A ;
 wire \l_fifo.genblk1[26].entry.input_buf[3].X ;
 wire \l_fifo.genblk1[26].entry.input_buf[3].genblk1[0].mid ;
 wire \l_fifo.genblk1[26].entry.input_buf[4].A ;
 wire \l_fifo.genblk1[26].entry.input_buf[4].X ;
 wire \l_fifo.genblk1[26].entry.input_buf[4].genblk1[0].mid ;
 wire \l_fifo.genblk1[26].entry.input_buf[5].A ;
 wire \l_fifo.genblk1[26].entry.input_buf[5].X ;
 wire \l_fifo.genblk1[26].entry.input_buf[5].genblk1[0].mid ;
 wire \l_fifo.genblk1[27].entry.empty ;
 wire \l_fifo.genblk1[27].entry.input_buf[0].A ;
 wire \l_fifo.genblk1[27].entry.input_buf[0].X ;
 wire \l_fifo.genblk1[27].entry.input_buf[0].genblk1[0].mid ;
 wire \l_fifo.genblk1[27].entry.input_buf[1].A ;
 wire \l_fifo.genblk1[27].entry.input_buf[1].X ;
 wire \l_fifo.genblk1[27].entry.input_buf[1].genblk1[0].mid ;
 wire \l_fifo.genblk1[27].entry.input_buf[2].A ;
 wire \l_fifo.genblk1[27].entry.input_buf[2].X ;
 wire \l_fifo.genblk1[27].entry.input_buf[2].genblk1[0].mid ;
 wire \l_fifo.genblk1[27].entry.input_buf[3].A ;
 wire \l_fifo.genblk1[27].entry.input_buf[3].X ;
 wire \l_fifo.genblk1[27].entry.input_buf[3].genblk1[0].mid ;
 wire \l_fifo.genblk1[27].entry.input_buf[4].A ;
 wire \l_fifo.genblk1[27].entry.input_buf[4].X ;
 wire \l_fifo.genblk1[27].entry.input_buf[4].genblk1[0].mid ;
 wire \l_fifo.genblk1[27].entry.input_buf[5].A ;
 wire \l_fifo.genblk1[27].entry.input_buf[5].X ;
 wire \l_fifo.genblk1[27].entry.input_buf[5].genblk1[0].mid ;
 wire \l_fifo.genblk1[28].entry.empty ;
 wire \l_fifo.genblk1[28].entry.input_buf[0].A ;
 wire \l_fifo.genblk1[28].entry.input_buf[0].X ;
 wire \l_fifo.genblk1[28].entry.input_buf[0].genblk1[0].mid ;
 wire \l_fifo.genblk1[28].entry.input_buf[1].A ;
 wire \l_fifo.genblk1[28].entry.input_buf[1].X ;
 wire \l_fifo.genblk1[28].entry.input_buf[1].genblk1[0].mid ;
 wire \l_fifo.genblk1[28].entry.input_buf[2].A ;
 wire \l_fifo.genblk1[28].entry.input_buf[2].X ;
 wire \l_fifo.genblk1[28].entry.input_buf[2].genblk1[0].mid ;
 wire \l_fifo.genblk1[28].entry.input_buf[3].A ;
 wire \l_fifo.genblk1[28].entry.input_buf[3].X ;
 wire \l_fifo.genblk1[28].entry.input_buf[3].genblk1[0].mid ;
 wire \l_fifo.genblk1[28].entry.input_buf[4].A ;
 wire \l_fifo.genblk1[28].entry.input_buf[4].X ;
 wire \l_fifo.genblk1[28].entry.input_buf[4].genblk1[0].mid ;
 wire \l_fifo.genblk1[28].entry.input_buf[5].A ;
 wire \l_fifo.genblk1[28].entry.input_buf[5].X ;
 wire \l_fifo.genblk1[28].entry.input_buf[5].genblk1[0].mid ;
 wire \l_fifo.genblk1[29].entry.empty ;
 wire \l_fifo.genblk1[29].entry.input_buf[0].A ;
 wire \l_fifo.genblk1[29].entry.input_buf[0].X ;
 wire \l_fifo.genblk1[29].entry.input_buf[0].genblk1[0].mid ;
 wire \l_fifo.genblk1[29].entry.input_buf[1].A ;
 wire \l_fifo.genblk1[29].entry.input_buf[1].X ;
 wire \l_fifo.genblk1[29].entry.input_buf[1].genblk1[0].mid ;
 wire \l_fifo.genblk1[29].entry.input_buf[2].A ;
 wire \l_fifo.genblk1[29].entry.input_buf[2].X ;
 wire \l_fifo.genblk1[29].entry.input_buf[2].genblk1[0].mid ;
 wire \l_fifo.genblk1[29].entry.input_buf[3].A ;
 wire \l_fifo.genblk1[29].entry.input_buf[3].X ;
 wire \l_fifo.genblk1[29].entry.input_buf[3].genblk1[0].mid ;
 wire \l_fifo.genblk1[29].entry.input_buf[4].A ;
 wire \l_fifo.genblk1[29].entry.input_buf[4].X ;
 wire \l_fifo.genblk1[29].entry.input_buf[4].genblk1[0].mid ;
 wire \l_fifo.genblk1[29].entry.input_buf[5].A ;
 wire \l_fifo.genblk1[29].entry.input_buf[5].X ;
 wire \l_fifo.genblk1[29].entry.input_buf[5].genblk1[0].mid ;
 wire \l_fifo.genblk1[2].entry.empty ;
 wire \l_fifo.genblk1[2].entry.input_buf[0].A ;
 wire \l_fifo.genblk1[2].entry.input_buf[0].X ;
 wire \l_fifo.genblk1[2].entry.input_buf[0].genblk1[0].mid ;
 wire \l_fifo.genblk1[2].entry.input_buf[1].A ;
 wire \l_fifo.genblk1[2].entry.input_buf[1].X ;
 wire \l_fifo.genblk1[2].entry.input_buf[1].genblk1[0].mid ;
 wire \l_fifo.genblk1[2].entry.input_buf[2].A ;
 wire \l_fifo.genblk1[2].entry.input_buf[2].X ;
 wire \l_fifo.genblk1[2].entry.input_buf[2].genblk1[0].mid ;
 wire \l_fifo.genblk1[2].entry.input_buf[3].A ;
 wire \l_fifo.genblk1[2].entry.input_buf[3].X ;
 wire \l_fifo.genblk1[2].entry.input_buf[3].genblk1[0].mid ;
 wire \l_fifo.genblk1[2].entry.input_buf[4].A ;
 wire \l_fifo.genblk1[2].entry.input_buf[4].X ;
 wire \l_fifo.genblk1[2].entry.input_buf[4].genblk1[0].mid ;
 wire \l_fifo.genblk1[2].entry.input_buf[5].A ;
 wire \l_fifo.genblk1[2].entry.input_buf[5].X ;
 wire \l_fifo.genblk1[2].entry.input_buf[5].genblk1[0].mid ;
 wire \l_fifo.genblk1[30].entry.empty ;
 wire \l_fifo.genblk1[30].entry.input_buf[0].A ;
 wire \l_fifo.genblk1[30].entry.input_buf[0].X ;
 wire \l_fifo.genblk1[30].entry.input_buf[0].genblk1[0].mid ;
 wire \l_fifo.genblk1[30].entry.input_buf[1].A ;
 wire \l_fifo.genblk1[30].entry.input_buf[1].X ;
 wire \l_fifo.genblk1[30].entry.input_buf[1].genblk1[0].mid ;
 wire \l_fifo.genblk1[30].entry.input_buf[2].A ;
 wire \l_fifo.genblk1[30].entry.input_buf[2].X ;
 wire \l_fifo.genblk1[30].entry.input_buf[2].genblk1[0].mid ;
 wire \l_fifo.genblk1[30].entry.input_buf[3].A ;
 wire \l_fifo.genblk1[30].entry.input_buf[3].X ;
 wire \l_fifo.genblk1[30].entry.input_buf[3].genblk1[0].mid ;
 wire \l_fifo.genblk1[30].entry.input_buf[4].A ;
 wire \l_fifo.genblk1[30].entry.input_buf[4].X ;
 wire \l_fifo.genblk1[30].entry.input_buf[4].genblk1[0].mid ;
 wire \l_fifo.genblk1[30].entry.input_buf[5].A ;
 wire \l_fifo.genblk1[30].entry.input_buf[5].X ;
 wire \l_fifo.genblk1[30].entry.input_buf[5].genblk1[0].mid ;
 wire \l_fifo.genblk1[31].entry.empty ;
 wire \l_fifo.genblk1[31].entry.input_buf[0].A ;
 wire \l_fifo.genblk1[31].entry.input_buf[0].X ;
 wire \l_fifo.genblk1[31].entry.input_buf[0].genblk1[0].mid ;
 wire \l_fifo.genblk1[31].entry.input_buf[1].A ;
 wire \l_fifo.genblk1[31].entry.input_buf[1].X ;
 wire \l_fifo.genblk1[31].entry.input_buf[1].genblk1[0].mid ;
 wire \l_fifo.genblk1[31].entry.input_buf[2].A ;
 wire \l_fifo.genblk1[31].entry.input_buf[2].X ;
 wire \l_fifo.genblk1[31].entry.input_buf[2].genblk1[0].mid ;
 wire \l_fifo.genblk1[31].entry.input_buf[3].A ;
 wire \l_fifo.genblk1[31].entry.input_buf[3].X ;
 wire \l_fifo.genblk1[31].entry.input_buf[3].genblk1[0].mid ;
 wire \l_fifo.genblk1[31].entry.input_buf[4].A ;
 wire \l_fifo.genblk1[31].entry.input_buf[4].X ;
 wire \l_fifo.genblk1[31].entry.input_buf[4].genblk1[0].mid ;
 wire \l_fifo.genblk1[31].entry.input_buf[5].A ;
 wire \l_fifo.genblk1[31].entry.input_buf[5].X ;
 wire \l_fifo.genblk1[31].entry.input_buf[5].genblk1[0].mid ;
 wire \l_fifo.genblk1[32].entry.empty ;
 wire \l_fifo.genblk1[32].entry.input_buf[0].A ;
 wire \l_fifo.genblk1[32].entry.input_buf[0].X ;
 wire \l_fifo.genblk1[32].entry.input_buf[0].genblk1[0].mid ;
 wire \l_fifo.genblk1[32].entry.input_buf[1].A ;
 wire \l_fifo.genblk1[32].entry.input_buf[1].X ;
 wire \l_fifo.genblk1[32].entry.input_buf[1].genblk1[0].mid ;
 wire \l_fifo.genblk1[32].entry.input_buf[2].A ;
 wire \l_fifo.genblk1[32].entry.input_buf[2].X ;
 wire \l_fifo.genblk1[32].entry.input_buf[2].genblk1[0].mid ;
 wire \l_fifo.genblk1[32].entry.input_buf[3].A ;
 wire \l_fifo.genblk1[32].entry.input_buf[3].X ;
 wire \l_fifo.genblk1[32].entry.input_buf[3].genblk1[0].mid ;
 wire \l_fifo.genblk1[32].entry.input_buf[4].A ;
 wire \l_fifo.genblk1[32].entry.input_buf[4].X ;
 wire \l_fifo.genblk1[32].entry.input_buf[4].genblk1[0].mid ;
 wire \l_fifo.genblk1[32].entry.input_buf[5].A ;
 wire \l_fifo.genblk1[32].entry.input_buf[5].X ;
 wire \l_fifo.genblk1[32].entry.input_buf[5].genblk1[0].mid ;
 wire \l_fifo.genblk1[33].entry.empty ;
 wire \l_fifo.genblk1[33].entry.input_buf[0].A ;
 wire \l_fifo.genblk1[33].entry.input_buf[0].X ;
 wire \l_fifo.genblk1[33].entry.input_buf[0].genblk1[0].mid ;
 wire \l_fifo.genblk1[33].entry.input_buf[1].A ;
 wire \l_fifo.genblk1[33].entry.input_buf[1].X ;
 wire \l_fifo.genblk1[33].entry.input_buf[1].genblk1[0].mid ;
 wire \l_fifo.genblk1[33].entry.input_buf[2].A ;
 wire \l_fifo.genblk1[33].entry.input_buf[2].X ;
 wire \l_fifo.genblk1[33].entry.input_buf[2].genblk1[0].mid ;
 wire \l_fifo.genblk1[33].entry.input_buf[3].A ;
 wire \l_fifo.genblk1[33].entry.input_buf[3].X ;
 wire \l_fifo.genblk1[33].entry.input_buf[3].genblk1[0].mid ;
 wire \l_fifo.genblk1[33].entry.input_buf[4].A ;
 wire \l_fifo.genblk1[33].entry.input_buf[4].X ;
 wire \l_fifo.genblk1[33].entry.input_buf[4].genblk1[0].mid ;
 wire \l_fifo.genblk1[33].entry.input_buf[5].A ;
 wire \l_fifo.genblk1[33].entry.input_buf[5].X ;
 wire \l_fifo.genblk1[33].entry.input_buf[5].genblk1[0].mid ;
 wire \l_fifo.genblk1[34].entry.empty ;
 wire \l_fifo.genblk1[34].entry.input_buf[0].A ;
 wire \l_fifo.genblk1[34].entry.input_buf[0].X ;
 wire \l_fifo.genblk1[34].entry.input_buf[0].genblk1[0].mid ;
 wire \l_fifo.genblk1[34].entry.input_buf[1].A ;
 wire \l_fifo.genblk1[34].entry.input_buf[1].X ;
 wire \l_fifo.genblk1[34].entry.input_buf[1].genblk1[0].mid ;
 wire \l_fifo.genblk1[34].entry.input_buf[2].A ;
 wire \l_fifo.genblk1[34].entry.input_buf[2].X ;
 wire \l_fifo.genblk1[34].entry.input_buf[2].genblk1[0].mid ;
 wire \l_fifo.genblk1[34].entry.input_buf[3].A ;
 wire \l_fifo.genblk1[34].entry.input_buf[3].X ;
 wire \l_fifo.genblk1[34].entry.input_buf[3].genblk1[0].mid ;
 wire \l_fifo.genblk1[34].entry.input_buf[4].A ;
 wire \l_fifo.genblk1[34].entry.input_buf[4].X ;
 wire \l_fifo.genblk1[34].entry.input_buf[4].genblk1[0].mid ;
 wire \l_fifo.genblk1[34].entry.input_buf[5].A ;
 wire \l_fifo.genblk1[34].entry.input_buf[5].X ;
 wire \l_fifo.genblk1[34].entry.input_buf[5].genblk1[0].mid ;
 wire \l_fifo.genblk1[35].entry.empty ;
 wire \l_fifo.genblk1[35].entry.input_buf[0].A ;
 wire \l_fifo.genblk1[35].entry.input_buf[0].X ;
 wire \l_fifo.genblk1[35].entry.input_buf[0].genblk1[0].mid ;
 wire \l_fifo.genblk1[35].entry.input_buf[1].A ;
 wire \l_fifo.genblk1[35].entry.input_buf[1].X ;
 wire \l_fifo.genblk1[35].entry.input_buf[1].genblk1[0].mid ;
 wire \l_fifo.genblk1[35].entry.input_buf[2].A ;
 wire \l_fifo.genblk1[35].entry.input_buf[2].X ;
 wire \l_fifo.genblk1[35].entry.input_buf[2].genblk1[0].mid ;
 wire \l_fifo.genblk1[35].entry.input_buf[3].A ;
 wire \l_fifo.genblk1[35].entry.input_buf[3].X ;
 wire \l_fifo.genblk1[35].entry.input_buf[3].genblk1[0].mid ;
 wire \l_fifo.genblk1[35].entry.input_buf[4].A ;
 wire \l_fifo.genblk1[35].entry.input_buf[4].X ;
 wire \l_fifo.genblk1[35].entry.input_buf[4].genblk1[0].mid ;
 wire \l_fifo.genblk1[35].entry.input_buf[5].A ;
 wire \l_fifo.genblk1[35].entry.input_buf[5].X ;
 wire \l_fifo.genblk1[35].entry.input_buf[5].genblk1[0].mid ;
 wire \l_fifo.genblk1[36].entry.empty ;
 wire \l_fifo.genblk1[36].entry.input_buf[0].A ;
 wire \l_fifo.genblk1[36].entry.input_buf[0].X ;
 wire \l_fifo.genblk1[36].entry.input_buf[0].genblk1[0].mid ;
 wire \l_fifo.genblk1[36].entry.input_buf[1].A ;
 wire \l_fifo.genblk1[36].entry.input_buf[1].X ;
 wire \l_fifo.genblk1[36].entry.input_buf[1].genblk1[0].mid ;
 wire \l_fifo.genblk1[36].entry.input_buf[2].A ;
 wire \l_fifo.genblk1[36].entry.input_buf[2].X ;
 wire \l_fifo.genblk1[36].entry.input_buf[2].genblk1[0].mid ;
 wire \l_fifo.genblk1[36].entry.input_buf[3].A ;
 wire \l_fifo.genblk1[36].entry.input_buf[3].X ;
 wire \l_fifo.genblk1[36].entry.input_buf[3].genblk1[0].mid ;
 wire \l_fifo.genblk1[36].entry.input_buf[4].A ;
 wire \l_fifo.genblk1[36].entry.input_buf[4].X ;
 wire \l_fifo.genblk1[36].entry.input_buf[4].genblk1[0].mid ;
 wire \l_fifo.genblk1[36].entry.input_buf[5].A ;
 wire \l_fifo.genblk1[36].entry.input_buf[5].X ;
 wire \l_fifo.genblk1[36].entry.input_buf[5].genblk1[0].mid ;
 wire \l_fifo.genblk1[37].entry.empty ;
 wire \l_fifo.genblk1[37].entry.input_buf[0].A ;
 wire \l_fifo.genblk1[37].entry.input_buf[0].X ;
 wire \l_fifo.genblk1[37].entry.input_buf[0].genblk1[0].mid ;
 wire \l_fifo.genblk1[37].entry.input_buf[1].A ;
 wire \l_fifo.genblk1[37].entry.input_buf[1].X ;
 wire \l_fifo.genblk1[37].entry.input_buf[1].genblk1[0].mid ;
 wire \l_fifo.genblk1[37].entry.input_buf[2].A ;
 wire \l_fifo.genblk1[37].entry.input_buf[2].X ;
 wire \l_fifo.genblk1[37].entry.input_buf[2].genblk1[0].mid ;
 wire \l_fifo.genblk1[37].entry.input_buf[3].A ;
 wire \l_fifo.genblk1[37].entry.input_buf[3].X ;
 wire \l_fifo.genblk1[37].entry.input_buf[3].genblk1[0].mid ;
 wire \l_fifo.genblk1[37].entry.input_buf[4].A ;
 wire \l_fifo.genblk1[37].entry.input_buf[4].X ;
 wire \l_fifo.genblk1[37].entry.input_buf[4].genblk1[0].mid ;
 wire \l_fifo.genblk1[37].entry.input_buf[5].A ;
 wire \l_fifo.genblk1[37].entry.input_buf[5].X ;
 wire \l_fifo.genblk1[37].entry.input_buf[5].genblk1[0].mid ;
 wire \l_fifo.genblk1[38].entry.empty ;
 wire \l_fifo.genblk1[38].entry.input_buf[0].A ;
 wire \l_fifo.genblk1[38].entry.input_buf[0].X ;
 wire \l_fifo.genblk1[38].entry.input_buf[0].genblk1[0].mid ;
 wire \l_fifo.genblk1[38].entry.input_buf[1].A ;
 wire \l_fifo.genblk1[38].entry.input_buf[1].X ;
 wire \l_fifo.genblk1[38].entry.input_buf[1].genblk1[0].mid ;
 wire \l_fifo.genblk1[38].entry.input_buf[2].A ;
 wire \l_fifo.genblk1[38].entry.input_buf[2].X ;
 wire \l_fifo.genblk1[38].entry.input_buf[2].genblk1[0].mid ;
 wire \l_fifo.genblk1[38].entry.input_buf[3].A ;
 wire \l_fifo.genblk1[38].entry.input_buf[3].X ;
 wire \l_fifo.genblk1[38].entry.input_buf[3].genblk1[0].mid ;
 wire \l_fifo.genblk1[38].entry.input_buf[4].A ;
 wire \l_fifo.genblk1[38].entry.input_buf[4].X ;
 wire \l_fifo.genblk1[38].entry.input_buf[4].genblk1[0].mid ;
 wire \l_fifo.genblk1[38].entry.input_buf[5].A ;
 wire \l_fifo.genblk1[38].entry.input_buf[5].X ;
 wire \l_fifo.genblk1[38].entry.input_buf[5].genblk1[0].mid ;
 wire \l_fifo.genblk1[39].entry.empty ;
 wire \l_fifo.genblk1[39].entry.input_buf[0].A ;
 wire \l_fifo.genblk1[39].entry.input_buf[0].X ;
 wire \l_fifo.genblk1[39].entry.input_buf[0].genblk1[0].mid ;
 wire \l_fifo.genblk1[39].entry.input_buf[1].A ;
 wire \l_fifo.genblk1[39].entry.input_buf[1].X ;
 wire \l_fifo.genblk1[39].entry.input_buf[1].genblk1[0].mid ;
 wire \l_fifo.genblk1[39].entry.input_buf[2].A ;
 wire \l_fifo.genblk1[39].entry.input_buf[2].X ;
 wire \l_fifo.genblk1[39].entry.input_buf[2].genblk1[0].mid ;
 wire \l_fifo.genblk1[39].entry.input_buf[3].A ;
 wire \l_fifo.genblk1[39].entry.input_buf[3].X ;
 wire \l_fifo.genblk1[39].entry.input_buf[3].genblk1[0].mid ;
 wire \l_fifo.genblk1[39].entry.input_buf[4].A ;
 wire \l_fifo.genblk1[39].entry.input_buf[4].X ;
 wire \l_fifo.genblk1[39].entry.input_buf[4].genblk1[0].mid ;
 wire \l_fifo.genblk1[39].entry.input_buf[5].A ;
 wire \l_fifo.genblk1[39].entry.input_buf[5].X ;
 wire \l_fifo.genblk1[39].entry.input_buf[5].genblk1[0].mid ;
 wire \l_fifo.genblk1[3].entry.empty ;
 wire \l_fifo.genblk1[3].entry.input_buf[0].A ;
 wire \l_fifo.genblk1[3].entry.input_buf[0].X ;
 wire \l_fifo.genblk1[3].entry.input_buf[0].genblk1[0].mid ;
 wire \l_fifo.genblk1[3].entry.input_buf[1].A ;
 wire \l_fifo.genblk1[3].entry.input_buf[1].X ;
 wire \l_fifo.genblk1[3].entry.input_buf[1].genblk1[0].mid ;
 wire \l_fifo.genblk1[3].entry.input_buf[2].A ;
 wire \l_fifo.genblk1[3].entry.input_buf[2].X ;
 wire \l_fifo.genblk1[3].entry.input_buf[2].genblk1[0].mid ;
 wire \l_fifo.genblk1[3].entry.input_buf[3].A ;
 wire \l_fifo.genblk1[3].entry.input_buf[3].X ;
 wire \l_fifo.genblk1[3].entry.input_buf[3].genblk1[0].mid ;
 wire \l_fifo.genblk1[3].entry.input_buf[4].A ;
 wire \l_fifo.genblk1[3].entry.input_buf[4].X ;
 wire \l_fifo.genblk1[3].entry.input_buf[4].genblk1[0].mid ;
 wire \l_fifo.genblk1[3].entry.input_buf[5].A ;
 wire \l_fifo.genblk1[3].entry.input_buf[5].X ;
 wire \l_fifo.genblk1[3].entry.input_buf[5].genblk1[0].mid ;
 wire \l_fifo.genblk1[40].entry.empty ;
 wire \l_fifo.genblk1[40].entry.input_buf[0].A ;
 wire \l_fifo.genblk1[40].entry.input_buf[0].X ;
 wire \l_fifo.genblk1[40].entry.input_buf[0].genblk1[0].mid ;
 wire \l_fifo.genblk1[40].entry.input_buf[1].A ;
 wire \l_fifo.genblk1[40].entry.input_buf[1].X ;
 wire \l_fifo.genblk1[40].entry.input_buf[1].genblk1[0].mid ;
 wire \l_fifo.genblk1[40].entry.input_buf[2].A ;
 wire \l_fifo.genblk1[40].entry.input_buf[2].X ;
 wire \l_fifo.genblk1[40].entry.input_buf[2].genblk1[0].mid ;
 wire \l_fifo.genblk1[40].entry.input_buf[3].A ;
 wire \l_fifo.genblk1[40].entry.input_buf[3].X ;
 wire \l_fifo.genblk1[40].entry.input_buf[3].genblk1[0].mid ;
 wire \l_fifo.genblk1[40].entry.input_buf[4].A ;
 wire \l_fifo.genblk1[40].entry.input_buf[4].X ;
 wire \l_fifo.genblk1[40].entry.input_buf[4].genblk1[0].mid ;
 wire \l_fifo.genblk1[40].entry.input_buf[5].A ;
 wire \l_fifo.genblk1[40].entry.input_buf[5].X ;
 wire \l_fifo.genblk1[40].entry.input_buf[5].genblk1[0].mid ;
 wire \l_fifo.genblk1[41].entry.empty ;
 wire \l_fifo.genblk1[41].entry.input_buf[0].A ;
 wire \l_fifo.genblk1[41].entry.input_buf[0].X ;
 wire \l_fifo.genblk1[41].entry.input_buf[0].genblk1[0].mid ;
 wire \l_fifo.genblk1[41].entry.input_buf[1].A ;
 wire \l_fifo.genblk1[41].entry.input_buf[1].X ;
 wire \l_fifo.genblk1[41].entry.input_buf[1].genblk1[0].mid ;
 wire \l_fifo.genblk1[41].entry.input_buf[2].A ;
 wire \l_fifo.genblk1[41].entry.input_buf[2].X ;
 wire \l_fifo.genblk1[41].entry.input_buf[2].genblk1[0].mid ;
 wire \l_fifo.genblk1[41].entry.input_buf[3].A ;
 wire \l_fifo.genblk1[41].entry.input_buf[3].X ;
 wire \l_fifo.genblk1[41].entry.input_buf[3].genblk1[0].mid ;
 wire \l_fifo.genblk1[41].entry.input_buf[4].A ;
 wire \l_fifo.genblk1[41].entry.input_buf[4].X ;
 wire \l_fifo.genblk1[41].entry.input_buf[4].genblk1[0].mid ;
 wire \l_fifo.genblk1[41].entry.input_buf[5].A ;
 wire \l_fifo.genblk1[41].entry.input_buf[5].X ;
 wire \l_fifo.genblk1[41].entry.input_buf[5].genblk1[0].mid ;
 wire \l_fifo.genblk1[42].entry.empty ;
 wire \l_fifo.genblk1[42].entry.input_buf[0].A ;
 wire \l_fifo.genblk1[42].entry.input_buf[0].X ;
 wire \l_fifo.genblk1[42].entry.input_buf[0].genblk1[0].mid ;
 wire \l_fifo.genblk1[42].entry.input_buf[1].A ;
 wire \l_fifo.genblk1[42].entry.input_buf[1].X ;
 wire \l_fifo.genblk1[42].entry.input_buf[1].genblk1[0].mid ;
 wire \l_fifo.genblk1[42].entry.input_buf[2].A ;
 wire \l_fifo.genblk1[42].entry.input_buf[2].X ;
 wire \l_fifo.genblk1[42].entry.input_buf[2].genblk1[0].mid ;
 wire \l_fifo.genblk1[42].entry.input_buf[3].A ;
 wire \l_fifo.genblk1[42].entry.input_buf[3].X ;
 wire \l_fifo.genblk1[42].entry.input_buf[3].genblk1[0].mid ;
 wire \l_fifo.genblk1[42].entry.input_buf[4].A ;
 wire \l_fifo.genblk1[42].entry.input_buf[4].X ;
 wire \l_fifo.genblk1[42].entry.input_buf[4].genblk1[0].mid ;
 wire \l_fifo.genblk1[42].entry.input_buf[5].A ;
 wire \l_fifo.genblk1[42].entry.input_buf[5].X ;
 wire \l_fifo.genblk1[42].entry.input_buf[5].genblk1[0].mid ;
 wire \l_fifo.genblk1[43].entry.empty ;
 wire \l_fifo.genblk1[43].entry.input_buf[0].A ;
 wire \l_fifo.genblk1[43].entry.input_buf[0].X ;
 wire \l_fifo.genblk1[43].entry.input_buf[0].genblk1[0].mid ;
 wire \l_fifo.genblk1[43].entry.input_buf[1].A ;
 wire \l_fifo.genblk1[43].entry.input_buf[1].X ;
 wire \l_fifo.genblk1[43].entry.input_buf[1].genblk1[0].mid ;
 wire \l_fifo.genblk1[43].entry.input_buf[2].A ;
 wire \l_fifo.genblk1[43].entry.input_buf[2].X ;
 wire \l_fifo.genblk1[43].entry.input_buf[2].genblk1[0].mid ;
 wire \l_fifo.genblk1[43].entry.input_buf[3].A ;
 wire \l_fifo.genblk1[43].entry.input_buf[3].X ;
 wire \l_fifo.genblk1[43].entry.input_buf[3].genblk1[0].mid ;
 wire \l_fifo.genblk1[43].entry.input_buf[4].A ;
 wire \l_fifo.genblk1[43].entry.input_buf[4].X ;
 wire \l_fifo.genblk1[43].entry.input_buf[4].genblk1[0].mid ;
 wire \l_fifo.genblk1[43].entry.input_buf[5].A ;
 wire \l_fifo.genblk1[43].entry.input_buf[5].X ;
 wire \l_fifo.genblk1[43].entry.input_buf[5].genblk1[0].mid ;
 wire \l_fifo.genblk1[44].entry.empty ;
 wire \l_fifo.genblk1[44].entry.input_buf[0].A ;
 wire \l_fifo.genblk1[44].entry.input_buf[0].X ;
 wire \l_fifo.genblk1[44].entry.input_buf[0].genblk1[0].mid ;
 wire \l_fifo.genblk1[44].entry.input_buf[1].A ;
 wire \l_fifo.genblk1[44].entry.input_buf[1].X ;
 wire \l_fifo.genblk1[44].entry.input_buf[1].genblk1[0].mid ;
 wire \l_fifo.genblk1[44].entry.input_buf[2].A ;
 wire \l_fifo.genblk1[44].entry.input_buf[2].X ;
 wire \l_fifo.genblk1[44].entry.input_buf[2].genblk1[0].mid ;
 wire \l_fifo.genblk1[44].entry.input_buf[3].A ;
 wire \l_fifo.genblk1[44].entry.input_buf[3].X ;
 wire \l_fifo.genblk1[44].entry.input_buf[3].genblk1[0].mid ;
 wire \l_fifo.genblk1[44].entry.input_buf[4].A ;
 wire \l_fifo.genblk1[44].entry.input_buf[4].X ;
 wire \l_fifo.genblk1[44].entry.input_buf[4].genblk1[0].mid ;
 wire \l_fifo.genblk1[44].entry.input_buf[5].A ;
 wire \l_fifo.genblk1[44].entry.input_buf[5].X ;
 wire \l_fifo.genblk1[44].entry.input_buf[5].genblk1[0].mid ;
 wire \l_fifo.genblk1[45].entry.empty ;
 wire \l_fifo.genblk1[45].entry.input_buf[0].A ;
 wire \l_fifo.genblk1[45].entry.input_buf[0].X ;
 wire \l_fifo.genblk1[45].entry.input_buf[0].genblk1[0].mid ;
 wire \l_fifo.genblk1[45].entry.input_buf[1].A ;
 wire \l_fifo.genblk1[45].entry.input_buf[1].X ;
 wire \l_fifo.genblk1[45].entry.input_buf[1].genblk1[0].mid ;
 wire \l_fifo.genblk1[45].entry.input_buf[2].A ;
 wire \l_fifo.genblk1[45].entry.input_buf[2].X ;
 wire \l_fifo.genblk1[45].entry.input_buf[2].genblk1[0].mid ;
 wire \l_fifo.genblk1[45].entry.input_buf[3].A ;
 wire \l_fifo.genblk1[45].entry.input_buf[3].X ;
 wire \l_fifo.genblk1[45].entry.input_buf[3].genblk1[0].mid ;
 wire \l_fifo.genblk1[45].entry.input_buf[4].A ;
 wire \l_fifo.genblk1[45].entry.input_buf[4].X ;
 wire \l_fifo.genblk1[45].entry.input_buf[4].genblk1[0].mid ;
 wire \l_fifo.genblk1[45].entry.input_buf[5].A ;
 wire \l_fifo.genblk1[45].entry.input_buf[5].X ;
 wire \l_fifo.genblk1[45].entry.input_buf[5].genblk1[0].mid ;
 wire \l_fifo.genblk1[46].entry.empty ;
 wire \l_fifo.genblk1[46].entry.input_buf[0].A ;
 wire \l_fifo.genblk1[46].entry.input_buf[0].X ;
 wire \l_fifo.genblk1[46].entry.input_buf[0].genblk1[0].mid ;
 wire \l_fifo.genblk1[46].entry.input_buf[1].A ;
 wire \l_fifo.genblk1[46].entry.input_buf[1].X ;
 wire \l_fifo.genblk1[46].entry.input_buf[1].genblk1[0].mid ;
 wire \l_fifo.genblk1[46].entry.input_buf[2].A ;
 wire \l_fifo.genblk1[46].entry.input_buf[2].X ;
 wire \l_fifo.genblk1[46].entry.input_buf[2].genblk1[0].mid ;
 wire \l_fifo.genblk1[46].entry.input_buf[3].A ;
 wire \l_fifo.genblk1[46].entry.input_buf[3].X ;
 wire \l_fifo.genblk1[46].entry.input_buf[3].genblk1[0].mid ;
 wire \l_fifo.genblk1[46].entry.input_buf[4].A ;
 wire \l_fifo.genblk1[46].entry.input_buf[4].X ;
 wire \l_fifo.genblk1[46].entry.input_buf[4].genblk1[0].mid ;
 wire \l_fifo.genblk1[46].entry.input_buf[5].A ;
 wire \l_fifo.genblk1[46].entry.input_buf[5].X ;
 wire \l_fifo.genblk1[46].entry.input_buf[5].genblk1[0].mid ;
 wire \l_fifo.genblk1[47].entry.empty ;
 wire \l_fifo.genblk1[47].entry.input_buf[0].X ;
 wire \l_fifo.genblk1[47].entry.input_buf[0].genblk1[0].mid ;
 wire \l_fifo.genblk1[47].entry.input_buf[1].X ;
 wire \l_fifo.genblk1[47].entry.input_buf[1].genblk1[0].mid ;
 wire \l_fifo.genblk1[47].entry.input_buf[2].X ;
 wire \l_fifo.genblk1[47].entry.input_buf[2].genblk1[0].mid ;
 wire \l_fifo.genblk1[47].entry.input_buf[3].X ;
 wire \l_fifo.genblk1[47].entry.input_buf[3].genblk1[0].mid ;
 wire \l_fifo.genblk1[47].entry.input_buf[4].X ;
 wire \l_fifo.genblk1[47].entry.input_buf[4].genblk1[0].mid ;
 wire \l_fifo.genblk1[47].entry.input_buf[5].X ;
 wire \l_fifo.genblk1[47].entry.input_buf[5].genblk1[0].mid ;
 wire \l_fifo.genblk1[47].entry.write_in ;
 wire \l_fifo.genblk1[4].entry.empty ;
 wire \l_fifo.genblk1[4].entry.input_buf[0].A ;
 wire \l_fifo.genblk1[4].entry.input_buf[0].X ;
 wire \l_fifo.genblk1[4].entry.input_buf[0].genblk1[0].mid ;
 wire \l_fifo.genblk1[4].entry.input_buf[1].A ;
 wire \l_fifo.genblk1[4].entry.input_buf[1].X ;
 wire \l_fifo.genblk1[4].entry.input_buf[1].genblk1[0].mid ;
 wire \l_fifo.genblk1[4].entry.input_buf[2].A ;
 wire \l_fifo.genblk1[4].entry.input_buf[2].X ;
 wire \l_fifo.genblk1[4].entry.input_buf[2].genblk1[0].mid ;
 wire \l_fifo.genblk1[4].entry.input_buf[3].A ;
 wire \l_fifo.genblk1[4].entry.input_buf[3].X ;
 wire \l_fifo.genblk1[4].entry.input_buf[3].genblk1[0].mid ;
 wire \l_fifo.genblk1[4].entry.input_buf[4].A ;
 wire \l_fifo.genblk1[4].entry.input_buf[4].X ;
 wire \l_fifo.genblk1[4].entry.input_buf[4].genblk1[0].mid ;
 wire \l_fifo.genblk1[4].entry.input_buf[5].A ;
 wire \l_fifo.genblk1[4].entry.input_buf[5].X ;
 wire \l_fifo.genblk1[4].entry.input_buf[5].genblk1[0].mid ;
 wire \l_fifo.genblk1[5].entry.empty ;
 wire \l_fifo.genblk1[5].entry.input_buf[0].A ;
 wire \l_fifo.genblk1[5].entry.input_buf[0].X ;
 wire \l_fifo.genblk1[5].entry.input_buf[0].genblk1[0].mid ;
 wire \l_fifo.genblk1[5].entry.input_buf[1].A ;
 wire \l_fifo.genblk1[5].entry.input_buf[1].X ;
 wire \l_fifo.genblk1[5].entry.input_buf[1].genblk1[0].mid ;
 wire \l_fifo.genblk1[5].entry.input_buf[2].A ;
 wire \l_fifo.genblk1[5].entry.input_buf[2].X ;
 wire \l_fifo.genblk1[5].entry.input_buf[2].genblk1[0].mid ;
 wire \l_fifo.genblk1[5].entry.input_buf[3].A ;
 wire \l_fifo.genblk1[5].entry.input_buf[3].X ;
 wire \l_fifo.genblk1[5].entry.input_buf[3].genblk1[0].mid ;
 wire \l_fifo.genblk1[5].entry.input_buf[4].A ;
 wire \l_fifo.genblk1[5].entry.input_buf[4].X ;
 wire \l_fifo.genblk1[5].entry.input_buf[4].genblk1[0].mid ;
 wire \l_fifo.genblk1[5].entry.input_buf[5].A ;
 wire \l_fifo.genblk1[5].entry.input_buf[5].X ;
 wire \l_fifo.genblk1[5].entry.input_buf[5].genblk1[0].mid ;
 wire \l_fifo.genblk1[6].entry.empty ;
 wire \l_fifo.genblk1[6].entry.input_buf[0].A ;
 wire \l_fifo.genblk1[6].entry.input_buf[0].X ;
 wire \l_fifo.genblk1[6].entry.input_buf[0].genblk1[0].mid ;
 wire \l_fifo.genblk1[6].entry.input_buf[1].A ;
 wire \l_fifo.genblk1[6].entry.input_buf[1].X ;
 wire \l_fifo.genblk1[6].entry.input_buf[1].genblk1[0].mid ;
 wire \l_fifo.genblk1[6].entry.input_buf[2].A ;
 wire \l_fifo.genblk1[6].entry.input_buf[2].X ;
 wire \l_fifo.genblk1[6].entry.input_buf[2].genblk1[0].mid ;
 wire \l_fifo.genblk1[6].entry.input_buf[3].A ;
 wire \l_fifo.genblk1[6].entry.input_buf[3].X ;
 wire \l_fifo.genblk1[6].entry.input_buf[3].genblk1[0].mid ;
 wire \l_fifo.genblk1[6].entry.input_buf[4].A ;
 wire \l_fifo.genblk1[6].entry.input_buf[4].X ;
 wire \l_fifo.genblk1[6].entry.input_buf[4].genblk1[0].mid ;
 wire \l_fifo.genblk1[6].entry.input_buf[5].A ;
 wire \l_fifo.genblk1[6].entry.input_buf[5].X ;
 wire \l_fifo.genblk1[6].entry.input_buf[5].genblk1[0].mid ;
 wire \l_fifo.genblk1[7].entry.empty ;
 wire \l_fifo.genblk1[7].entry.input_buf[0].A ;
 wire \l_fifo.genblk1[7].entry.input_buf[0].X ;
 wire \l_fifo.genblk1[7].entry.input_buf[0].genblk1[0].mid ;
 wire \l_fifo.genblk1[7].entry.input_buf[1].A ;
 wire \l_fifo.genblk1[7].entry.input_buf[1].X ;
 wire \l_fifo.genblk1[7].entry.input_buf[1].genblk1[0].mid ;
 wire \l_fifo.genblk1[7].entry.input_buf[2].A ;
 wire \l_fifo.genblk1[7].entry.input_buf[2].X ;
 wire \l_fifo.genblk1[7].entry.input_buf[2].genblk1[0].mid ;
 wire \l_fifo.genblk1[7].entry.input_buf[3].A ;
 wire \l_fifo.genblk1[7].entry.input_buf[3].X ;
 wire \l_fifo.genblk1[7].entry.input_buf[3].genblk1[0].mid ;
 wire \l_fifo.genblk1[7].entry.input_buf[4].A ;
 wire \l_fifo.genblk1[7].entry.input_buf[4].X ;
 wire \l_fifo.genblk1[7].entry.input_buf[4].genblk1[0].mid ;
 wire \l_fifo.genblk1[7].entry.input_buf[5].A ;
 wire \l_fifo.genblk1[7].entry.input_buf[5].X ;
 wire \l_fifo.genblk1[7].entry.input_buf[5].genblk1[0].mid ;
 wire \l_fifo.genblk1[8].entry.empty ;
 wire \l_fifo.genblk1[8].entry.input_buf[0].A ;
 wire \l_fifo.genblk1[8].entry.input_buf[0].X ;
 wire \l_fifo.genblk1[8].entry.input_buf[0].genblk1[0].mid ;
 wire \l_fifo.genblk1[8].entry.input_buf[1].A ;
 wire \l_fifo.genblk1[8].entry.input_buf[1].X ;
 wire \l_fifo.genblk1[8].entry.input_buf[1].genblk1[0].mid ;
 wire \l_fifo.genblk1[8].entry.input_buf[2].A ;
 wire \l_fifo.genblk1[8].entry.input_buf[2].X ;
 wire \l_fifo.genblk1[8].entry.input_buf[2].genblk1[0].mid ;
 wire \l_fifo.genblk1[8].entry.input_buf[3].A ;
 wire \l_fifo.genblk1[8].entry.input_buf[3].X ;
 wire \l_fifo.genblk1[8].entry.input_buf[3].genblk1[0].mid ;
 wire \l_fifo.genblk1[8].entry.input_buf[4].A ;
 wire \l_fifo.genblk1[8].entry.input_buf[4].X ;
 wire \l_fifo.genblk1[8].entry.input_buf[4].genblk1[0].mid ;
 wire \l_fifo.genblk1[8].entry.input_buf[5].A ;
 wire \l_fifo.genblk1[8].entry.input_buf[5].X ;
 wire \l_fifo.genblk1[8].entry.input_buf[5].genblk1[0].mid ;
 wire \l_fifo.genblk1[9].entry.input_buf[0].A ;
 wire \l_fifo.genblk1[9].entry.input_buf[0].X ;
 wire \l_fifo.genblk1[9].entry.input_buf[0].genblk1[0].mid ;
 wire \l_fifo.genblk1[9].entry.input_buf[1].A ;
 wire \l_fifo.genblk1[9].entry.input_buf[1].X ;
 wire \l_fifo.genblk1[9].entry.input_buf[1].genblk1[0].mid ;
 wire \l_fifo.genblk1[9].entry.input_buf[2].A ;
 wire \l_fifo.genblk1[9].entry.input_buf[2].X ;
 wire \l_fifo.genblk1[9].entry.input_buf[2].genblk1[0].mid ;
 wire \l_fifo.genblk1[9].entry.input_buf[3].A ;
 wire \l_fifo.genblk1[9].entry.input_buf[3].X ;
 wire \l_fifo.genblk1[9].entry.input_buf[3].genblk1[0].mid ;
 wire \l_fifo.genblk1[9].entry.input_buf[4].A ;
 wire \l_fifo.genblk1[9].entry.input_buf[4].X ;
 wire \l_fifo.genblk1[9].entry.input_buf[4].genblk1[0].mid ;
 wire \l_fifo.genblk1[9].entry.input_buf[5].A ;
 wire \l_fifo.genblk1[9].entry.input_buf[5].X ;
 wire \l_fifo.genblk1[9].entry.input_buf[5].genblk1[0].mid ;
 wire \l_fifo.ready ;
 wire net1;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net2;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net3;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net4;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire reset_n_in;
 wire [0:0] clknet_0_io_in;
 wire [0:0] clknet_3_0__leaf_io_in;
 wire [0:0] clknet_3_1__leaf_io_in;
 wire [0:0] clknet_3_2__leaf_io_in;
 wire [0:0] clknet_3_3__leaf_io_in;
 wire [0:0] clknet_3_4__leaf_io_in;
 wire [0:0] clknet_3_5__leaf_io_in;
 wire [0:0] clknet_3_6__leaf_io_in;
 wire [0:0] clknet_3_7__leaf_io_in;

 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(_005_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_10 (.DIODE(_056_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_11 (.DIODE(_078_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_12 (.DIODE(_081_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_13 (.DIODE(_083_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_14 (.DIODE(\l_fifo.genblk1[2].entry.input_buf[5].X ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_15 (.DIODE(_000_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_16 (.DIODE(\l_fifo.genblk1[47].entry.input_buf[5].X ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(_008_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_3 (.DIODE(_034_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_4 (.DIODE(_037_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_5 (.DIODE(_042_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_6 (.DIODE(_043_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_7 (.DIODE(_049_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_8 (.DIODE(_050_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_9 (.DIODE(_055_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_101 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_110 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_0_113 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_121 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_125 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_137 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_141 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_153 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_165 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_169 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_181 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_193 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_197 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_209 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_0_21 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_221 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_225 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_232 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_239 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_0_246 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_253 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_258 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_0_265 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_27 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_273 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_278 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_281 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_0_286 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_29 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_292 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_296 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_41 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_53 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_57 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_69 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_75 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_82 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_85 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_0_92 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_10_102 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_10_113 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_10_128 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_10_132 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_10_138 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_10_141 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_10_162 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_10_179 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_10_186 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_10_193 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_10_197 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_10_216 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_10_22 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_10_223 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_10_230 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_10_237 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_10_245 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_10_250 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_10_253 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_10_257 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_10_271 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_10_278 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_10_285 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_10_29 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_10_292 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_10_298 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_10_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_10_48 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_10_60 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_10_72 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_10_76 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_10_82 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_10_85 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_10_94 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_11_110 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_11_113 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_11_119 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_11_127 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_11_138 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_11_144 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_11_15 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_11_152 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_11_161 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_11_167 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_11_169 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_11_174 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_11_178 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_11_192 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_11_209 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_11_216 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_11_225 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_11_229 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_11_243 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_11_247 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_11_251 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_11_270 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_11_277 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_11_281 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_11_286 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_11_293 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_11_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_11_36 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_11_48 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_11_57 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_11_69 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_11_77 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_11_83 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_11_95 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_12_102 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_12_106 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_12_114 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_12_121 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_12_132 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_12_141 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_12_150 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_12_157 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_12_174 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_12_181 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_12_188 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_12_197 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_12_203 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_12_224 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_12_241 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_12_25 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_12_250 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_12_253 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_12_268 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_12_287 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_12_29 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_12_294 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_12_298 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_12_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_12_43 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_12_65 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_12_7 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_12_77 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_12_83 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_12_85 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_12_91 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_12_98 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_13_105 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_13_110 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_13_113 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_13_121 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_13_133 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_13_140 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_13_144 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_13_158 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_13_165 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_13_169 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_13_175 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_13_192 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_13_209 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_13_216 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_13_225 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_13_230 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_13_249 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_13_256 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_13_26 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_13_265 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_13_272 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_13_281 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_13_286 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_13_293 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_13_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_13_46 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_13_54 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_13_57 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_13_76 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_13_88 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_13_97 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_14_102 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_14_113 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_14_121 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_14_126 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_14_137 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_14_141 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_14_148 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_14_157 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_14_174 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_14_178 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_14_182 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_14_189 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_14_195 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_14_197 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_14_202 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_14_21 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_14_219 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_14_226 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_14_243 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_14_25 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_14_250 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_14_253 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_14_268 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_14_285 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_14_29 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_14_292 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_14_298 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_14_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_14_41 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_14_59 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_14_82 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_14_85 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_14_97 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_15_105 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_15_111 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_15_113 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_15_122 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_15_128 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_15_134 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_15_143 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_15_147 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_15_151 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_15_158 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_15_166 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_15_169 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_15_182 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_15_186 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_15_20 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_15_200 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_15_217 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_15_223 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_15_225 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_15_24 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_15_240 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_15_257 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_15_276 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_15_281 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_15_296 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_15_43 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_15_55 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_15_57 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_15_65 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_15_84 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_16_106 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_16_115 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_16_125 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_16_138 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_16_141 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_16_150 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_16_158 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_16_162 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_16_169 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_16_190 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_16_197 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_16_213 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_16_221 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_16_23 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_16_235 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_16_249 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_16_253 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_16_258 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_16_265 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_16_27 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_16_272 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_16_280 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_16_29 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_16_297 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_16_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_16_50 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_16_54 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_16_72 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_16_85 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_16_97 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_17_105 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_17_110 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_17_113 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_17_120 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_17_131 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_17_138 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_17_145 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_17_152 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_17_159 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_17_166 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_17_169 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_17_184 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_17_191 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_17_195 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_17_199 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_17_20 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_17_206 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_17_213 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_17_220 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_17_225 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_17_235 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_17_239 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_17_24 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_17_253 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_17_257 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_17_271 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_17_278 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_17_281 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_17_286 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_17_293 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_17_43 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_17_50 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_17_57 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_17_69 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_17_81 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_17_93 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_18_101 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_18_107 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_18_116 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_18_126 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_18_138 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_18_141 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_18_149 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_18_153 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_18_159 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_18_165 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_18_169 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_18_177 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_18_191 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_18_195 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_18_197 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_18_212 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_18_219 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_18_22 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_18_225 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_18_239 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_18_246 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_18_253 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_18_259 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_18_26 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_18_273 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_18_280 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_18_287 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_18_29 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_18_294 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_18_298 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_18_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_18_41 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_18_48 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_18_55 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_18_62 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_18_74 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_18_82 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_18_85 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_18_97 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_19_107 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_19_111 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_19_113 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_19_121 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_19_127 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_19_135 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_19_139 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_19_148 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_19_157 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_19_166 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_19_169 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_19_184 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_19_201 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_19_218 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_19_225 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_19_230 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_19_236 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_19_25 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_19_250 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_19_254 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_19_268 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_19_275 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_19_279 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_19_281 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_19_296 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_19_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_19_32 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_19_54 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_19_57 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_19_7 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_19_75 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_19_83 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_19_90 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_1_110 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_1_113 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_1_122 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_1_133 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_1_145 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_1_151 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_1_159 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_1_167 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_1_169 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_1_174 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_1_186 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_1_198 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_1_210 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_1_218 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_1_22 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_1_222 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_1_225 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_1_236 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_1_243 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_1_249 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_1_253 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_1_260 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_1_267 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_1_278 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_1_281 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_1_286 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_1_295 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_1_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_1_34 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_1_54 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_1_57 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_1_65 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_1_85 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_1_93 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_1_99 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_20_104 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_20_110 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_20_118 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_20_122 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_20_131 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_20_138 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_20_141 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_20_147 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_20_153 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_20_162 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_20_174 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_20_181 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_20_188 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_20_197 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_20_202 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_20_210 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_20_224 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_20_24 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_20_241 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_20_248 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_20_253 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_20_258 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_20_265 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_20_284 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_20_29 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_20_291 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_20_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_20_36 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_20_55 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_20_75 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_20_82 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_20_85 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_20_95 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_20_99 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_21_109 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_21_113 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_21_120 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_21_130 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_21_136 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_21_142 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_21_151 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_21_155 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_21_161 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_21_167 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_21_169 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_21_190 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_21_197 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_21_216 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_21_225 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_21_229 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_21_234 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_21_24 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_21_241 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_21_260 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_21_267 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_21_274 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_21_281 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_21_286 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_21_293 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_21_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_21_30 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_21_48 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_21_57 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_21_63 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_21_80 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_21_88 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_21_99 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_22_103 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_22_109 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_22_121 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_22_138 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_22_141 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_22_155 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_22_172 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_22_178 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_22_192 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_22_197 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_22_214 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_22_218 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_22_232 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_22_249 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_22_25 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_22_253 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_22_258 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_22_265 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_22_273 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_22_288 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_22_29 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_22_295 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_22_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_22_34 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_22_41 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_22_65 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_22_74 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_22_82 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_22_85 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_22_95 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_23_102 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_23_108 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_23_113 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_23_120 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_23_131 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_23_140 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_23_144 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_23_154 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_23_162 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_23_166 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_23_169 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_23_184 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_23_191 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_23_198 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_23_205 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_23_212 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_23_219 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_23_223 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_23_225 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_23_24 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_23_240 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_23_244 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_23_258 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_23_275 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_23_279 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_23_281 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_23_286 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_23_292 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_23_296 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_23_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_23_45 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_23_52 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_23_57 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_23_61 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_23_79 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_23_83 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_23_88 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_23_98 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_24_108 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_24_116 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_24_125 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_24_133 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_24_138 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_24_141 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_24_147 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_24_151 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_24_155 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_24_172 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_24_183 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_24_190 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_24_197 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_24_212 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_24_22 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_24_229 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_24_246 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_24_253 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_24_258 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_24_266 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_24_280 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_24_287 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_24_29 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_24_294 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_24_298 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_24_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_24_34 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_24_42 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_24_59 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_24_66 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_24_73 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_24_82 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_24_85 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_24_99 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_25_110 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_25_113 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_25_117 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_25_123 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_25_13 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_25_131 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_25_136 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_25_143 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_25_152 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_25_159 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_25_166 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_25_169 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_25_174 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_25_193 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_25_200 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_25_207 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_25_214 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_25_221 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_25_225 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_25_230 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_25_237 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_25_244 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_25_251 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_25_258 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_25_265 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_25_272 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_25_281 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_25_286 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_25_293 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_25_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_25_34 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_25_54 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_25_57 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_25_77 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_25_9 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_25_91 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_25_98 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_26_105 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_26_113 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_26_121 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_26_138 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_26_141 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_26_152 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_26_160 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_26_177 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_26_184 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_26_191 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_26_195 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_26_197 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_26_212 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_26_216 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_26_230 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_26_237 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_26_244 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_26_253 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_26_258 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_26_26 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_26_266 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_26_281 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_26_288 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_26_29 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_26_295 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_26_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_26_34 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_26_41 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_26_65 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_26_71 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_26_75 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_26_8 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_26_82 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_26_85 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_26_92 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_26_96 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_27_100 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_27_108 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_27_113 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_27_124 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_27_143 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_27_147 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_27_161 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_27_167 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_27_169 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_27_184 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_27_191 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_27_198 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_27_202 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_27_216 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_27_225 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_27_229 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_27_243 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_27_25 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_27_250 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_27_254 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_27_268 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_27_275 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_27_279 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_27_281 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_27_286 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_27_293 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_27_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_27_33 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_27_51 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_27_55 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_27_57 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_27_75 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_27_84 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_27_92 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_28_103 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_28_121 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_28_138 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_28_141 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_28_147 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_28_161 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_28_169 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_28_188 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_28_197 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_28_202 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_28_21 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_28_219 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_28_226 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_28_233 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_28_250 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_28_253 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_28_268 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_28_27 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_28_275 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_28_282 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_28_289 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_28_29 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_28_296 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_28_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_28_34 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_28_40 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_28_61 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_28_82 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_28_85 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_28_94 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_29_107 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_29_111 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_29_113 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_29_123 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_29_142 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_29_159 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_29_166 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_29_169 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_29_184 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_29_190 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_29_204 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_29_21 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_29_221 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_29_225 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_29_231 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_29_239 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_29_246 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_29_253 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_29_272 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_29_28 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_29_281 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_29_296 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_29_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_29_52 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_29_57 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_29_65 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_29_82 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_29_90 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_2_103 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_2_111 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_2_115 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_2_121 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_2_130 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_2_138 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_2_141 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_2_147 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_2_159 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_2_168 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_2_180 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_2_187 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_2_195 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_2_197 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_2_209 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_2_21 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_2_213 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_2_217 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_2_224 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_2_233 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_2_240 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_2_247 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_2_251 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_2_253 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_2_259 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_2_266 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_2_27 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_2_270 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_2_274 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_2_278 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_2_282 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_2_29 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_2_293 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_2_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_2_48 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_2_69 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_2_82 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_2_85 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_2_90 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_2_94 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_30_106 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_30_110 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_30_117 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_30_124 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_30_131 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_30_138 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_30_141 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_30_148 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_30_156 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_30_171 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_30_178 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_30_185 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_30_192 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_30_197 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_30_202 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_30_208 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_30_212 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_30_22 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_30_220 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_30_235 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_30_243 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_30_250 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_30_253 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_30_268 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_30_285 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_30_29 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_30_292 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_30_298 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_30_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_30_34 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_30_38 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_30_55 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_30_59 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_30_63 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_30_70 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_30_81 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_30_85 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_30_98 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_31_109 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_31_113 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_31_119 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_31_123 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_31_140 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_31_144 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_31_148 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_31_155 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_31_162 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_31_169 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_31_174 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_31_181 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_31_188 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_31_195 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_31_201 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_31_21 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_31_215 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_31_222 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_31_225 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_31_246 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_31_25 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_31_253 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_31_260 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_31_267 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_31_274 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_31_281 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_31_286 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_31_293 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_31_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_31_43 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_31_54 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_31_57 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_31_64 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_31_74 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_31_91 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_31_98 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_32_100 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_32_108 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_32_125 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_32_133 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_32_138 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_32_141 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_32_145 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_32_159 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_32_163 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_32_177 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_32_194 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_32_197 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_32_21 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_32_212 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_32_231 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_32_250 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_32_253 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_32_259 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_32_27 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_32_273 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_32_29 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_32_292 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_32_298 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_32_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_32_34 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_32_41 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_32_62 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_32_73 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_32_82 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_32_85 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_33_101 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_33_109 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_33_113 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_33_119 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_33_125 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_33_139 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_33_156 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_33_165 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_33_169 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_33_184 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_33_191 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_33_198 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_33_205 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_33_212 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_33_219 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_33_223 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_33_225 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_33_24 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_33_240 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_33_248 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_33_255 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_33_263 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_33_277 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_33_281 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_33_286 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_33_293 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_33_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_33_44 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_33_50 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_33_54 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_33_57 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_33_69 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_33_76 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_33_87 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_33_95 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_34_105 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_34_122 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_34_133 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_34_139 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_34_141 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_34_146 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_34_152 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_34_156 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_34_164 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_34_172 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_34_187 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_34_194 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_34_197 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_34_202 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_34_208 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_34_22 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_34_222 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_34_240 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_34_247 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_34_251 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_34_253 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_34_268 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_34_275 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_34_282 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_34_289 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_34_29 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_34_296 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_34_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_34_36 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_34_44 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_34_62 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_34_78 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_34_85 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_34_98 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_35_110 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_35_113 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_35_118 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_35_135 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_35_142 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_35_148 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_35_162 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_35_169 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_35_184 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_35_205 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_35_22 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_35_222 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_35_225 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_35_241 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_35_258 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_35_274 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_35_281 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_35_297 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_35_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_35_42 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_35_50 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_35_54 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_35_57 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_35_76 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_35_88 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_35_96 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_36_102 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_36_119 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_36_136 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_36_141 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_36_156 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_36_164 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_36_185 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_36_192 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_36_197 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_36_202 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_36_209 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_36_230 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_36_236 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_36_241 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_36_248 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_36_25 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_36_253 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_36_257 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_36_271 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_36_288 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_36_29 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_36_295 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_36_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_36_34 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_36_41 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_36_65 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_36_72 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_36_82 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_36_85 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_37_101 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_37_110 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_37_113 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_37_122 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_37_128 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_37_132 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_37_139 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_37_143 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_37_147 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_37_166 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_37_169 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_37_174 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_37_182 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_37_196 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_37_20 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_37_203 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_37_207 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_37_221 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_37_225 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_37_24 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_37_240 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_37_246 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_37_260 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_37_267 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_37_274 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_37_281 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_37_297 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_37_42 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_37_50 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_37_54 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_37_57 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_37_66 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_37_74 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_37_83 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_37_94 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_38_109 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_38_113 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_38_127 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_38_138 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_38_141 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_38_148 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_38_155 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_38_162 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_38_170 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_38_191 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_38_195 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_38_197 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_38_218 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_38_22 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_38_225 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_38_232 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_38_236 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_38_250 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_38_253 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_38_258 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_38_265 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_38_272 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_38_289 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_38_29 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_38_296 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_38_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_38_35 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_38_52 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_38_72 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_38_78 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_38_82 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_38_85 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_38_94 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_39_104 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_39_113 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_39_119 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_39_126 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_39_133 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_39_140 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_39_147 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_39_166 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_39_169 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_39_185 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_39_206 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_39_214 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_39_221 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_39_225 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_39_230 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_39_237 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_39_244 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_39_251 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_39_270 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_39_277 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_39_281 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_39_296 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_39_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_39_30 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_39_54 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_39_57 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_39_62 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_39_72 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_39_76 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_39_80 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_39_89 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_39_9 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_3_109 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_3_113 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_3_122 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_3_130 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_3_136 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_3_144 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_3_15 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_3_159 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_3_166 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_3_169 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_3_177 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_3_183 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_3_194 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_3_201 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_3_208 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_3_215 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_3_222 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_3_225 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_3_241 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_3_249 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_3_264 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_3_273 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_3_279 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_3_281 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_3_286 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_3_293 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_3_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_3_34 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_3_46 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_3_54 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_3_57 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_3_69 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_3_77 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_3_82 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_3_94 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_40_100 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_40_104 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_40_110 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_40_12 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_40_121 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_40_138 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_40_141 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_40_156 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_40_162 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_40_176 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_40_183 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_40_19 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_40_190 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_40_197 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_40_202 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_40_209 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_40_213 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_40_227 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_40_234 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_40_241 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_40_248 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_40_253 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_40_258 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_40_26 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_40_265 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_40_284 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_40_29 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_40_291 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_40_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_40_35 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_40_47 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_40_54 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_40_62 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_40_66 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_40_73 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_40_82 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_40_85 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_40_91 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_41_106 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_41_113 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_41_12 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_41_128 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_41_132 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_41_136 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_41_142 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_41_146 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_41_153 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_41_160 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_41_169 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_41_174 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_41_181 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_41_185 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_41_189 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_41_197 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_41_20 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_41_211 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_41_218 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_41_225 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_41_24 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_41_244 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_41_261 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_41_267 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_41_27 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_41_271 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_41_278 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_41_281 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_41_286 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_41_297 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_41_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_41_46 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_41_53 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_41_57 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_41_66 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_41_87 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_41_94 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_42_100 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_42_108 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_42_119 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_42_127 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_42_133 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_42_139 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_42_141 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_42_146 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_42_153 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_42_170 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_42_177 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_42_184 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_42_191 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_42_195 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_42_197 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_42_202 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_42_209 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_42_21 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_42_226 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_42_233 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_42_240 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_42_247 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_42_251 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_42_253 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_42_258 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_42_264 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_42_268 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_42_27 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_42_276 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_42_29 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_42_290 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_42_297 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_42_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_42_34 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_42_42 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_42_60 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_42_67 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_42_71 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_42_75 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_42_82 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_42_85 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_43_103 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_43_110 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_43_113 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_43_117 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_43_12 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_43_131 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_43_148 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_43_152 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_43_166 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_43_169 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_43_185 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_43_19 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_43_192 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_43_199 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_43_203 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_43_217 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_43_223 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_43_225 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_43_240 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_43_257 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_43_278 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_43_28 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_43_281 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_43_286 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_43_293 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_43_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_43_36 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_43_40 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_43_47 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_43_54 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_43_57 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_43_63 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_43_67 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_43_76 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_43_83 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_43_92 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_44_100 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_44_121 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_44_138 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_44_141 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_44_157 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_44_161 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_44_165 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_44_172 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_44_179 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_44_186 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_44_193 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_44_197 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_44_212 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_44_219 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_44_226 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_44_23 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_44_233 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_44_241 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_44_249 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_44_253 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_44_27 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_44_270 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_44_277 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_44_284 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_44_29 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_44_291 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_44_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_44_52 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_44_61 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_44_68 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_44_75 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_44_82 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_44_85 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_45_101 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_45_110 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_45_113 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_45_128 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_45_145 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_45_152 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_45_16 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_45_160 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_45_165 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_45_169 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_45_184 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_45_191 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_45_197 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_45_211 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_45_218 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_45_225 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_45_230 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_45_237 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_45_244 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_45_248 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_45_25 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_45_262 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_45_269 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_45_276 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_45_281 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_45_286 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_45_293 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_45_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_45_37 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_45_43 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_45_47 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_45_54 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_45_57 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_45_64 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_45_75 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_45_8 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_45_84 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_46_116 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_46_122 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_46_126 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_46_133 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_46_139 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_46_141 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_46_147 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_46_15 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_46_151 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_46_159 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_46_165 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_46_172 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_46_180 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_46_194 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_46_197 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_46_201 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_46_215 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_46_22 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_46_232 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_46_249 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_46_253 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_46_258 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_46_264 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_46_278 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_46_285 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_46_29 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_46_292 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_46_298 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_46_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_46_45 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_46_60 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_46_73 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_46_82 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_46_85 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_46_9 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_46_91 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_46_99 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_47_103 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_47_110 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_47_113 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_47_119 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_47_133 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_47_141 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_47_146 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_47_163 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_47_167 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_47_169 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_47_174 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_47_182 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_47_186 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_47_193 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_47_200 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_47_207 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_47_21 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_47_214 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_47_221 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_47_225 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_47_242 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_47_263 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_47_270 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_47_277 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_47_281 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_47_296 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_47_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_47_37 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_47_48 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_47_57 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_47_64 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_47_68 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_47_76 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_47_93 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_47_99 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_48_100 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_48_117 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_48_126 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_48_133 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_48_139 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_48_141 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_48_156 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_48_160 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_48_165 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_48_172 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_48_179 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_48_186 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_48_193 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_48_197 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_48_212 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_48_229 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_48_235 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_48_24 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_48_249 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_48_253 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_48_258 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_48_266 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_48_280 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_48_289 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_48_29 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_48_296 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_48_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_48_34 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_48_41 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_48_52 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_48_59 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_48_65 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_48_69 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_48_80 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_48_85 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_49_103 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_49_110 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_49_113 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_49_119 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_49_12 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_49_123 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_49_140 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_49_147 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_49_164 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_49_169 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_49_175 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_49_18 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_49_189 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_49_196 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_49_203 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_49_210 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_49_217 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_49_223 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_49_225 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_49_240 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_49_248 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_49_262 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_49_269 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_49_27 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_49_276 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_49_281 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_49_286 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_49_292 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_49_296 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_49_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_49_34 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_49_42 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_49_47 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_49_54 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_49_57 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_49_62 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_49_8 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_49_83 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_49_91 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_49_96 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_4_105 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_4_116 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_4_123 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_4_134 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_4_141 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_4_150 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_4_171 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_4_188 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_4_197 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_4_212 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_4_22 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_4_229 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_4_236 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_4_243 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_4_250 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_4_253 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_4_258 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_4_265 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_4_282 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_4_289 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_4_29 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_4_296 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_4_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_4_41 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_4_53 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_4_65 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_4_82 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_4_85 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_4_95 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_4_99 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_50_101 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_50_118 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_50_130 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_50_134 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_50_138 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_50_141 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_50_156 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_50_163 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_50_167 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_50_181 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_50_188 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_50_197 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_50_212 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_50_229 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_50_246 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_50_253 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_50_258 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_50_26 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_50_265 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_50_272 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_50_279 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_50_286 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_50_29 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_50_293 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_50_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_50_40 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_50_47 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_50_54 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_50_61 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_50_82 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_50_85 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_50_9 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_51_103 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_51_110 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_51_113 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_51_12 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_51_129 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_51_135 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_51_149 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_51_166 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_51_169 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_51_175 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_51_183 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_51_197 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_51_216 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_51_225 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_51_230 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_51_237 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_51_254 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_51_27 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_51_271 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_51_278 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_51_281 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_51_286 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_51_293 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_51_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_51_44 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_51_50 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_51_54 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_51_57 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_51_66 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_51_73 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_51_8 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_51_85 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_51_96 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_52_100 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_52_104 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_52_118 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_52_124 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_52_138 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_52_14 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_52_141 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_52_146 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_52_154 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_52_159 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_52_166 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_52_18 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_52_183 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_52_190 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_52_197 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_52_203 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_52_211 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_52_225 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_52_242 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_52_249 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_52_253 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_52_258 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_52_26 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_52_265 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_52_272 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_52_279 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_52_286 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_52_29 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_52_293 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_52_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_52_33 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_52_44 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_52_58 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_52_65 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_52_8 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_52_82 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_52_85 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_53_108 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_53_113 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_53_132 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_53_149 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_53_155 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_53_159 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_53_166 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_53_169 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_53_175 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_53_189 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_53_196 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_53_21 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_53_215 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_53_222 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_53_225 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_53_230 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_53_237 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_53_244 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_53_252 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_53_266 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_53_273 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_53_279 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_53_281 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_53_286 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_53_293 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_53_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_53_40 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_53_47 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_53_54 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_53_57 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_53_68 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_53_7 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_53_85 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_53_93 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_54_107 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_54_111 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_54_118 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_54_125 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_54_133 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_54_138 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_54_141 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_54_157 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_54_16 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_54_174 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_54_181 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_54_188 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_54_197 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_54_212 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_54_219 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_54_22 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_54_226 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_54_232 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_54_246 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_54_253 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_54_258 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_54_26 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_54_265 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_54_272 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_54_279 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_54_286 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_54_29 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_54_293 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_54_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_54_34 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_54_38 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_54_52 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_54_69 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_54_77 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_54_82 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_54_85 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_54_9 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_54_91 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_54_99 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_55_10 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_55_105 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_55_110 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_55_113 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_55_128 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_55_132 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_55_136 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_55_14 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_55_140 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_55_144 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_55_150 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_55_154 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_55_161 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_55_167 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_55_169 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_55_174 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_55_18 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_55_181 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_55_198 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_55_204 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_55_218 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_55_225 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_55_230 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_55_237 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_55_244 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_55_251 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_55_258 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_55_26 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_55_265 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_55_272 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_55_281 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_55_286 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_55_293 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_55_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_55_41 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_55_49 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_55_54 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_55_57 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_55_76 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_55_97 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_56_103 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_56_11 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_56_120 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_56_137 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_56_141 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_56_147 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_56_15 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_56_151 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_56_168 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_56_172 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_56_186 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_56_19 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_56_193 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_56_197 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_56_213 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_56_220 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_56_227 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_56_231 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_56_245 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_56_251 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_56_253 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_56_258 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_56_26 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_56_265 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_56_272 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_56_279 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_56_286 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_56_29 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_56_293 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_56_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_56_38 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_56_45 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_56_62 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_56_67 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_56_7 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_56_82 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_56_85 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_56_89 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_57_103 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_57_110 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_57_113 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_57_119 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_57_12 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_57_126 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_57_134 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_57_138 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_57_141 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_57_146 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_57_150 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_57_154 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_57_162 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_57_166 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_57_169 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_57_174 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_57_178 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_57_182 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_57_19 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_57_190 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_57_194 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_57_197 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_57_202 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_57_210 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_57_215 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_57_222 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_57_225 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_57_230 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_57_237 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_57_244 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_57_253 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_57_258 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_57_26 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_57_265 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_57_272 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_57_281 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_57_286 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_57_29 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_57_293 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_57_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_57_40 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_57_47 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_57_54 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_57_57 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_57_68 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_57_75 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_57_82 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_57_85 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_57_96 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_5_108 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_5_113 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_5_117 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_5_125 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_5_138 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_5_149 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_5_15 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_5_155 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_5_159 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_5_166 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_5_169 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_5_173 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_5_187 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_5_194 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_5_201 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_5_208 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_5_215 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_5_222 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_5_225 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_5_240 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_5_247 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_5_254 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_5_258 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_5_272 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_5_281 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_5_286 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_5_295 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_5_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_5_32 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_5_44 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_5_57 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_5_68 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_5_79 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_5_9 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_5_90 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_5_97 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_6_100 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_6_113 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_6_117 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_6_126 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_6_133 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_6_139 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_6_141 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_6_148 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_6_165 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_6_172 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_6_179 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_6_186 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_6_193 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_6_197 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_6_203 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_6_207 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_6_214 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_6_221 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_6_229 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_6_234 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_6_241 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_6_250 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_6_253 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_6_258 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_6_26 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_6_277 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_6_285 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_6_289 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_6_29 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_6_296 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_6_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_6_33 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_6_52 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_6_61 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_6_82 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_6_85 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_6_9 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_7_101 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_7_109 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_7_113 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_7_119 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_7_125 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_7_136 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_7_147 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_7_166 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_7_169 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_7_188 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_7_195 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_7_202 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_7_208 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_7_222 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_7_225 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_7_229 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_7_233 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_7_237 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_7_25 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_7_251 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_7_268 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_7_275 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_7_279 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_7_281 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_7_297 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_7_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_7_37 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_7_54 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_7_57 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_7_63 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_7_82 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_7_93 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_8_108 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_8_114 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_8_123 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_8_134 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_8_141 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_8_148 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_8_152 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_8_156 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_8_163 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_8_171 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_8_178 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_8_182 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_8_186 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_8_193 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_8_197 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_8_213 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_8_22 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_8_230 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_8_237 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_8_246 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_8_253 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_8_258 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_8_265 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_8_286 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_8_29 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_8_293 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_8_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_8_41 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_8_49 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_8_69 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_8_82 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_8_85 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_8_97 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_9_101 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_9_110 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_9_113 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_9_122 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_9_128 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_9_136 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_9_147 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_9_156 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_9_163 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_9_167 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_9_169 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_9_185 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_9_192 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_9_199 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_9_206 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_9_213 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_9_22 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_9_220 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_9_225 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_9_231 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_9_245 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_9_253 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_9_274 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_9_281 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_9_286 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_9_293 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_9_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_9_34 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_9_46 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_9_54 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_9_57 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_9_65 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_9_70 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_9_79 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_9_93 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_0 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_1 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_10 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_100 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_101 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_102 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_103 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_104 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_105 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_106 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_107 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_108 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_109 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_11 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_110 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_111 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_112 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_113 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_114 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_115 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_12 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_13 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_14 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_15 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_16 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_17 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_18 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_19 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_2 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_20 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_21 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_22 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_23 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_24 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_25 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_26 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_27 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_28 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_29 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_30 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_31 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_32 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_33 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_34 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_35 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_36 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_37 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_38 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_39 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_4 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_40 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_41 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_42 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_43 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_44 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_45 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_46 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_47 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_48 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_49 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_5 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_50 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_51 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_52 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_53 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_54 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_55 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_56 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_57 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_58 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_59 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_6 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_60 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_61 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_62 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_63 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_64 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_65 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_66 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_67 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_68 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_69 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_7 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_70 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_71 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_72 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_73 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_74 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_75 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_76 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_77 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_78 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_79 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_8 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_80 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_81 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_82 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_83 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_84 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_85 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_86 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_87 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_88 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_89 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_9 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_90 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_91 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_92 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_93 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_94 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_95 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_96 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_97 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_98 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_99 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_116 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_117 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_118 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_119 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_120 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_121 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_122 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_123 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_124 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_125 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_126 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_127 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_128 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_129 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_130 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_131 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_132 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_133 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_134 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_135 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_136 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_137 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_138 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_139 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_140 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_141 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_142 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_143 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_144 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_145 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_146 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_147 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_148 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_149 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_150 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_151 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_152 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_153 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_154 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_155 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_156 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_157 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_158 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_159 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_160 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_161 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_162 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_163 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_164 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_165 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_166 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_167 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_168 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_169 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_170 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_171 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_172 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_173 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_174 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_175 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_176 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_177 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_178 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_179 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_180 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_181 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_182 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_183 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_184 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_185 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_186 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_187 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_188 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_189 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_190 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_191 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_192 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_193 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_194 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_195 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_196 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_197 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_198 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_199 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_200 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_201 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_202 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_203 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_204 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_205 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_206 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_207 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_208 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_209 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_210 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_211 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_212 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_213 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_214 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_215 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_216 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_217 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_218 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_219 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_220 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_221 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_222 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_223 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_224 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_225 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_226 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_227 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_228 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_229 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_230 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_231 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_232 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_233 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_234 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_235 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_236 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_237 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_238 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_239 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_240 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_241 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_242 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_243 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_244 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_245 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_246 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_247 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_248 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_249 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_250 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_251 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_252 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_253 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_254 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_255 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_256 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_257 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_258 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_259 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_260 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_261 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_262 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_263 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_264 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_265 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_266 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_267 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_268 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_269 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_270 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_271 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_272 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_273 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_274 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_275 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_276 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_277 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_278 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_279 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_280 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_281 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_282 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_283 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_284 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_285 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_286 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_287 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_288 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_289 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_290 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_291 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_292 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_293 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_294 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_295 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_296 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_297 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_298 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_299 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_300 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_301 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_302 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_303 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_304 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_305 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_306 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_307 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_308 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_309 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_310 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_311 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_312 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_313 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_314 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_315 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_316 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_317 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_318 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_319 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_320 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_321 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_322 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_323 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_324 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_325 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_326 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_327 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_328 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_329 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_330 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_331 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_332 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_333 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_334 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_335 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_336 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_337 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_338 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_339 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_340 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_341 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_342 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_343 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_344 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_345 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_346 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_347 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_348 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_349 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_350 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_351 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_352 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_353 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_354 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_355 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_356 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_357 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_358 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_359 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_360 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_361 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_362 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_363 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_364 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_365 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_366 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_367 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_368 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_369 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_370 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_371 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_372 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_373 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_374 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_375 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_376 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_377 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_378 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_379 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_380 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_381 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_382 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_383 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_384 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_385 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_386 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_387 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_388 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_389 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_390 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_391 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_392 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_393 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_394 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_395 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_396 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_397 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_398 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_399 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_400 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_401 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_402 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_403 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_404 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_405 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_406 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_407 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_408 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_409 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_410 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_411 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_412 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_413 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_414 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_415 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_1 _252_ (.A(\l_fifo.genblk1[46].entry.empty ),
    .B(net29),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_089_));
 sky130_fd_sc_hd__clkbuf_1 _253_ (.A(_089_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.ready ));
 sky130_fd_sc_hd__or2_1 _254_ (.A(net1),
    .B(net2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_090_));
 sky130_fd_sc_hd__clkbuf_1 _255_ (.A(_090_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(reset_n_in));
 sky130_fd_sc_hd__and4b_1 _256_ (.A_N(\l_fifo.genblk1[47].entry.write_in ),
    .B(\l_fifo.genblk1[47].entry.empty ),
    .C(\l_fifo.genblk1[46].entry.empty ),
    .D(\l_fifo.genblk1[45].entry.empty ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_091_));
 sky130_fd_sc_hd__and4_1 _257_ (.A(\l_fifo.genblk1[44].entry.empty ),
    .B(\l_fifo.genblk1[43].entry.empty ),
    .C(\l_fifo.genblk1[42].entry.empty ),
    .D(_091_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_092_));
 sky130_fd_sc_hd__and4_1 _258_ (.A(\l_fifo.genblk1[41].entry.empty ),
    .B(\l_fifo.genblk1[40].entry.empty ),
    .C(\l_fifo.genblk1[39].entry.empty ),
    .D(_092_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_093_));
 sky130_fd_sc_hd__and4_1 _259_ (.A(\l_fifo.genblk1[38].entry.empty ),
    .B(\l_fifo.genblk1[37].entry.empty ),
    .C(\l_fifo.genblk1[36].entry.empty ),
    .D(_093_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_094_));
 sky130_fd_sc_hd__and4_1 _260_ (.A(\l_fifo.genblk1[35].entry.empty ),
    .B(\l_fifo.genblk1[34].entry.empty ),
    .C(\l_fifo.genblk1[33].entry.empty ),
    .D(_094_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_095_));
 sky130_fd_sc_hd__and4_1 _261_ (.A(\l_fifo.genblk1[32].entry.empty ),
    .B(\l_fifo.genblk1[31].entry.empty ),
    .C(\l_fifo.genblk1[30].entry.empty ),
    .D(_095_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_096_));
 sky130_fd_sc_hd__and4_1 _262_ (.A(\l_fifo.genblk1[29].entry.empty ),
    .B(\l_fifo.genblk1[28].entry.empty ),
    .C(\l_fifo.genblk1[27].entry.empty ),
    .D(_096_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_097_));
 sky130_fd_sc_hd__and4_1 _263_ (.A(\l_fifo.genblk1[26].entry.empty ),
    .B(\l_fifo.genblk1[25].entry.empty ),
    .C(\l_fifo.genblk1[24].entry.empty ),
    .D(_097_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_098_));
 sky130_fd_sc_hd__and4_1 _264_ (.A(\l_fifo.genblk1[23].entry.empty ),
    .B(\l_fifo.genblk1[22].entry.empty ),
    .C(\l_fifo.genblk1[21].entry.empty ),
    .D(_098_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_099_));
 sky130_fd_sc_hd__and4_1 _265_ (.A(\l_fifo.genblk1[20].entry.empty ),
    .B(\l_fifo.genblk1[19].entry.empty ),
    .C(\l_fifo.genblk1[18].entry.empty ),
    .D(_099_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_100_));
 sky130_fd_sc_hd__and4_1 _266_ (.A(\l_fifo.genblk1[17].entry.empty ),
    .B(\l_fifo.genblk1[16].entry.empty ),
    .C(\l_fifo.genblk1[15].entry.empty ),
    .D(_100_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_101_));
 sky130_fd_sc_hd__inv_2 _267_ (.A(net9),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_102_));
 sky130_fd_sc_hd__clkbuf_4 _268_ (.A(_102_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_103_));
 sky130_fd_sc_hd__a311o_1 _269_ (.A1(\l_fifo.genblk1[14].entry.empty ),
    .A2(\l_fifo.genblk1[13].entry.empty ),
    .A3(_101_),
    .B1(_103_),
    .C1(\l_fifo.genblk1[12].entry.empty ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_000_));
 sky130_fd_sc_hd__buf_2 _270_ (.A(_102_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_104_));
 sky130_fd_sc_hd__and4_1 _271_ (.A(\l_fifo.genblk1[14].entry.empty ),
    .B(\l_fifo.genblk1[13].entry.empty ),
    .C(\l_fifo.genblk1[12].entry.empty ),
    .D(_101_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_105_));
 sky130_fd_sc_hd__or3_1 _272_ (.A(\l_fifo.genblk1[11].entry.empty ),
    .B(_104_),
    .C(_105_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_106_));
 sky130_fd_sc_hd__clkbuf_1 _273_ (.A(_106_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_001_));
 sky130_fd_sc_hd__clkbuf_4 _274_ (.A(_104_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_107_));
 sky130_fd_sc_hd__a211o_1 _275_ (.A1(\l_fifo.genblk1[11].entry.empty ),
    .A2(_105_),
    .B1(_107_),
    .C1(\l_fifo.genblk1[10].entry.empty ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_002_));
 sky130_fd_sc_hd__a311o_1 _276_ (.A1(\l_fifo.genblk1[11].entry.empty ),
    .A2(\l_fifo.genblk1[10].entry.empty ),
    .A3(_105_),
    .B1(_103_),
    .C1(\l_fifo.genblk1[10].entry.next_is_empty ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_003_));
 sky130_fd_sc_hd__and4_1 _277_ (.A(\l_fifo.genblk1[11].entry.empty ),
    .B(\l_fifo.genblk1[10].entry.empty ),
    .C(\l_fifo.genblk1[10].entry.next_is_empty ),
    .D(_105_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_108_));
 sky130_fd_sc_hd__and4_1 _278_ (.A(\l_fifo.genblk1[8].entry.empty ),
    .B(\l_fifo.genblk1[7].entry.empty ),
    .C(\l_fifo.genblk1[6].entry.empty ),
    .D(_108_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_109_));
 sky130_fd_sc_hd__and4_1 _279_ (.A(\l_fifo.genblk1[5].entry.empty ),
    .B(\l_fifo.genblk1[4].entry.empty ),
    .C(\l_fifo.genblk1[3].entry.empty ),
    .D(_109_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_110_));
 sky130_fd_sc_hd__and3_1 _280_ (.A(\l_fifo.genblk1[2].entry.empty ),
    .B(\l_fifo.genblk1[1].entry.empty ),
    .C(_110_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_111_));
 sky130_fd_sc_hd__buf_2 _281_ (.A(net12),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_112_));
 sky130_fd_sc_hd__clkinv_2 _282_ (.A(\f_fifo.write_addr[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_113_));
 sky130_fd_sc_hd__and2_1 _283_ (.A(_113_),
    .B(\f_fifo.read_addr[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_114_));
 sky130_fd_sc_hd__nor2_1 _284_ (.A(_113_),
    .B(\f_fifo.read_addr[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_115_));
 sky130_fd_sc_hd__xnor2_1 _285_ (.A(\f_fifo.write_addr[1] ),
    .B(\f_fifo.read_addr[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_116_));
 sky130_fd_sc_hd__and4bb_1 _286_ (.A_N(_114_),
    .B_N(_115_),
    .C(\f_fifo.empty_n ),
    .D(_116_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_117_));
 sky130_fd_sc_hd__nand2_1 _287_ (.A(_112_),
    .B(_117_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_118_));
 sky130_fd_sc_hd__a21o_1 _288_ (.A1(\l_fifo.genblk1[0].entry.empty ),
    .A2(_111_),
    .B1(_118_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_004_));
 sky130_fd_sc_hd__a211o_1 _289_ (.A1(\l_fifo.genblk1[8].entry.empty ),
    .A2(_108_),
    .B1(_107_),
    .C1(\l_fifo.genblk1[7].entry.empty ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_005_));
 sky130_fd_sc_hd__a311o_1 _290_ (.A1(\l_fifo.genblk1[8].entry.empty ),
    .A2(\l_fifo.genblk1[7].entry.empty ),
    .A3(_108_),
    .B1(_103_),
    .C1(\l_fifo.genblk1[6].entry.empty ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_006_));
 sky130_fd_sc_hd__or3_1 _291_ (.A(\l_fifo.genblk1[5].entry.empty ),
    .B(_104_),
    .C(_109_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_119_));
 sky130_fd_sc_hd__clkbuf_1 _292_ (.A(_119_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_007_));
 sky130_fd_sc_hd__a211o_1 _293_ (.A1(\l_fifo.genblk1[5].entry.empty ),
    .A2(_109_),
    .B1(_107_),
    .C1(\l_fifo.genblk1[4].entry.empty ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_008_));
 sky130_fd_sc_hd__clkbuf_4 _294_ (.A(_102_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_120_));
 sky130_fd_sc_hd__a311o_1 _295_ (.A1(\l_fifo.genblk1[5].entry.empty ),
    .A2(\l_fifo.genblk1[4].entry.empty ),
    .A3(_109_),
    .B1(_120_),
    .C1(\l_fifo.genblk1[3].entry.empty ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_009_));
 sky130_fd_sc_hd__and2b_1 _296_ (.A_N(\l_fifo.genblk1[47].entry.write_in ),
    .B(\l_fifo.genblk1[47].entry.empty ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_121_));
 sky130_fd_sc_hd__or3_1 _297_ (.A(\l_fifo.genblk1[46].entry.empty ),
    .B(_104_),
    .C(_121_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_122_));
 sky130_fd_sc_hd__clkbuf_1 _298_ (.A(_122_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_010_));
 sky130_fd_sc_hd__or3_1 _299_ (.A(\l_fifo.genblk1[38].entry.empty ),
    .B(_104_),
    .C(_093_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_123_));
 sky130_fd_sc_hd__clkbuf_1 _300_ (.A(_123_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_011_));
 sky130_fd_sc_hd__a211o_1 _301_ (.A1(\l_fifo.genblk1[29].entry.empty ),
    .A2(_096_),
    .B1(_107_),
    .C1(\l_fifo.genblk1[28].entry.empty ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_012_));
 sky130_fd_sc_hd__a311o_1 _302_ (.A1(\l_fifo.genblk1[20].entry.empty ),
    .A2(\l_fifo.genblk1[19].entry.empty ),
    .A3(_099_),
    .B1(_120_),
    .C1(\l_fifo.genblk1[18].entry.empty ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_013_));
 sky130_fd_sc_hd__and2_1 _303_ (.A(net1),
    .B(net2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_124_));
 sky130_fd_sc_hd__clkbuf_1 _304_ (.A(_124_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_014_));
 sky130_fd_sc_hd__and2_1 _305_ (.A(net3),
    .B(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_125_));
 sky130_fd_sc_hd__clkbuf_1 _306_ (.A(_125_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_015_));
 sky130_fd_sc_hd__and2_1 _307_ (.A(net1),
    .B(net4),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_126_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _308_ (.A(_126_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_016_));
 sky130_fd_sc_hd__and2_1 _309_ (.A(net1),
    .B(net5),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_127_));
 sky130_fd_sc_hd__clkbuf_1 _310_ (.A(_127_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_017_));
 sky130_fd_sc_hd__and2_1 _311_ (.A(net1),
    .B(net6),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_128_));
 sky130_fd_sc_hd__clkbuf_1 _312_ (.A(_128_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_018_));
 sky130_fd_sc_hd__and2_1 _313_ (.A(net1),
    .B(net7),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_129_));
 sky130_fd_sc_hd__clkbuf_1 _314_ (.A(_129_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_019_));
 sky130_fd_sc_hd__inv_2 _315_ (.A(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_130_));
 sky130_fd_sc_hd__and3_1 _316_ (.A(\f_fifo.empty_n ),
    .B(net3),
    .C(_130_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_131_));
 sky130_fd_sc_hd__and2_1 _317_ (.A(\f_fifo.read_addr[0] ),
    .B(_131_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_132_));
 sky130_fd_sc_hd__o21ai_1 _318_ (.A1(\f_fifo.read_addr[0] ),
    .A2(_131_),
    .B1(_112_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_133_));
 sky130_fd_sc_hd__nor2_1 _319_ (.A(_132_),
    .B(_133_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_020_));
 sky130_fd_sc_hd__a31o_1 _320_ (.A1(\f_fifo.read_addr[1] ),
    .A2(\f_fifo.read_addr[0] ),
    .A3(_131_),
    .B1(_104_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_134_));
 sky130_fd_sc_hd__o21ba_1 _321_ (.A1(\f_fifo.read_addr[1] ),
    .A2(_132_),
    .B1_N(_134_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_021_));
 sky130_fd_sc_hd__a41o_1 _322_ (.A1(\l_fifo.genblk1[2].entry.empty ),
    .A2(\l_fifo.genblk1[1].entry.empty ),
    .A3(\l_fifo.genblk1[0].entry.empty ),
    .A4(_110_),
    .B1(_117_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_135_));
 sky130_fd_sc_hd__clkbuf_4 _323_ (.A(_135_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_136_));
 sky130_fd_sc_hd__o21ai_1 _324_ (.A1(_113_),
    .A2(_136_),
    .B1(_112_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_137_));
 sky130_fd_sc_hd__a21oi_1 _325_ (.A1(_113_),
    .A2(_136_),
    .B1(_137_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_022_));
 sky130_fd_sc_hd__nor2_2 _326_ (.A(\f_fifo.write_addr[1] ),
    .B(\f_fifo.write_addr[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_138_));
 sky130_fd_sc_hd__and2_2 _327_ (.A(\f_fifo.write_addr[1] ),
    .B(\f_fifo.write_addr[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_139_));
 sky130_fd_sc_hd__nor2_1 _328_ (.A(_138_),
    .B(_139_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_140_));
 sky130_fd_sc_hd__mux2_1 _329_ (.A0(_140_),
    .A1(\f_fifo.write_addr[1] ),
    .S(_136_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_141_));
 sky130_fd_sc_hd__and2_1 _330_ (.A(_112_),
    .B(_141_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_142_));
 sky130_fd_sc_hd__clkbuf_1 _331_ (.A(_142_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_023_));
 sky130_fd_sc_hd__mux2_1 _332_ (.A0(_114_),
    .A1(_115_),
    .S(_116_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_143_));
 sky130_fd_sc_hd__nand2_2 _333_ (.A(_131_),
    .B(_143_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_144_));
 sky130_fd_sc_hd__nand2_1 _334_ (.A(\f_fifo.empty_n ),
    .B(_144_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_145_));
 sky130_fd_sc_hd__a21oi_1 _335_ (.A1(_136_),
    .A2(_145_),
    .B1(_107_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_024_));
 sky130_fd_sc_hd__clkbuf_2 _336_ (.A(net8),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_146_));
 sky130_fd_sc_hd__a21bo_2 _337_ (.A1(_135_),
    .A2(_144_),
    .B1_N(_138_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_147_));
 sky130_fd_sc_hd__inv_2 _338_ (.A(\f_fifo.data_in[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_148_));
 sky130_fd_sc_hd__nor2_1 _339_ (.A(_148_),
    .B(_136_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_149_));
 sky130_fd_sc_hd__a22o_1 _340_ (.A1(\f_fifo.fifo_data[0][0] ),
    .A2(_147_),
    .B1(_149_),
    .B2(_138_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_150_));
 sky130_fd_sc_hd__and2_1 _341_ (.A(_146_),
    .B(_150_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_151_));
 sky130_fd_sc_hd__clkbuf_1 _342_ (.A(_151_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_025_));
 sky130_fd_sc_hd__inv_2 _343_ (.A(\f_fifo.data_in[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_152_));
 sky130_fd_sc_hd__nor2_2 _344_ (.A(_152_),
    .B(_136_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_153_));
 sky130_fd_sc_hd__a22o_1 _345_ (.A1(\f_fifo.fifo_data[0][1] ),
    .A2(_147_),
    .B1(_153_),
    .B2(_138_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_154_));
 sky130_fd_sc_hd__and2_1 _346_ (.A(_146_),
    .B(_154_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_155_));
 sky130_fd_sc_hd__clkbuf_1 _347_ (.A(_155_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_026_));
 sky130_fd_sc_hd__inv_2 _348_ (.A(\f_fifo.data_in[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_156_));
 sky130_fd_sc_hd__nor2_2 _349_ (.A(_156_),
    .B(_136_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_157_));
 sky130_fd_sc_hd__a22o_1 _350_ (.A1(\f_fifo.fifo_data[0][2] ),
    .A2(_147_),
    .B1(_157_),
    .B2(_138_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_158_));
 sky130_fd_sc_hd__and2_1 _351_ (.A(_146_),
    .B(_158_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_159_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _352_ (.A(_159_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_027_));
 sky130_fd_sc_hd__inv_2 _353_ (.A(\f_fifo.data_in[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_160_));
 sky130_fd_sc_hd__nor2_2 _354_ (.A(_160_),
    .B(_136_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_161_));
 sky130_fd_sc_hd__a22o_1 _355_ (.A1(\f_fifo.fifo_data[0][3] ),
    .A2(_147_),
    .B1(_161_),
    .B2(_138_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_162_));
 sky130_fd_sc_hd__and2_1 _356_ (.A(_146_),
    .B(_162_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_163_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _357_ (.A(_163_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_028_));
 sky130_fd_sc_hd__inv_2 _358_ (.A(\f_fifo.data_in[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_164_));
 sky130_fd_sc_hd__nor2_2 _359_ (.A(_164_),
    .B(_136_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_165_));
 sky130_fd_sc_hd__a22o_1 _360_ (.A1(\f_fifo.fifo_data[0][4] ),
    .A2(_147_),
    .B1(_165_),
    .B2(_138_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_166_));
 sky130_fd_sc_hd__and2_1 _361_ (.A(_146_),
    .B(_166_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_167_));
 sky130_fd_sc_hd__clkbuf_1 _362_ (.A(_167_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_029_));
 sky130_fd_sc_hd__inv_2 _363_ (.A(\f_fifo.data_in[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_168_));
 sky130_fd_sc_hd__nor2_2 _364_ (.A(_168_),
    .B(_136_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_169_));
 sky130_fd_sc_hd__a22o_1 _365_ (.A1(\f_fifo.fifo_data[0][5] ),
    .A2(_147_),
    .B1(_169_),
    .B2(_138_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_170_));
 sky130_fd_sc_hd__and2_1 _366_ (.A(_146_),
    .B(_170_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_171_));
 sky130_fd_sc_hd__clkbuf_1 _367_ (.A(_171_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_030_));
 sky130_fd_sc_hd__nor2_2 _368_ (.A(\f_fifo.write_addr[1] ),
    .B(_113_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_172_));
 sky130_fd_sc_hd__a21bo_2 _369_ (.A1(_135_),
    .A2(_144_),
    .B1_N(_172_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_173_));
 sky130_fd_sc_hd__a22o_1 _370_ (.A1(_149_),
    .A2(_172_),
    .B1(_173_),
    .B2(\f_fifo.fifo_data[1][0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_174_));
 sky130_fd_sc_hd__and2_1 _371_ (.A(_146_),
    .B(_174_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_175_));
 sky130_fd_sc_hd__clkbuf_1 _372_ (.A(_175_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_031_));
 sky130_fd_sc_hd__a22o_1 _373_ (.A1(_153_),
    .A2(_172_),
    .B1(_173_),
    .B2(\f_fifo.fifo_data[1][1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_176_));
 sky130_fd_sc_hd__and2_1 _374_ (.A(_146_),
    .B(_176_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_177_));
 sky130_fd_sc_hd__clkbuf_1 _375_ (.A(_177_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_032_));
 sky130_fd_sc_hd__a22o_1 _376_ (.A1(_157_),
    .A2(_172_),
    .B1(_173_),
    .B2(\f_fifo.fifo_data[1][2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_178_));
 sky130_fd_sc_hd__and2_1 _377_ (.A(_146_),
    .B(_178_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_179_));
 sky130_fd_sc_hd__clkbuf_1 _378_ (.A(_179_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_033_));
 sky130_fd_sc_hd__a22o_1 _379_ (.A1(_161_),
    .A2(_172_),
    .B1(_173_),
    .B2(\f_fifo.fifo_data[1][3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_180_));
 sky130_fd_sc_hd__and2_1 _380_ (.A(_146_),
    .B(_180_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_181_));
 sky130_fd_sc_hd__clkbuf_1 _381_ (.A(_181_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_034_));
 sky130_fd_sc_hd__clkbuf_2 _382_ (.A(net8),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_182_));
 sky130_fd_sc_hd__a22o_1 _383_ (.A1(_165_),
    .A2(_172_),
    .B1(_173_),
    .B2(\f_fifo.fifo_data[1][4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_183_));
 sky130_fd_sc_hd__and2_1 _384_ (.A(_182_),
    .B(_183_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_184_));
 sky130_fd_sc_hd__clkbuf_1 _385_ (.A(_184_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_035_));
 sky130_fd_sc_hd__a22o_1 _386_ (.A1(_169_),
    .A2(_172_),
    .B1(_173_),
    .B2(\f_fifo.fifo_data[1][5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_185_));
 sky130_fd_sc_hd__and2_1 _387_ (.A(_182_),
    .B(_185_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_186_));
 sky130_fd_sc_hd__clkbuf_1 _388_ (.A(_186_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_036_));
 sky130_fd_sc_hd__and2_2 _389_ (.A(\f_fifo.write_addr[1] ),
    .B(_113_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_187_));
 sky130_fd_sc_hd__a21bo_1 _390_ (.A1(_135_),
    .A2(_144_),
    .B1_N(_187_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_188_));
 sky130_fd_sc_hd__a22o_1 _391_ (.A1(_149_),
    .A2(_187_),
    .B1(_188_),
    .B2(\f_fifo.fifo_data[2][0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_189_));
 sky130_fd_sc_hd__and2_1 _392_ (.A(_182_),
    .B(_189_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_190_));
 sky130_fd_sc_hd__clkbuf_1 _393_ (.A(_190_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_037_));
 sky130_fd_sc_hd__a22o_1 _394_ (.A1(_153_),
    .A2(_187_),
    .B1(_188_),
    .B2(\f_fifo.fifo_data[2][1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_191_));
 sky130_fd_sc_hd__and2_1 _395_ (.A(_182_),
    .B(_191_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_192_));
 sky130_fd_sc_hd__clkbuf_1 _396_ (.A(_192_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_038_));
 sky130_fd_sc_hd__a22o_1 _397_ (.A1(_157_),
    .A2(_187_),
    .B1(_188_),
    .B2(\f_fifo.fifo_data[2][2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_193_));
 sky130_fd_sc_hd__and2_1 _398_ (.A(_182_),
    .B(_193_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_194_));
 sky130_fd_sc_hd__clkbuf_1 _399_ (.A(_194_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_039_));
 sky130_fd_sc_hd__a22o_1 _400_ (.A1(_161_),
    .A2(_187_),
    .B1(_188_),
    .B2(\f_fifo.fifo_data[2][3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_195_));
 sky130_fd_sc_hd__and2_1 _401_ (.A(_182_),
    .B(_195_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_196_));
 sky130_fd_sc_hd__clkbuf_1 _402_ (.A(_196_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_040_));
 sky130_fd_sc_hd__a22o_1 _403_ (.A1(_165_),
    .A2(_187_),
    .B1(_188_),
    .B2(\f_fifo.fifo_data[2][4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_197_));
 sky130_fd_sc_hd__and2_1 _404_ (.A(_182_),
    .B(_197_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_198_));
 sky130_fd_sc_hd__clkbuf_1 _405_ (.A(_198_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_041_));
 sky130_fd_sc_hd__a22o_1 _406_ (.A1(_169_),
    .A2(_187_),
    .B1(_188_),
    .B2(\f_fifo.fifo_data[2][5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_199_));
 sky130_fd_sc_hd__and2_1 _407_ (.A(_182_),
    .B(_199_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_200_));
 sky130_fd_sc_hd__clkbuf_1 _408_ (.A(_200_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_042_));
 sky130_fd_sc_hd__a21bo_2 _409_ (.A1(_135_),
    .A2(_144_),
    .B1_N(_139_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_201_));
 sky130_fd_sc_hd__a22o_1 _410_ (.A1(_139_),
    .A2(_149_),
    .B1(_201_),
    .B2(\f_fifo.fifo_data[3][0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_202_));
 sky130_fd_sc_hd__and2_1 _411_ (.A(_182_),
    .B(_202_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_203_));
 sky130_fd_sc_hd__clkbuf_1 _412_ (.A(_203_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_043_));
 sky130_fd_sc_hd__a22o_1 _413_ (.A1(_139_),
    .A2(_153_),
    .B1(_201_),
    .B2(\f_fifo.fifo_data[3][1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_204_));
 sky130_fd_sc_hd__and2_1 _414_ (.A(_182_),
    .B(_204_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_205_));
 sky130_fd_sc_hd__clkbuf_1 _415_ (.A(_205_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_044_));
 sky130_fd_sc_hd__a22o_1 _416_ (.A1(_139_),
    .A2(_157_),
    .B1(_201_),
    .B2(\f_fifo.fifo_data[3][2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_206_));
 sky130_fd_sc_hd__and2_1 _417_ (.A(net9),
    .B(_206_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_207_));
 sky130_fd_sc_hd__clkbuf_1 _418_ (.A(_207_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_045_));
 sky130_fd_sc_hd__a22o_1 _419_ (.A1(_139_),
    .A2(_161_),
    .B1(_201_),
    .B2(\f_fifo.fifo_data[3][3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_208_));
 sky130_fd_sc_hd__and2_1 _420_ (.A(net8),
    .B(_208_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_209_));
 sky130_fd_sc_hd__clkbuf_1 _421_ (.A(_209_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_046_));
 sky130_fd_sc_hd__a22o_1 _422_ (.A1(_139_),
    .A2(_165_),
    .B1(_201_),
    .B2(\f_fifo.fifo_data[3][4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_210_));
 sky130_fd_sc_hd__and2_1 _423_ (.A(net8),
    .B(_210_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_211_));
 sky130_fd_sc_hd__clkbuf_1 _424_ (.A(_211_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_047_));
 sky130_fd_sc_hd__a22o_1 _425_ (.A1(_139_),
    .A2(_169_),
    .B1(_201_),
    .B2(\f_fifo.fifo_data[3][5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_212_));
 sky130_fd_sc_hd__and2_1 _426_ (.A(net8),
    .B(_212_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_213_));
 sky130_fd_sc_hd__clkbuf_1 _427_ (.A(_213_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_048_));
 sky130_fd_sc_hd__and2_1 _428_ (.A(_130_),
    .B(net5),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_214_));
 sky130_fd_sc_hd__xnor2_2 _429_ (.A(\f_fifo.read_addr[1] ),
    .B(_214_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_215_));
 sky130_fd_sc_hd__inv_2 _430_ (.A(_215_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_216_));
 sky130_fd_sc_hd__a21oi_1 _431_ (.A1(_130_),
    .A2(net4),
    .B1(\f_fifo.read_addr[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_217_));
 sky130_fd_sc_hd__and3_1 _432_ (.A(\f_fifo.read_addr[0] ),
    .B(_130_),
    .C(net4),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_218_));
 sky130_fd_sc_hd__or2_1 _433_ (.A(_215_),
    .B(_218_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_219_));
 sky130_fd_sc_hd__o21ai_2 _434_ (.A1(_216_),
    .A2(_217_),
    .B1(_219_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_220_));
 sky130_fd_sc_hd__or2_1 _435_ (.A(_217_),
    .B(_218_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_221_));
 sky130_fd_sc_hd__buf_2 _436_ (.A(_221_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_222_));
 sky130_fd_sc_hd__o21a_1 _437_ (.A1(_216_),
    .A2(_217_),
    .B1(_219_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_223_));
 sky130_fd_sc_hd__a21o_1 _438_ (.A1(\f_fifo.fifo_data[2][0] ),
    .A2(_222_),
    .B1(_223_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_224_));
 sky130_fd_sc_hd__nor2_2 _439_ (.A(_215_),
    .B(_222_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_225_));
 sky130_fd_sc_hd__nor2_2 _440_ (.A(_216_),
    .B(_222_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_226_));
 sky130_fd_sc_hd__a22o_1 _441_ (.A1(\f_fifo.fifo_data[3][0] ),
    .A2(_225_),
    .B1(_226_),
    .B2(\f_fifo.fifo_data[1][0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_227_));
 sky130_fd_sc_hd__o221a_1 _442_ (.A1(\f_fifo.fifo_data[0][0] ),
    .A2(_220_),
    .B1(_224_),
    .B2(_227_),
    .C1(_112_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_049_));
 sky130_fd_sc_hd__a22o_1 _443_ (.A1(\f_fifo.fifo_data[3][1] ),
    .A2(_225_),
    .B1(_226_),
    .B2(\f_fifo.fifo_data[1][1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_228_));
 sky130_fd_sc_hd__a21o_1 _444_ (.A1(\f_fifo.fifo_data[2][1] ),
    .A2(_222_),
    .B1(_223_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_229_));
 sky130_fd_sc_hd__o221a_1 _445_ (.A1(\f_fifo.fifo_data[0][1] ),
    .A2(_220_),
    .B1(_228_),
    .B2(_229_),
    .C1(_112_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_050_));
 sky130_fd_sc_hd__a22o_1 _446_ (.A1(\f_fifo.fifo_data[3][2] ),
    .A2(_225_),
    .B1(_226_),
    .B2(\f_fifo.fifo_data[1][2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_230_));
 sky130_fd_sc_hd__a21o_1 _447_ (.A1(\f_fifo.fifo_data[2][2] ),
    .A2(_222_),
    .B1(_223_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_231_));
 sky130_fd_sc_hd__o221a_1 _448_ (.A1(\f_fifo.fifo_data[0][2] ),
    .A2(_220_),
    .B1(_230_),
    .B2(_231_),
    .C1(_112_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_051_));
 sky130_fd_sc_hd__a22o_1 _449_ (.A1(\f_fifo.fifo_data[3][3] ),
    .A2(_225_),
    .B1(_226_),
    .B2(\f_fifo.fifo_data[1][3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_232_));
 sky130_fd_sc_hd__a21o_1 _450_ (.A1(\f_fifo.fifo_data[2][3] ),
    .A2(_222_),
    .B1(_223_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_233_));
 sky130_fd_sc_hd__o221a_1 _451_ (.A1(\f_fifo.fifo_data[0][3] ),
    .A2(_220_),
    .B1(_232_),
    .B2(_233_),
    .C1(_112_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_052_));
 sky130_fd_sc_hd__a22o_1 _452_ (.A1(\f_fifo.fifo_data[3][4] ),
    .A2(_225_),
    .B1(_226_),
    .B2(\f_fifo.fifo_data[1][4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_234_));
 sky130_fd_sc_hd__a21o_1 _453_ (.A1(\f_fifo.fifo_data[2][4] ),
    .A2(_222_),
    .B1(_223_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_235_));
 sky130_fd_sc_hd__o221a_1 _454_ (.A1(\f_fifo.fifo_data[0][4] ),
    .A2(_220_),
    .B1(_234_),
    .B2(_235_),
    .C1(_112_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_053_));
 sky130_fd_sc_hd__a221o_1 _455_ (.A1(\f_fifo.fifo_data[2][5] ),
    .A2(_222_),
    .B1(_225_),
    .B2(\f_fifo.fifo_data[3][5] ),
    .C1(_223_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_236_));
 sky130_fd_sc_hd__a21o_1 _456_ (.A1(\f_fifo.fifo_data[1][5] ),
    .A2(_226_),
    .B1(_236_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_237_));
 sky130_fd_sc_hd__o211a_1 _457_ (.A1(\f_fifo.fifo_data[0][5] ),
    .A2(_220_),
    .B1(_237_),
    .C1(_112_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_054_));
 sky130_fd_sc_hd__or3_1 _458_ (.A(\l_fifo.genblk1[8].entry.empty ),
    .B(_104_),
    .C(_108_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_238_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _459_ (.A(_238_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_055_));
 sky130_fd_sc_hd__a211o_1 _460_ (.A1(\l_fifo.genblk1[46].entry.empty ),
    .A2(_121_),
    .B1(_107_),
    .C1(\l_fifo.genblk1[45].entry.empty ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_056_));
 sky130_fd_sc_hd__or3_1 _461_ (.A(\l_fifo.genblk1[44].entry.empty ),
    .B(_104_),
    .C(_091_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_239_));
 sky130_fd_sc_hd__clkbuf_1 _462_ (.A(_239_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_057_));
 sky130_fd_sc_hd__a211o_1 _463_ (.A1(\l_fifo.genblk1[44].entry.empty ),
    .A2(_091_),
    .B1(_107_),
    .C1(\l_fifo.genblk1[43].entry.empty ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_058_));
 sky130_fd_sc_hd__a311o_1 _464_ (.A1(\l_fifo.genblk1[44].entry.empty ),
    .A2(\l_fifo.genblk1[43].entry.empty ),
    .A3(_091_),
    .B1(_120_),
    .C1(\l_fifo.genblk1[42].entry.empty ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_059_));
 sky130_fd_sc_hd__or3_1 _465_ (.A(\l_fifo.genblk1[41].entry.empty ),
    .B(_104_),
    .C(_092_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_240_));
 sky130_fd_sc_hd__clkbuf_1 _466_ (.A(_240_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_060_));
 sky130_fd_sc_hd__a211o_1 _467_ (.A1(\l_fifo.genblk1[41].entry.empty ),
    .A2(_092_),
    .B1(_107_),
    .C1(\l_fifo.genblk1[40].entry.empty ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_061_));
 sky130_fd_sc_hd__a311o_1 _468_ (.A1(\l_fifo.genblk1[41].entry.empty ),
    .A2(\l_fifo.genblk1[40].entry.empty ),
    .A3(_092_),
    .B1(_120_),
    .C1(\l_fifo.genblk1[39].entry.empty ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_062_));
 sky130_fd_sc_hd__buf_2 _469_ (.A(_102_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_241_));
 sky130_fd_sc_hd__or3_1 _470_ (.A(\l_fifo.genblk1[2].entry.empty ),
    .B(_241_),
    .C(_110_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_242_));
 sky130_fd_sc_hd__clkbuf_1 _471_ (.A(_242_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_063_));
 sky130_fd_sc_hd__a211o_1 _472_ (.A1(\l_fifo.genblk1[38].entry.empty ),
    .A2(_093_),
    .B1(_107_),
    .C1(\l_fifo.genblk1[37].entry.empty ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_064_));
 sky130_fd_sc_hd__a311o_1 _473_ (.A1(\l_fifo.genblk1[38].entry.empty ),
    .A2(\l_fifo.genblk1[37].entry.empty ),
    .A3(_093_),
    .B1(_120_),
    .C1(\l_fifo.genblk1[36].entry.empty ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_065_));
 sky130_fd_sc_hd__or3_1 _474_ (.A(\l_fifo.genblk1[35].entry.empty ),
    .B(_241_),
    .C(_094_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_243_));
 sky130_fd_sc_hd__clkbuf_1 _475_ (.A(_243_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_066_));
 sky130_fd_sc_hd__a211o_1 _476_ (.A1(\l_fifo.genblk1[35].entry.empty ),
    .A2(_094_),
    .B1(_107_),
    .C1(\l_fifo.genblk1[34].entry.empty ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_067_));
 sky130_fd_sc_hd__a311o_1 _477_ (.A1(\l_fifo.genblk1[35].entry.empty ),
    .A2(\l_fifo.genblk1[34].entry.empty ),
    .A3(_094_),
    .B1(_120_),
    .C1(\l_fifo.genblk1[33].entry.empty ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_068_));
 sky130_fd_sc_hd__or3_1 _478_ (.A(\l_fifo.genblk1[32].entry.empty ),
    .B(_241_),
    .C(_095_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_244_));
 sky130_fd_sc_hd__clkbuf_1 _479_ (.A(_244_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_069_));
 sky130_fd_sc_hd__a211o_1 _480_ (.A1(\l_fifo.genblk1[32].entry.empty ),
    .A2(_095_),
    .B1(_103_),
    .C1(\l_fifo.genblk1[31].entry.empty ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_070_));
 sky130_fd_sc_hd__a311o_1 _481_ (.A1(\l_fifo.genblk1[32].entry.empty ),
    .A2(\l_fifo.genblk1[31].entry.empty ),
    .A3(_095_),
    .B1(_120_),
    .C1(\l_fifo.genblk1[30].entry.empty ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_071_));
 sky130_fd_sc_hd__or3_1 _482_ (.A(\l_fifo.genblk1[29].entry.empty ),
    .B(_241_),
    .C(_096_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_245_));
 sky130_fd_sc_hd__clkbuf_1 _483_ (.A(_245_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_072_));
 sky130_fd_sc_hd__a211o_1 _484_ (.A1(\l_fifo.genblk1[2].entry.empty ),
    .A2(_110_),
    .B1(_103_),
    .C1(\l_fifo.genblk1[1].entry.empty ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_073_));
 sky130_fd_sc_hd__a311o_1 _485_ (.A1(\l_fifo.genblk1[29].entry.empty ),
    .A2(\l_fifo.genblk1[28].entry.empty ),
    .A3(_096_),
    .B1(_120_),
    .C1(\l_fifo.genblk1[27].entry.empty ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_074_));
 sky130_fd_sc_hd__or3_1 _486_ (.A(\l_fifo.genblk1[26].entry.empty ),
    .B(_241_),
    .C(_097_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_246_));
 sky130_fd_sc_hd__clkbuf_1 _487_ (.A(_246_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_075_));
 sky130_fd_sc_hd__a211o_1 _488_ (.A1(\l_fifo.genblk1[26].entry.empty ),
    .A2(_097_),
    .B1(_103_),
    .C1(\l_fifo.genblk1[25].entry.empty ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_076_));
 sky130_fd_sc_hd__a311o_1 _489_ (.A1(\l_fifo.genblk1[26].entry.empty ),
    .A2(\l_fifo.genblk1[25].entry.empty ),
    .A3(_097_),
    .B1(_120_),
    .C1(\l_fifo.genblk1[24].entry.empty ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_077_));
 sky130_fd_sc_hd__or3_1 _490_ (.A(\l_fifo.genblk1[23].entry.empty ),
    .B(_241_),
    .C(_098_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_247_));
 sky130_fd_sc_hd__clkbuf_1 _491_ (.A(_247_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_078_));
 sky130_fd_sc_hd__a211o_1 _492_ (.A1(\l_fifo.genblk1[23].entry.empty ),
    .A2(_098_),
    .B1(_103_),
    .C1(\l_fifo.genblk1[22].entry.empty ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_079_));
 sky130_fd_sc_hd__a311o_1 _493_ (.A1(\l_fifo.genblk1[23].entry.empty ),
    .A2(\l_fifo.genblk1[22].entry.empty ),
    .A3(_098_),
    .B1(_120_),
    .C1(\l_fifo.genblk1[21].entry.empty ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_080_));
 sky130_fd_sc_hd__or3_1 _494_ (.A(\l_fifo.genblk1[20].entry.empty ),
    .B(_241_),
    .C(_099_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_248_));
 sky130_fd_sc_hd__clkbuf_1 _495_ (.A(_248_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_081_));
 sky130_fd_sc_hd__a211o_1 _496_ (.A1(\l_fifo.genblk1[20].entry.empty ),
    .A2(_099_),
    .B1(_103_),
    .C1(\l_fifo.genblk1[19].entry.empty ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_082_));
 sky130_fd_sc_hd__or3_1 _497_ (.A(\l_fifo.genblk1[0].entry.empty ),
    .B(_241_),
    .C(_111_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_249_));
 sky130_fd_sc_hd__clkbuf_1 _498_ (.A(_249_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_083_));
 sky130_fd_sc_hd__or3_1 _499_ (.A(\l_fifo.genblk1[17].entry.empty ),
    .B(_241_),
    .C(_100_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_250_));
 sky130_fd_sc_hd__clkbuf_1 _500_ (.A(_250_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_084_));
 sky130_fd_sc_hd__a211o_1 _501_ (.A1(\l_fifo.genblk1[17].entry.empty ),
    .A2(_100_),
    .B1(_103_),
    .C1(\l_fifo.genblk1[16].entry.empty ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_085_));
 sky130_fd_sc_hd__a311o_1 _502_ (.A1(\l_fifo.genblk1[17].entry.empty ),
    .A2(\l_fifo.genblk1[16].entry.empty ),
    .A3(_100_),
    .B1(_104_),
    .C1(\l_fifo.genblk1[15].entry.empty ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_086_));
 sky130_fd_sc_hd__or3_1 _503_ (.A(\l_fifo.genblk1[14].entry.empty ),
    .B(_241_),
    .C(_101_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_251_));
 sky130_fd_sc_hd__clkbuf_1 _504_ (.A(_251_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_087_));
 sky130_fd_sc_hd__a211o_1 _505_ (.A1(\l_fifo.genblk1[14].entry.empty ),
    .A2(_101_),
    .B1(_103_),
    .C1(\l_fifo.genblk1[13].entry.empty ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_088_));
 sky130_fd_sc_hd__dfxtp_2 _506_ (.CLK(clknet_3_0__leaf_io_in[0]),
    .D(_000_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[13].entry.empty ));
 sky130_fd_sc_hd__dfxtp_2 _507_ (.CLK(clknet_3_0__leaf_io_in[0]),
    .D(_001_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[12].entry.empty ));
 sky130_fd_sc_hd__dfxtp_4 _508_ (.CLK(clknet_3_0__leaf_io_in[0]),
    .D(_002_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[11].entry.empty ));
 sky130_fd_sc_hd__dfxtp_2 _509_ (.CLK(clknet_3_1__leaf_io_in[0]),
    .D(_003_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[10].entry.empty ));
 sky130_fd_sc_hd__dfxtp_2 _510_ (.CLK(clknet_3_7__leaf_io_in[0]),
    .D(_004_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[0].entry.empty ));
 sky130_fd_sc_hd__dfxtp_2 _511_ (.CLK(clknet_3_1__leaf_io_in[0]),
    .D(_005_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[8].entry.empty ));
 sky130_fd_sc_hd__dfxtp_2 _512_ (.CLK(clknet_3_4__leaf_io_in[0]),
    .D(_006_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[7].entry.empty ));
 sky130_fd_sc_hd__dfxtp_2 _513_ (.CLK(clknet_3_4__leaf_io_in[0]),
    .D(_007_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[6].entry.empty ));
 sky130_fd_sc_hd__dfxtp_2 _514_ (.CLK(clknet_3_0__leaf_io_in[0]),
    .D(_008_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[5].entry.empty ));
 sky130_fd_sc_hd__dfxtp_2 _515_ (.CLK(clknet_3_7__leaf_io_in[0]),
    .D(_009_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[4].entry.empty ));
 sky130_fd_sc_hd__dfxtp_2 _516_ (.CLK(clknet_3_7__leaf_io_in[0]),
    .D(_010_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[47].entry.empty ));
 sky130_fd_sc_hd__dfxtp_2 _517_ (.CLK(clknet_3_2__leaf_io_in[0]),
    .D(_011_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[39].entry.empty ));
 sky130_fd_sc_hd__dfxtp_2 _518_ (.CLK(clknet_3_0__leaf_io_in[0]),
    .D(_012_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[29].entry.empty ));
 sky130_fd_sc_hd__dfxtp_2 _519_ (.CLK(clknet_3_1__leaf_io_in[0]),
    .D(_013_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[19].entry.empty ));
 sky130_fd_sc_hd__dfxtp_1 _520_ (.CLK(clknet_3_7__leaf_io_in[0]),
    .D(_014_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\data_in_buffer[0].A ));
 sky130_fd_sc_hd__dfxtp_1 _521_ (.CLK(clknet_3_0__leaf_io_in[0]),
    .D(_015_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\data_in_buffer[1].A ));
 sky130_fd_sc_hd__dfxtp_1 _522_ (.CLK(clknet_3_0__leaf_io_in[0]),
    .D(_016_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\data_in_buffer[2].A ));
 sky130_fd_sc_hd__dfxtp_1 _523_ (.CLK(clknet_3_5__leaf_io_in[0]),
    .D(_017_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\data_in_buffer[3].A ));
 sky130_fd_sc_hd__dfxtp_1 _524_ (.CLK(clknet_3_2__leaf_io_in[0]),
    .D(_018_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\data_in_buffer[4].A ));
 sky130_fd_sc_hd__dfxtp_1 _525_ (.CLK(clknet_3_5__leaf_io_in[0]),
    .D(_019_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\data_in_buffer[5].A ));
 sky130_fd_sc_hd__dfxtp_1 _526_ (.CLK(clknet_3_6__leaf_io_in[0]),
    .D(_020_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\f_fifo.read_addr[0] ));
 sky130_fd_sc_hd__dfxtp_2 _527_ (.CLK(clknet_3_2__leaf_io_in[0]),
    .D(_021_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\f_fifo.read_addr[1] ));
 sky130_fd_sc_hd__dfxtp_1 _528_ (.CLK(clknet_3_0__leaf_io_in[0]),
    .D(_022_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\f_fifo.write_addr[0] ));
 sky130_fd_sc_hd__dfxtp_2 _529_ (.CLK(clknet_3_7__leaf_io_in[0]),
    .D(_023_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\f_fifo.write_addr[1] ));
 sky130_fd_sc_hd__dfxtp_2 _530_ (.CLK(clknet_3_2__leaf_io_in[0]),
    .D(_024_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\f_fifo.empty_n ));
 sky130_fd_sc_hd__dfxtp_1 _531_ (.CLK(clknet_3_5__leaf_io_in[0]),
    .D(_025_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\f_fifo.fifo_data[0][0] ));
 sky130_fd_sc_hd__dfxtp_1 _532_ (.CLK(clknet_3_0__leaf_io_in[0]),
    .D(_026_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\f_fifo.fifo_data[0][1] ));
 sky130_fd_sc_hd__dfxtp_1 _533_ (.CLK(clknet_3_5__leaf_io_in[0]),
    .D(_027_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\f_fifo.fifo_data[0][2] ));
 sky130_fd_sc_hd__dfxtp_1 _534_ (.CLK(clknet_3_5__leaf_io_in[0]),
    .D(_028_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\f_fifo.fifo_data[0][3] ));
 sky130_fd_sc_hd__dfxtp_1 _535_ (.CLK(clknet_3_6__leaf_io_in[0]),
    .D(_029_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\f_fifo.fifo_data[0][4] ));
 sky130_fd_sc_hd__dfxtp_1 _536_ (.CLK(clknet_3_3__leaf_io_in[0]),
    .D(_030_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\f_fifo.fifo_data[0][5] ));
 sky130_fd_sc_hd__dfxtp_1 _537_ (.CLK(clknet_3_6__leaf_io_in[0]),
    .D(_031_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\f_fifo.fifo_data[1][0] ));
 sky130_fd_sc_hd__dfxtp_1 _538_ (.CLK(clknet_3_1__leaf_io_in[0]),
    .D(_032_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\f_fifo.fifo_data[1][1] ));
 sky130_fd_sc_hd__dfxtp_1 _539_ (.CLK(clknet_3_0__leaf_io_in[0]),
    .D(_033_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\f_fifo.fifo_data[1][2] ));
 sky130_fd_sc_hd__dfxtp_1 _540_ (.CLK(clknet_3_4__leaf_io_in[0]),
    .D(_034_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\f_fifo.fifo_data[1][3] ));
 sky130_fd_sc_hd__dfxtp_1 _541_ (.CLK(clknet_3_3__leaf_io_in[0]),
    .D(_035_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\f_fifo.fifo_data[1][4] ));
 sky130_fd_sc_hd__dfxtp_1 _542_ (.CLK(clknet_3_0__leaf_io_in[0]),
    .D(_036_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\f_fifo.fifo_data[1][5] ));
 sky130_fd_sc_hd__dfxtp_1 _543_ (.CLK(clknet_3_1__leaf_io_in[0]),
    .D(_037_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\f_fifo.fifo_data[2][0] ));
 sky130_fd_sc_hd__dfxtp_1 _544_ (.CLK(clknet_3_7__leaf_io_in[0]),
    .D(_038_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\f_fifo.fifo_data[2][1] ));
 sky130_fd_sc_hd__dfxtp_1 _545_ (.CLK(clknet_3_7__leaf_io_in[0]),
    .D(_039_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\f_fifo.fifo_data[2][2] ));
 sky130_fd_sc_hd__dfxtp_1 _546_ (.CLK(clknet_3_0__leaf_io_in[0]),
    .D(_040_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\f_fifo.fifo_data[2][3] ));
 sky130_fd_sc_hd__dfxtp_1 _547_ (.CLK(clknet_3_3__leaf_io_in[0]),
    .D(_041_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\f_fifo.fifo_data[2][4] ));
 sky130_fd_sc_hd__dfxtp_1 _548_ (.CLK(clknet_3_4__leaf_io_in[0]),
    .D(_042_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\f_fifo.fifo_data[2][5] ));
 sky130_fd_sc_hd__dfxtp_1 _549_ (.CLK(clknet_3_5__leaf_io_in[0]),
    .D(_043_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\f_fifo.fifo_data[3][0] ));
 sky130_fd_sc_hd__dfxtp_1 _550_ (.CLK(clknet_3_0__leaf_io_in[0]),
    .D(_044_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\f_fifo.fifo_data[3][1] ));
 sky130_fd_sc_hd__dfxtp_1 _551_ (.CLK(clknet_3_0__leaf_io_in[0]),
    .D(_045_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\f_fifo.fifo_data[3][2] ));
 sky130_fd_sc_hd__dfxtp_1 _552_ (.CLK(clknet_3_3__leaf_io_in[0]),
    .D(_046_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\f_fifo.fifo_data[3][3] ));
 sky130_fd_sc_hd__dfxtp_1 _553_ (.CLK(clknet_3_3__leaf_io_in[0]),
    .D(_047_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\f_fifo.fifo_data[3][4] ));
 sky130_fd_sc_hd__dfxtp_1 _554_ (.CLK(clknet_3_4__leaf_io_in[0]),
    .D(_048_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\f_fifo.fifo_data[3][5] ));
 sky130_fd_sc_hd__dfxtp_1 _555_ (.CLK(clknet_3_6__leaf_io_in[0]),
    .D(reset_n_in),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\f_fifo.reset_n ));
 sky130_fd_sc_hd__dfxtp_1 _556_ (.CLK(clknet_3_2__leaf_io_in[0]),
    .D(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[47].entry.write_in ));
 sky130_fd_sc_hd__dfxtp_2 _557_ (.CLK(clknet_3_7__leaf_io_in[0]),
    .D(_049_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(io_out[2]));
 sky130_fd_sc_hd__dfxtp_2 _558_ (.CLK(clknet_3_7__leaf_io_in[0]),
    .D(_050_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(io_out[3]));
 sky130_fd_sc_hd__dfxtp_2 _559_ (.CLK(clknet_3_6__leaf_io_in[0]),
    .D(_051_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(io_out[4]));
 sky130_fd_sc_hd__dfxtp_2 _560_ (.CLK(clknet_3_6__leaf_io_in[0]),
    .D(_052_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(io_out[5]));
 sky130_fd_sc_hd__dfxtp_2 _561_ (.CLK(clknet_3_2__leaf_io_in[0]),
    .D(_053_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(io_out[6]));
 sky130_fd_sc_hd__dfxtp_2 _562_ (.CLK(clknet_3_0__leaf_io_in[0]),
    .D(_054_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(io_out[7]));
 sky130_fd_sc_hd__dfxtp_2 _563_ (.CLK(clknet_3_2__leaf_io_in[0]),
    .D(_055_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[10].entry.next_is_empty ));
 sky130_fd_sc_hd__dfxtp_2 _564_ (.CLK(clknet_3_2__leaf_io_in[0]),
    .D(_056_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[46].entry.empty ));
 sky130_fd_sc_hd__dfxtp_2 _565_ (.CLK(clknet_3_6__leaf_io_in[0]),
    .D(_057_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[45].entry.empty ));
 sky130_fd_sc_hd__dfxtp_2 _566_ (.CLK(clknet_3_5__leaf_io_in[0]),
    .D(_058_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[44].entry.empty ));
 sky130_fd_sc_hd__dfxtp_2 _567_ (.CLK(clknet_3_3__leaf_io_in[0]),
    .D(_059_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[43].entry.empty ));
 sky130_fd_sc_hd__dfxtp_2 _568_ (.CLK(clknet_3_0__leaf_io_in[0]),
    .D(_060_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[42].entry.empty ));
 sky130_fd_sc_hd__dfxtp_2 _569_ (.CLK(clknet_3_3__leaf_io_in[0]),
    .D(_061_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[41].entry.empty ));
 sky130_fd_sc_hd__dfxtp_2 _570_ (.CLK(clknet_3_2__leaf_io_in[0]),
    .D(_062_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[40].entry.empty ));
 sky130_fd_sc_hd__dfxtp_2 _571_ (.CLK(clknet_3_1__leaf_io_in[0]),
    .D(_063_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[3].entry.empty ));
 sky130_fd_sc_hd__dfxtp_2 _572_ (.CLK(clknet_3_1__leaf_io_in[0]),
    .D(_064_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[38].entry.empty ));
 sky130_fd_sc_hd__dfxtp_2 _573_ (.CLK(clknet_3_2__leaf_io_in[0]),
    .D(_065_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[37].entry.empty ));
 sky130_fd_sc_hd__dfxtp_2 _574_ (.CLK(clknet_3_4__leaf_io_in[0]),
    .D(_066_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[36].entry.empty ));
 sky130_fd_sc_hd__dfxtp_2 _575_ (.CLK(clknet_3_1__leaf_io_in[0]),
    .D(_067_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[35].entry.empty ));
 sky130_fd_sc_hd__dfxtp_4 _576_ (.CLK(clknet_3_5__leaf_io_in[0]),
    .D(_068_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[34].entry.empty ));
 sky130_fd_sc_hd__dfxtp_2 _577_ (.CLK(clknet_3_3__leaf_io_in[0]),
    .D(_069_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[33].entry.empty ));
 sky130_fd_sc_hd__dfxtp_2 _578_ (.CLK(clknet_3_3__leaf_io_in[0]),
    .D(_070_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[32].entry.empty ));
 sky130_fd_sc_hd__dfxtp_2 _579_ (.CLK(clknet_3_2__leaf_io_in[0]),
    .D(_071_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[31].entry.empty ));
 sky130_fd_sc_hd__dfxtp_2 _580_ (.CLK(clknet_3_1__leaf_io_in[0]),
    .D(_072_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[30].entry.empty ));
 sky130_fd_sc_hd__dfxtp_2 _581_ (.CLK(clknet_3_7__leaf_io_in[0]),
    .D(_073_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[2].entry.empty ));
 sky130_fd_sc_hd__dfxtp_2 _582_ (.CLK(clknet_3_2__leaf_io_in[0]),
    .D(_074_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[28].entry.empty ));
 sky130_fd_sc_hd__dfxtp_2 _583_ (.CLK(clknet_3_2__leaf_io_in[0]),
    .D(_075_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[27].entry.empty ));
 sky130_fd_sc_hd__dfxtp_2 _584_ (.CLK(clknet_3_0__leaf_io_in[0]),
    .D(_076_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[26].entry.empty ));
 sky130_fd_sc_hd__dfxtp_2 _585_ (.CLK(clknet_3_4__leaf_io_in[0]),
    .D(_077_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[25].entry.empty ));
 sky130_fd_sc_hd__dfxtp_2 _586_ (.CLK(clknet_3_1__leaf_io_in[0]),
    .D(_078_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[24].entry.empty ));
 sky130_fd_sc_hd__dfxtp_2 _587_ (.CLK(clknet_3_5__leaf_io_in[0]),
    .D(_079_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[23].entry.empty ));
 sky130_fd_sc_hd__dfxtp_2 _588_ (.CLK(clknet_3_1__leaf_io_in[0]),
    .D(_080_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[22].entry.empty ));
 sky130_fd_sc_hd__dfxtp_2 _589_ (.CLK(clknet_3_1__leaf_io_in[0]),
    .D(_081_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[21].entry.empty ));
 sky130_fd_sc_hd__dfxtp_2 _590_ (.CLK(clknet_3_2__leaf_io_in[0]),
    .D(_082_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[20].entry.empty ));
 sky130_fd_sc_hd__dfxtp_2 _591_ (.CLK(clknet_3_2__leaf_io_in[0]),
    .D(_083_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[1].entry.empty ));
 sky130_fd_sc_hd__dfxtp_2 _592_ (.CLK(clknet_3_5__leaf_io_in[0]),
    .D(_084_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[18].entry.empty ));
 sky130_fd_sc_hd__dfxtp_4 _593_ (.CLK(clknet_3_2__leaf_io_in[0]),
    .D(_085_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[17].entry.empty ));
 sky130_fd_sc_hd__dfxtp_2 _594_ (.CLK(clknet_3_0__leaf_io_in[0]),
    .D(_086_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[16].entry.empty ));
 sky130_fd_sc_hd__dfxtp_2 _595_ (.CLK(clknet_3_4__leaf_io_in[0]),
    .D(_087_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[15].entry.empty ));
 sky130_fd_sc_hd__dfxtp_2 _596_ (.CLK(clknet_3_6__leaf_io_in[0]),
    .D(_088_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[14].entry.empty ));
 sky130_fd_sc_hd__buf_2 _597_ (.A(\l_fifo.ready ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(io_out[0]));
 sky130_fd_sc_hd__buf_2 _598_ (.A(\f_fifo.empty_n ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(io_out[1]));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_io_in[0]  (.A(io_in[0]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(clknet_0_io_in[0]));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_3_0__f_io_in[0]  (.A(clknet_0_io_in[0]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(clknet_3_0__leaf_io_in[0]));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_3_1__f_io_in[0]  (.A(clknet_0_io_in[0]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(clknet_3_1__leaf_io_in[0]));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_3_2__f_io_in[0]  (.A(clknet_0_io_in[0]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(clknet_3_2__leaf_io_in[0]));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_3_3__f_io_in[0]  (.A(clknet_0_io_in[0]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(clknet_3_3__leaf_io_in[0]));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_3_4__f_io_in[0]  (.A(clknet_0_io_in[0]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(clknet_3_4__leaf_io_in[0]));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_3_5__f_io_in[0]  (.A(clknet_0_io_in[0]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(clknet_3_5__leaf_io_in[0]));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_3_6__f_io_in[0]  (.A(clknet_0_io_in[0]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(clknet_3_6__leaf_io_in[0]));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_3_7__f_io_in[0]  (.A(clknet_0_io_in[0]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(clknet_3_7__leaf_io_in[0]));
 sky130_fd_sc_hd__clkbuf_1 \data_in_buffer[0].genblk1[0].genblk1.buf_first  (.A(\data_in_buffer[0].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\data_in_buffer[0].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \data_in_buffer[0].genblk1[0].genblk2.buf2  (.A(\data_in_buffer[0].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\data_in_buffer[0].b[0] ));
 sky130_fd_sc_hd__clkbuf_1 \data_in_buffer[0].genblk1[1].genblk1.buf1  (.A(\data_in_buffer[0].b[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\data_in_buffer[0].genblk1[1].mid ));
 sky130_fd_sc_hd__clkbuf_1 \data_in_buffer[0].genblk1[1].genblk2.buf_last  (.A(\data_in_buffer[0].genblk1[1].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\data_in_buffer[0].X ));
 sky130_fd_sc_hd__clkbuf_1 \data_in_buffer[1].genblk1[0].genblk1.buf_first  (.A(\data_in_buffer[1].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\data_in_buffer[1].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \data_in_buffer[1].genblk1[0].genblk2.buf2  (.A(\data_in_buffer[1].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\data_in_buffer[1].b[0] ));
 sky130_fd_sc_hd__clkbuf_1 \data_in_buffer[1].genblk1[1].genblk1.buf1  (.A(\data_in_buffer[1].b[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\data_in_buffer[1].genblk1[1].mid ));
 sky130_fd_sc_hd__clkbuf_1 \data_in_buffer[1].genblk1[1].genblk2.buf_last  (.A(\data_in_buffer[1].genblk1[1].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\data_in_buffer[1].X ));
 sky130_fd_sc_hd__clkbuf_1 \data_in_buffer[2].genblk1[0].genblk1.buf_first  (.A(\data_in_buffer[2].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\data_in_buffer[2].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \data_in_buffer[2].genblk1[0].genblk2.buf2  (.A(\data_in_buffer[2].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\data_in_buffer[2].b[0] ));
 sky130_fd_sc_hd__clkbuf_1 \data_in_buffer[2].genblk1[1].genblk1.buf1  (.A(\data_in_buffer[2].b[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\data_in_buffer[2].genblk1[1].mid ));
 sky130_fd_sc_hd__clkbuf_1 \data_in_buffer[2].genblk1[1].genblk2.buf_last  (.A(\data_in_buffer[2].genblk1[1].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\data_in_buffer[2].X ));
 sky130_fd_sc_hd__clkbuf_1 \data_in_buffer[3].genblk1[0].genblk1.buf_first  (.A(\data_in_buffer[3].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\data_in_buffer[3].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \data_in_buffer[3].genblk1[0].genblk2.buf2  (.A(\data_in_buffer[3].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\data_in_buffer[3].b[0] ));
 sky130_fd_sc_hd__clkbuf_1 \data_in_buffer[3].genblk1[1].genblk1.buf1  (.A(\data_in_buffer[3].b[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\data_in_buffer[3].genblk1[1].mid ));
 sky130_fd_sc_hd__clkbuf_1 \data_in_buffer[3].genblk1[1].genblk2.buf_last  (.A(\data_in_buffer[3].genblk1[1].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\data_in_buffer[3].X ));
 sky130_fd_sc_hd__clkbuf_1 \data_in_buffer[4].genblk1[0].genblk1.buf_first  (.A(\data_in_buffer[4].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\data_in_buffer[4].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \data_in_buffer[4].genblk1[0].genblk2.buf2  (.A(\data_in_buffer[4].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\data_in_buffer[4].b[0] ));
 sky130_fd_sc_hd__clkbuf_1 \data_in_buffer[4].genblk1[1].genblk1.buf1  (.A(\data_in_buffer[4].b[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\data_in_buffer[4].genblk1[1].mid ));
 sky130_fd_sc_hd__clkbuf_1 \data_in_buffer[4].genblk1[1].genblk2.buf_last  (.A(\data_in_buffer[4].genblk1[1].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\data_in_buffer[4].X ));
 sky130_fd_sc_hd__clkbuf_1 \data_in_buffer[5].genblk1[0].genblk1.buf_first  (.A(\data_in_buffer[5].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\data_in_buffer[5].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \data_in_buffer[5].genblk1[0].genblk2.buf2  (.A(\data_in_buffer[5].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\data_in_buffer[5].b[0] ));
 sky130_fd_sc_hd__clkbuf_1 \data_in_buffer[5].genblk1[1].genblk1.buf1  (.A(\data_in_buffer[5].b[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\data_in_buffer[5].genblk1[1].mid ));
 sky130_fd_sc_hd__clkbuf_1 \data_in_buffer[5].genblk1[1].genblk2.buf_last  (.A(\data_in_buffer[5].genblk1[1].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\data_in_buffer[5].X ));
 sky130_fd_sc_hd__buf_2 fanout10 (.A(net13),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net10));
 sky130_fd_sc_hd__buf_2 fanout11 (.A(net13),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net11));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout12 (.A(net13),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net12));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout13 (.A(net25),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net13));
 sky130_fd_sc_hd__buf_2 fanout14 (.A(net17),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net14));
 sky130_fd_sc_hd__buf_2 fanout15 (.A(net17),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_2 fanout16 (.A(net17),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net16));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout17 (.A(net25),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net17));
 sky130_fd_sc_hd__buf_2 fanout18 (.A(net21),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net18));
 sky130_fd_sc_hd__buf_2 fanout19 (.A(net21),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net19));
 sky130_fd_sc_hd__clkbuf_2 fanout20 (.A(net21),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net20));
 sky130_fd_sc_hd__clkbuf_2 fanout21 (.A(net25),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net21));
 sky130_fd_sc_hd__buf_2 fanout22 (.A(net24),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net22));
 sky130_fd_sc_hd__buf_2 fanout23 (.A(net24),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net23));
 sky130_fd_sc_hd__clkbuf_2 fanout24 (.A(net25),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net24));
 sky130_fd_sc_hd__clkbuf_2 fanout25 (.A(\f_fifo.reset_n ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net25));
 sky130_fd_sc_hd__buf_2 fanout26 (.A(net27),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net26));
 sky130_fd_sc_hd__buf_2 fanout27 (.A(net49),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net27));
 sky130_fd_sc_hd__buf_2 fanout28 (.A(net29),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net28));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout29 (.A(net34),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net29));
 sky130_fd_sc_hd__buf_2 fanout30 (.A(net34),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net30));
 sky130_fd_sc_hd__clkbuf_2 fanout31 (.A(net34),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net31));
 sky130_fd_sc_hd__buf_2 fanout32 (.A(net34),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net32));
 sky130_fd_sc_hd__clkbuf_2 fanout33 (.A(net34),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net33));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout34 (.A(net49),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net34));
 sky130_fd_sc_hd__buf_2 fanout35 (.A(net38),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net35));
 sky130_fd_sc_hd__buf_2 fanout36 (.A(net38),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net36));
 sky130_fd_sc_hd__clkbuf_2 fanout37 (.A(net38),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net37));
 sky130_fd_sc_hd__clkbuf_2 fanout38 (.A(net49),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net38));
 sky130_fd_sc_hd__buf_2 fanout39 (.A(net42),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net39));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout40 (.A(net42),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net40));
 sky130_fd_sc_hd__buf_2 fanout41 (.A(net42),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net41));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout42 (.A(net49),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net42));
 sky130_fd_sc_hd__buf_2 fanout43 (.A(net48),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net43));
 sky130_fd_sc_hd__buf_2 fanout44 (.A(net48),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net44));
 sky130_fd_sc_hd__clkbuf_2 fanout45 (.A(net48),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net45));
 sky130_fd_sc_hd__buf_2 fanout46 (.A(net47),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net46));
 sky130_fd_sc_hd__buf_2 fanout47 (.A(net48),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net47));
 sky130_fd_sc_hd__clkbuf_2 fanout48 (.A(net49),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net48));
 sky130_fd_sc_hd__buf_2 fanout49 (.A(\f_fifo.reset_n ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net49));
 sky130_fd_sc_hd__buf_2 fanout8 (.A(net25),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_2 fanout9 (.A(net25),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net9));
 sky130_fd_sc_hd__buf_2 input1 (.A(io_in[1]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1));
 sky130_fd_sc_hd__dlymetal6s2s_1 input2 (.A(io_in[2]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net2));
 sky130_fd_sc_hd__dlymetal6s2s_1 input3 (.A(io_in[3]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net3));
 sky130_fd_sc_hd__dlymetal6s2s_1 input4 (.A(io_in[4]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_1 input5 (.A(io_in[5]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_1 input6 (.A(io_in[6]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_1 input7 (.A(io_in[7]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[0].entry.input_buf[0].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[0].entry.input_buf[0].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[0].entry.input_buf[0].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[0].entry.input_buf[0].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[0].entry.input_buf[0].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[0].entry.input_buf[0].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[0].entry.input_buf[1].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[0].entry.input_buf[1].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[0].entry.input_buf[1].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[0].entry.input_buf[1].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[0].entry.input_buf[1].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[0].entry.input_buf[1].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[0].entry.input_buf[2].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[0].entry.input_buf[2].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[0].entry.input_buf[2].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[0].entry.input_buf[2].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[0].entry.input_buf[2].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[0].entry.input_buf[2].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[0].entry.input_buf[3].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[0].entry.input_buf[3].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[0].entry.input_buf[3].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[0].entry.input_buf[3].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[0].entry.input_buf[3].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[0].entry.input_buf[3].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[0].entry.input_buf[4].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[0].entry.input_buf[4].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[0].entry.input_buf[4].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[0].entry.input_buf[4].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[0].entry.input_buf[4].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[0].entry.input_buf[4].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[0].entry.input_buf[5].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[0].entry.input_buf[5].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[0].entry.input_buf[5].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[0].entry.input_buf[5].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[0].entry.input_buf[5].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[0].entry.input_buf[5].X ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[0].entry.latch[0]  (.D(\l_fifo.genblk1[0].entry.input_buf[0].X ),
    .GATE(\l_fifo.genblk1[0].entry.empty ),
    .RESET_B(net26),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\f_fifo.data_in[0] ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[0].entry.latch[1]  (.D(\l_fifo.genblk1[0].entry.input_buf[1].X ),
    .GATE(\l_fifo.genblk1[0].entry.empty ),
    .RESET_B(net35),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\f_fifo.data_in[1] ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[0].entry.latch[2]  (.D(\l_fifo.genblk1[0].entry.input_buf[2].X ),
    .GATE(\l_fifo.genblk1[0].entry.empty ),
    .RESET_B(net9),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\f_fifo.data_in[2] ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[0].entry.latch[3]  (.D(\l_fifo.genblk1[0].entry.input_buf[3].X ),
    .GATE(\l_fifo.genblk1[0].entry.empty ),
    .RESET_B(net8),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\f_fifo.data_in[3] ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[0].entry.latch[4]  (.D(\l_fifo.genblk1[0].entry.input_buf[4].X ),
    .GATE(\l_fifo.genblk1[0].entry.empty ),
    .RESET_B(net19),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\f_fifo.data_in[4] ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[0].entry.latch[5]  (.D(\l_fifo.genblk1[0].entry.input_buf[5].X ),
    .GATE(\l_fifo.genblk1[0].entry.empty ),
    .RESET_B(net26),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\f_fifo.data_in[5] ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[10].entry.input_buf[0].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[10].entry.input_buf[0].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[10].entry.input_buf[0].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[10].entry.input_buf[0].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[10].entry.input_buf[0].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[10].entry.input_buf[0].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[10].entry.input_buf[1].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[10].entry.input_buf[1].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[10].entry.input_buf[1].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[10].entry.input_buf[1].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[10].entry.input_buf[1].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[10].entry.input_buf[1].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[10].entry.input_buf[2].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[10].entry.input_buf[2].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[10].entry.input_buf[2].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[10].entry.input_buf[2].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[10].entry.input_buf[2].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[10].entry.input_buf[2].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[10].entry.input_buf[3].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[10].entry.input_buf[3].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[10].entry.input_buf[3].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[10].entry.input_buf[3].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[10].entry.input_buf[3].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[10].entry.input_buf[3].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[10].entry.input_buf[4].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[10].entry.input_buf[4].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[10].entry.input_buf[4].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[10].entry.input_buf[4].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[10].entry.input_buf[4].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[10].entry.input_buf[4].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[10].entry.input_buf[5].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[10].entry.input_buf[5].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[10].entry.input_buf[5].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[10].entry.input_buf[5].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[10].entry.input_buf[5].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[10].entry.input_buf[5].X ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[10].entry.latch[0]  (.D(\l_fifo.genblk1[10].entry.input_buf[0].X ),
    .GATE(\l_fifo.genblk1[10].entry.empty ),
    .RESET_B(net44),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[9].entry.input_buf[0].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[10].entry.latch[1]  (.D(\l_fifo.genblk1[10].entry.input_buf[1].X ),
    .GATE(\l_fifo.genblk1[10].entry.empty ),
    .RESET_B(net43),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[9].entry.input_buf[1].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[10].entry.latch[2]  (.D(\l_fifo.genblk1[10].entry.input_buf[2].X ),
    .GATE(\l_fifo.genblk1[10].entry.empty ),
    .RESET_B(net43),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[9].entry.input_buf[2].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[10].entry.latch[3]  (.D(\l_fifo.genblk1[10].entry.input_buf[3].X ),
    .GATE(\l_fifo.genblk1[10].entry.empty ),
    .RESET_B(net43),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[9].entry.input_buf[3].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[10].entry.latch[4]  (.D(\l_fifo.genblk1[10].entry.input_buf[4].X ),
    .GATE(\l_fifo.genblk1[10].entry.empty ),
    .RESET_B(net33),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[9].entry.input_buf[4].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[10].entry.latch[5]  (.D(\l_fifo.genblk1[10].entry.input_buf[5].X ),
    .GATE(\l_fifo.genblk1[10].entry.empty ),
    .RESET_B(net43),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[9].entry.input_buf[5].A ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[11].entry.input_buf[0].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[11].entry.input_buf[0].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[11].entry.input_buf[0].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[11].entry.input_buf[0].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[11].entry.input_buf[0].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[11].entry.input_buf[0].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[11].entry.input_buf[1].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[11].entry.input_buf[1].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[11].entry.input_buf[1].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[11].entry.input_buf[1].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[11].entry.input_buf[1].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[11].entry.input_buf[1].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[11].entry.input_buf[2].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[11].entry.input_buf[2].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[11].entry.input_buf[2].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[11].entry.input_buf[2].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[11].entry.input_buf[2].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[11].entry.input_buf[2].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[11].entry.input_buf[3].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[11].entry.input_buf[3].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[11].entry.input_buf[3].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[11].entry.input_buf[3].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[11].entry.input_buf[3].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[11].entry.input_buf[3].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[11].entry.input_buf[4].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[11].entry.input_buf[4].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[11].entry.input_buf[4].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[11].entry.input_buf[4].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[11].entry.input_buf[4].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[11].entry.input_buf[4].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[11].entry.input_buf[5].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[11].entry.input_buf[5].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[11].entry.input_buf[5].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[11].entry.input_buf[5].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[11].entry.input_buf[5].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[11].entry.input_buf[5].X ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[11].entry.latch[0]  (.D(\l_fifo.genblk1[11].entry.input_buf[0].X ),
    .GATE(\l_fifo.genblk1[11].entry.empty ),
    .RESET_B(net33),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[10].entry.input_buf[0].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[11].entry.latch[1]  (.D(\l_fifo.genblk1[11].entry.input_buf[1].X ),
    .GATE(\l_fifo.genblk1[11].entry.empty ),
    .RESET_B(net43),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[10].entry.input_buf[1].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[11].entry.latch[2]  (.D(\l_fifo.genblk1[11].entry.input_buf[2].X ),
    .GATE(\l_fifo.genblk1[11].entry.empty ),
    .RESET_B(net44),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[10].entry.input_buf[2].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[11].entry.latch[3]  (.D(\l_fifo.genblk1[11].entry.input_buf[3].X ),
    .GATE(\l_fifo.genblk1[11].entry.empty ),
    .RESET_B(net45),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[10].entry.input_buf[3].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[11].entry.latch[4]  (.D(\l_fifo.genblk1[11].entry.input_buf[4].X ),
    .GATE(\l_fifo.genblk1[11].entry.empty ),
    .RESET_B(net33),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[10].entry.input_buf[4].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[11].entry.latch[5]  (.D(\l_fifo.genblk1[11].entry.input_buf[5].X ),
    .GATE(\l_fifo.genblk1[11].entry.empty ),
    .RESET_B(net44),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[10].entry.input_buf[5].A ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[12].entry.input_buf[0].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[12].entry.input_buf[0].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[12].entry.input_buf[0].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[12].entry.input_buf[0].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[12].entry.input_buf[0].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[12].entry.input_buf[0].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[12].entry.input_buf[1].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[12].entry.input_buf[1].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[12].entry.input_buf[1].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[12].entry.input_buf[1].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[12].entry.input_buf[1].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[12].entry.input_buf[1].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[12].entry.input_buf[2].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[12].entry.input_buf[2].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[12].entry.input_buf[2].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[12].entry.input_buf[2].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[12].entry.input_buf[2].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[12].entry.input_buf[2].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[12].entry.input_buf[3].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[12].entry.input_buf[3].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[12].entry.input_buf[3].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[12].entry.input_buf[3].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[12].entry.input_buf[3].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[12].entry.input_buf[3].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[12].entry.input_buf[4].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[12].entry.input_buf[4].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[12].entry.input_buf[4].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[12].entry.input_buf[4].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[12].entry.input_buf[4].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[12].entry.input_buf[4].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[12].entry.input_buf[5].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[12].entry.input_buf[5].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[12].entry.input_buf[5].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[12].entry.input_buf[5].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[12].entry.input_buf[5].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[12].entry.input_buf[5].X ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[12].entry.latch[0]  (.D(\l_fifo.genblk1[12].entry.input_buf[0].X ),
    .GATE(\l_fifo.genblk1[12].entry.empty ),
    .RESET_B(net30),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[11].entry.input_buf[0].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[12].entry.latch[1]  (.D(\l_fifo.genblk1[12].entry.input_buf[1].X ),
    .GATE(\l_fifo.genblk1[12].entry.empty ),
    .RESET_B(net45),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[11].entry.input_buf[1].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[12].entry.latch[2]  (.D(\l_fifo.genblk1[12].entry.input_buf[2].X ),
    .GATE(\l_fifo.genblk1[12].entry.empty ),
    .RESET_B(net44),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[11].entry.input_buf[2].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[12].entry.latch[3]  (.D(\l_fifo.genblk1[12].entry.input_buf[3].X ),
    .GATE(\l_fifo.genblk1[12].entry.empty ),
    .RESET_B(net45),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[11].entry.input_buf[3].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[12].entry.latch[4]  (.D(\l_fifo.genblk1[12].entry.input_buf[4].X ),
    .GATE(\l_fifo.genblk1[12].entry.empty ),
    .RESET_B(net33),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[11].entry.input_buf[4].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[12].entry.latch[5]  (.D(\l_fifo.genblk1[12].entry.input_buf[5].X ),
    .GATE(\l_fifo.genblk1[12].entry.empty ),
    .RESET_B(net44),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[11].entry.input_buf[5].A ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[13].entry.input_buf[0].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[13].entry.input_buf[0].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[13].entry.input_buf[0].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[13].entry.input_buf[0].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[13].entry.input_buf[0].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[13].entry.input_buf[0].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[13].entry.input_buf[1].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[13].entry.input_buf[1].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[13].entry.input_buf[1].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[13].entry.input_buf[1].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[13].entry.input_buf[1].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[13].entry.input_buf[1].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[13].entry.input_buf[2].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[13].entry.input_buf[2].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[13].entry.input_buf[2].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[13].entry.input_buf[2].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[13].entry.input_buf[2].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[13].entry.input_buf[2].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[13].entry.input_buf[3].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[13].entry.input_buf[3].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[13].entry.input_buf[3].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[13].entry.input_buf[3].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[13].entry.input_buf[3].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[13].entry.input_buf[3].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[13].entry.input_buf[4].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[13].entry.input_buf[4].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[13].entry.input_buf[4].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[13].entry.input_buf[4].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[13].entry.input_buf[4].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[13].entry.input_buf[4].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[13].entry.input_buf[5].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[13].entry.input_buf[5].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[13].entry.input_buf[5].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[13].entry.input_buf[5].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[13].entry.input_buf[5].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[13].entry.input_buf[5].X ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[13].entry.latch[0]  (.D(\l_fifo.genblk1[13].entry.input_buf[0].X ),
    .GATE(\l_fifo.genblk1[13].entry.empty ),
    .RESET_B(net43),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[12].entry.input_buf[0].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[13].entry.latch[1]  (.D(\l_fifo.genblk1[13].entry.input_buf[1].X ),
    .GATE(\l_fifo.genblk1[13].entry.empty ),
    .RESET_B(net44),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[12].entry.input_buf[1].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[13].entry.latch[2]  (.D(\l_fifo.genblk1[13].entry.input_buf[2].X ),
    .GATE(\l_fifo.genblk1[13].entry.empty ),
    .RESET_B(net45),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[12].entry.input_buf[2].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[13].entry.latch[3]  (.D(\l_fifo.genblk1[13].entry.input_buf[3].X ),
    .GATE(\l_fifo.genblk1[13].entry.empty ),
    .RESET_B(net44),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[12].entry.input_buf[3].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[13].entry.latch[4]  (.D(\l_fifo.genblk1[13].entry.input_buf[4].X ),
    .GATE(\l_fifo.genblk1[13].entry.empty ),
    .RESET_B(net44),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[12].entry.input_buf[4].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[13].entry.latch[5]  (.D(\l_fifo.genblk1[13].entry.input_buf[5].X ),
    .GATE(\l_fifo.genblk1[13].entry.empty ),
    .RESET_B(net44),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[12].entry.input_buf[5].A ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[14].entry.input_buf[0].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[14].entry.input_buf[0].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[14].entry.input_buf[0].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[14].entry.input_buf[0].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[14].entry.input_buf[0].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[14].entry.input_buf[0].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[14].entry.input_buf[1].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[14].entry.input_buf[1].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[14].entry.input_buf[1].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[14].entry.input_buf[1].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[14].entry.input_buf[1].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[14].entry.input_buf[1].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[14].entry.input_buf[2].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[14].entry.input_buf[2].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[14].entry.input_buf[2].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[14].entry.input_buf[2].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[14].entry.input_buf[2].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[14].entry.input_buf[2].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[14].entry.input_buf[3].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[14].entry.input_buf[3].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[14].entry.input_buf[3].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[14].entry.input_buf[3].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[14].entry.input_buf[3].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[14].entry.input_buf[3].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[14].entry.input_buf[4].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[14].entry.input_buf[4].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[14].entry.input_buf[4].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[14].entry.input_buf[4].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[14].entry.input_buf[4].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[14].entry.input_buf[4].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[14].entry.input_buf[5].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[14].entry.input_buf[5].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[14].entry.input_buf[5].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[14].entry.input_buf[5].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[14].entry.input_buf[5].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[14].entry.input_buf[5].X ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[14].entry.latch[0]  (.D(\l_fifo.genblk1[14].entry.input_buf[0].X ),
    .GATE(\l_fifo.genblk1[14].entry.empty ),
    .RESET_B(net43),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[13].entry.input_buf[0].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[14].entry.latch[1]  (.D(\l_fifo.genblk1[14].entry.input_buf[1].X ),
    .GATE(\l_fifo.genblk1[14].entry.empty ),
    .RESET_B(net45),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[13].entry.input_buf[1].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[14].entry.latch[2]  (.D(\l_fifo.genblk1[14].entry.input_buf[2].X ),
    .GATE(\l_fifo.genblk1[14].entry.empty ),
    .RESET_B(net45),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[13].entry.input_buf[2].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[14].entry.latch[3]  (.D(\l_fifo.genblk1[14].entry.input_buf[3].X ),
    .GATE(\l_fifo.genblk1[14].entry.empty ),
    .RESET_B(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[13].entry.input_buf[3].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[14].entry.latch[4]  (.D(\l_fifo.genblk1[14].entry.input_buf[4].X ),
    .GATE(\l_fifo.genblk1[14].entry.empty ),
    .RESET_B(net45),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[13].entry.input_buf[4].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[14].entry.latch[5]  (.D(\l_fifo.genblk1[14].entry.input_buf[5].X ),
    .GATE(\l_fifo.genblk1[14].entry.empty ),
    .RESET_B(net43),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[13].entry.input_buf[5].A ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[15].entry.input_buf[0].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[15].entry.input_buf[0].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[15].entry.input_buf[0].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[15].entry.input_buf[0].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[15].entry.input_buf[0].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[15].entry.input_buf[0].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[15].entry.input_buf[1].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[15].entry.input_buf[1].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[15].entry.input_buf[1].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[15].entry.input_buf[1].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[15].entry.input_buf[1].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[15].entry.input_buf[1].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[15].entry.input_buf[2].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[15].entry.input_buf[2].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[15].entry.input_buf[2].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[15].entry.input_buf[2].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[15].entry.input_buf[2].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[15].entry.input_buf[2].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[15].entry.input_buf[3].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[15].entry.input_buf[3].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[15].entry.input_buf[3].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[15].entry.input_buf[3].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[15].entry.input_buf[3].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[15].entry.input_buf[3].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[15].entry.input_buf[4].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[15].entry.input_buf[4].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[15].entry.input_buf[4].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[15].entry.input_buf[4].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[15].entry.input_buf[4].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[15].entry.input_buf[4].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[15].entry.input_buf[5].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[15].entry.input_buf[5].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[15].entry.input_buf[5].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[15].entry.input_buf[5].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[15].entry.input_buf[5].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[15].entry.input_buf[5].X ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[15].entry.latch[0]  (.D(\l_fifo.genblk1[15].entry.input_buf[0].X ),
    .GATE(\l_fifo.genblk1[15].entry.empty ),
    .RESET_B(net47),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[14].entry.input_buf[0].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[15].entry.latch[1]  (.D(\l_fifo.genblk1[15].entry.input_buf[1].X ),
    .GATE(\l_fifo.genblk1[15].entry.empty ),
    .RESET_B(net48),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[14].entry.input_buf[1].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[15].entry.latch[2]  (.D(\l_fifo.genblk1[15].entry.input_buf[2].X ),
    .GATE(\l_fifo.genblk1[15].entry.empty ),
    .RESET_B(net47),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[14].entry.input_buf[2].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[15].entry.latch[3]  (.D(\l_fifo.genblk1[15].entry.input_buf[3].X ),
    .GATE(\l_fifo.genblk1[15].entry.empty ),
    .RESET_B(net46),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[14].entry.input_buf[3].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[15].entry.latch[4]  (.D(\l_fifo.genblk1[15].entry.input_buf[4].X ),
    .GATE(\l_fifo.genblk1[15].entry.empty ),
    .RESET_B(net47),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[14].entry.input_buf[4].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[15].entry.latch[5]  (.D(\l_fifo.genblk1[15].entry.input_buf[5].X ),
    .GATE(\l_fifo.genblk1[15].entry.empty ),
    .RESET_B(net37),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[14].entry.input_buf[5].A ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[16].entry.input_buf[0].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[16].entry.input_buf[0].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[16].entry.input_buf[0].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[16].entry.input_buf[0].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[16].entry.input_buf[0].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[16].entry.input_buf[0].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[16].entry.input_buf[1].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[16].entry.input_buf[1].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[16].entry.input_buf[1].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[16].entry.input_buf[1].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[16].entry.input_buf[1].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[16].entry.input_buf[1].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[16].entry.input_buf[2].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[16].entry.input_buf[2].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[16].entry.input_buf[2].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[16].entry.input_buf[2].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[16].entry.input_buf[2].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[16].entry.input_buf[2].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[16].entry.input_buf[3].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[16].entry.input_buf[3].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[16].entry.input_buf[3].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[16].entry.input_buf[3].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[16].entry.input_buf[3].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[16].entry.input_buf[3].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[16].entry.input_buf[4].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[16].entry.input_buf[4].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[16].entry.input_buf[4].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[16].entry.input_buf[4].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[16].entry.input_buf[4].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[16].entry.input_buf[4].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[16].entry.input_buf[5].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[16].entry.input_buf[5].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[16].entry.input_buf[5].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[16].entry.input_buf[5].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[16].entry.input_buf[5].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[16].entry.input_buf[5].X ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[16].entry.latch[0]  (.D(\l_fifo.genblk1[16].entry.input_buf[0].X ),
    .GATE(\l_fifo.genblk1[16].entry.empty ),
    .RESET_B(net47),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[15].entry.input_buf[0].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[16].entry.latch[1]  (.D(\l_fifo.genblk1[16].entry.input_buf[1].X ),
    .GATE(\l_fifo.genblk1[16].entry.empty ),
    .RESET_B(net47),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[15].entry.input_buf[1].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[16].entry.latch[2]  (.D(\l_fifo.genblk1[16].entry.input_buf[2].X ),
    .GATE(\l_fifo.genblk1[16].entry.empty ),
    .RESET_B(net46),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[15].entry.input_buf[2].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[16].entry.latch[3]  (.D(\l_fifo.genblk1[16].entry.input_buf[3].X ),
    .GATE(\l_fifo.genblk1[16].entry.empty ),
    .RESET_B(net47),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[15].entry.input_buf[3].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[16].entry.latch[4]  (.D(\l_fifo.genblk1[16].entry.input_buf[4].X ),
    .GATE(\l_fifo.genblk1[16].entry.empty ),
    .RESET_B(net47),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[15].entry.input_buf[4].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[16].entry.latch[5]  (.D(\l_fifo.genblk1[16].entry.input_buf[5].X ),
    .GATE(\l_fifo.genblk1[16].entry.empty ),
    .RESET_B(net46),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[15].entry.input_buf[5].A ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[17].entry.input_buf[0].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[17].entry.input_buf[0].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[17].entry.input_buf[0].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[17].entry.input_buf[0].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[17].entry.input_buf[0].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[17].entry.input_buf[0].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[17].entry.input_buf[1].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[17].entry.input_buf[1].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[17].entry.input_buf[1].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[17].entry.input_buf[1].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[17].entry.input_buf[1].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[17].entry.input_buf[1].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[17].entry.input_buf[2].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[17].entry.input_buf[2].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[17].entry.input_buf[2].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[17].entry.input_buf[2].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[17].entry.input_buf[2].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[17].entry.input_buf[2].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[17].entry.input_buf[3].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[17].entry.input_buf[3].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[17].entry.input_buf[3].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[17].entry.input_buf[3].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[17].entry.input_buf[3].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[17].entry.input_buf[3].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[17].entry.input_buf[4].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[17].entry.input_buf[4].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[17].entry.input_buf[4].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[17].entry.input_buf[4].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[17].entry.input_buf[4].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[17].entry.input_buf[4].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[17].entry.input_buf[5].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[17].entry.input_buf[5].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[17].entry.input_buf[5].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[17].entry.input_buf[5].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[17].entry.input_buf[5].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[17].entry.input_buf[5].X ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[17].entry.latch[0]  (.D(\l_fifo.genblk1[17].entry.input_buf[0].X ),
    .GATE(\l_fifo.genblk1[17].entry.empty ),
    .RESET_B(net46),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[16].entry.input_buf[0].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[17].entry.latch[1]  (.D(\l_fifo.genblk1[17].entry.input_buf[1].X ),
    .GATE(\l_fifo.genblk1[17].entry.empty ),
    .RESET_B(net47),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[16].entry.input_buf[1].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[17].entry.latch[2]  (.D(\l_fifo.genblk1[17].entry.input_buf[2].X ),
    .GATE(\l_fifo.genblk1[17].entry.empty ),
    .RESET_B(net48),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[16].entry.input_buf[2].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[17].entry.latch[3]  (.D(\l_fifo.genblk1[17].entry.input_buf[3].X ),
    .GATE(\l_fifo.genblk1[17].entry.empty ),
    .RESET_B(net46),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[16].entry.input_buf[3].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[17].entry.latch[4]  (.D(\l_fifo.genblk1[17].entry.input_buf[4].X ),
    .GATE(\l_fifo.genblk1[17].entry.empty ),
    .RESET_B(net46),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[16].entry.input_buf[4].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[17].entry.latch[5]  (.D(\l_fifo.genblk1[17].entry.input_buf[5].X ),
    .GATE(\l_fifo.genblk1[17].entry.empty ),
    .RESET_B(net46),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[16].entry.input_buf[5].A ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[18].entry.input_buf[0].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[18].entry.input_buf[0].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[18].entry.input_buf[0].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[18].entry.input_buf[0].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[18].entry.input_buf[0].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[18].entry.input_buf[0].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[18].entry.input_buf[1].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[18].entry.input_buf[1].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[18].entry.input_buf[1].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[18].entry.input_buf[1].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[18].entry.input_buf[1].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[18].entry.input_buf[1].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[18].entry.input_buf[2].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[18].entry.input_buf[2].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[18].entry.input_buf[2].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[18].entry.input_buf[2].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[18].entry.input_buf[2].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[18].entry.input_buf[2].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[18].entry.input_buf[3].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[18].entry.input_buf[3].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[18].entry.input_buf[3].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[18].entry.input_buf[3].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[18].entry.input_buf[3].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[18].entry.input_buf[3].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[18].entry.input_buf[4].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[18].entry.input_buf[4].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[18].entry.input_buf[4].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[18].entry.input_buf[4].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[18].entry.input_buf[4].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[18].entry.input_buf[4].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[18].entry.input_buf[5].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[18].entry.input_buf[5].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[18].entry.input_buf[5].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[18].entry.input_buf[5].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[18].entry.input_buf[5].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[18].entry.input_buf[5].X ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[18].entry.latch[0]  (.D(\l_fifo.genblk1[18].entry.input_buf[0].X ),
    .GATE(\l_fifo.genblk1[18].entry.empty ),
    .RESET_B(net46),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[17].entry.input_buf[0].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[18].entry.latch[1]  (.D(\l_fifo.genblk1[18].entry.input_buf[1].X ),
    .GATE(\l_fifo.genblk1[18].entry.empty ),
    .RESET_B(net41),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[17].entry.input_buf[1].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[18].entry.latch[2]  (.D(\l_fifo.genblk1[18].entry.input_buf[2].X ),
    .GATE(\l_fifo.genblk1[18].entry.empty ),
    .RESET_B(net46),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[17].entry.input_buf[2].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[18].entry.latch[3]  (.D(\l_fifo.genblk1[18].entry.input_buf[3].X ),
    .GATE(\l_fifo.genblk1[18].entry.empty ),
    .RESET_B(net47),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[17].entry.input_buf[3].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[18].entry.latch[4]  (.D(\l_fifo.genblk1[18].entry.input_buf[4].X ),
    .GATE(\l_fifo.genblk1[18].entry.empty ),
    .RESET_B(net46),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[17].entry.input_buf[4].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[18].entry.latch[5]  (.D(\l_fifo.genblk1[18].entry.input_buf[5].X ),
    .GATE(\l_fifo.genblk1[18].entry.empty ),
    .RESET_B(net41),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[17].entry.input_buf[5].A ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[19].entry.input_buf[0].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[19].entry.input_buf[0].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[19].entry.input_buf[0].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[19].entry.input_buf[0].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[19].entry.input_buf[0].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[19].entry.input_buf[0].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[19].entry.input_buf[1].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[19].entry.input_buf[1].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[19].entry.input_buf[1].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[19].entry.input_buf[1].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[19].entry.input_buf[1].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[19].entry.input_buf[1].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[19].entry.input_buf[2].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[19].entry.input_buf[2].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[19].entry.input_buf[2].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[19].entry.input_buf[2].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[19].entry.input_buf[2].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[19].entry.input_buf[2].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[19].entry.input_buf[3].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[19].entry.input_buf[3].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[19].entry.input_buf[3].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[19].entry.input_buf[3].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[19].entry.input_buf[3].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[19].entry.input_buf[3].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[19].entry.input_buf[4].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[19].entry.input_buf[4].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[19].entry.input_buf[4].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[19].entry.input_buf[4].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[19].entry.input_buf[4].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[19].entry.input_buf[4].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[19].entry.input_buf[5].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[19].entry.input_buf[5].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[19].entry.input_buf[5].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[19].entry.input_buf[5].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[19].entry.input_buf[5].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[19].entry.input_buf[5].X ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[19].entry.latch[0]  (.D(\l_fifo.genblk1[19].entry.input_buf[0].X ),
    .GATE(\l_fifo.genblk1[19].entry.empty ),
    .RESET_B(net41),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[18].entry.input_buf[0].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[19].entry.latch[1]  (.D(\l_fifo.genblk1[19].entry.input_buf[1].X ),
    .GATE(\l_fifo.genblk1[19].entry.empty ),
    .RESET_B(net39),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[18].entry.input_buf[1].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[19].entry.latch[2]  (.D(\l_fifo.genblk1[19].entry.input_buf[2].X ),
    .GATE(\l_fifo.genblk1[19].entry.empty ),
    .RESET_B(net41),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[18].entry.input_buf[2].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[19].entry.latch[3]  (.D(\l_fifo.genblk1[19].entry.input_buf[3].X ),
    .GATE(\l_fifo.genblk1[19].entry.empty ),
    .RESET_B(net42),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[18].entry.input_buf[3].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[19].entry.latch[4]  (.D(\l_fifo.genblk1[19].entry.input_buf[4].X ),
    .GATE(\l_fifo.genblk1[19].entry.empty ),
    .RESET_B(net41),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[18].entry.input_buf[4].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[19].entry.latch[5]  (.D(\l_fifo.genblk1[19].entry.input_buf[5].X ),
    .GATE(\l_fifo.genblk1[19].entry.empty ),
    .RESET_B(net37),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[18].entry.input_buf[5].A ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[1].entry.input_buf[0].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[1].entry.input_buf[0].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[1].entry.input_buf[0].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[1].entry.input_buf[0].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[1].entry.input_buf[0].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[1].entry.input_buf[0].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[1].entry.input_buf[1].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[1].entry.input_buf[1].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[1].entry.input_buf[1].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[1].entry.input_buf[1].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[1].entry.input_buf[1].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[1].entry.input_buf[1].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[1].entry.input_buf[2].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[1].entry.input_buf[2].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[1].entry.input_buf[2].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[1].entry.input_buf[2].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[1].entry.input_buf[2].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[1].entry.input_buf[2].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[1].entry.input_buf[3].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[1].entry.input_buf[3].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[1].entry.input_buf[3].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[1].entry.input_buf[3].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[1].entry.input_buf[3].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[1].entry.input_buf[3].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[1].entry.input_buf[4].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[1].entry.input_buf[4].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[1].entry.input_buf[4].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[1].entry.input_buf[4].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[1].entry.input_buf[4].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[1].entry.input_buf[4].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[1].entry.input_buf[5].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[1].entry.input_buf[5].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[1].entry.input_buf[5].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[1].entry.input_buf[5].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[1].entry.input_buf[5].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[1].entry.input_buf[5].X ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[1].entry.latch[0]  (.D(\l_fifo.genblk1[1].entry.input_buf[0].X ),
    .GATE(\l_fifo.genblk1[1].entry.empty ),
    .RESET_B(net28),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[0].entry.input_buf[0].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[1].entry.latch[1]  (.D(\l_fifo.genblk1[1].entry.input_buf[1].X ),
    .GATE(\l_fifo.genblk1[1].entry.empty ),
    .RESET_B(net28),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[0].entry.input_buf[1].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[1].entry.latch[2]  (.D(\l_fifo.genblk1[1].entry.input_buf[2].X ),
    .GATE(\l_fifo.genblk1[1].entry.empty ),
    .RESET_B(net28),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[0].entry.input_buf[2].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[1].entry.latch[3]  (.D(\l_fifo.genblk1[1].entry.input_buf[3].X ),
    .GATE(\l_fifo.genblk1[1].entry.empty ),
    .RESET_B(net27),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[0].entry.input_buf[3].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[1].entry.latch[4]  (.D(\l_fifo.genblk1[1].entry.input_buf[4].X ),
    .GATE(\l_fifo.genblk1[1].entry.empty ),
    .RESET_B(net27),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[0].entry.input_buf[4].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[1].entry.latch[5]  (.D(\l_fifo.genblk1[1].entry.input_buf[5].X ),
    .GATE(\l_fifo.genblk1[1].entry.empty ),
    .RESET_B(net27),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[0].entry.input_buf[5].A ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[20].entry.input_buf[0].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[20].entry.input_buf[0].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[20].entry.input_buf[0].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[20].entry.input_buf[0].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[20].entry.input_buf[0].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[20].entry.input_buf[0].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[20].entry.input_buf[1].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[20].entry.input_buf[1].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[20].entry.input_buf[1].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[20].entry.input_buf[1].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[20].entry.input_buf[1].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[20].entry.input_buf[1].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[20].entry.input_buf[2].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[20].entry.input_buf[2].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[20].entry.input_buf[2].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[20].entry.input_buf[2].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[20].entry.input_buf[2].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[20].entry.input_buf[2].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[20].entry.input_buf[3].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[20].entry.input_buf[3].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[20].entry.input_buf[3].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[20].entry.input_buf[3].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[20].entry.input_buf[3].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[20].entry.input_buf[3].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[20].entry.input_buf[4].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[20].entry.input_buf[4].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[20].entry.input_buf[4].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[20].entry.input_buf[4].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[20].entry.input_buf[4].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[20].entry.input_buf[4].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[20].entry.input_buf[5].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[20].entry.input_buf[5].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[20].entry.input_buf[5].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[20].entry.input_buf[5].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[20].entry.input_buf[5].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[20].entry.input_buf[5].X ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[20].entry.latch[0]  (.D(\l_fifo.genblk1[20].entry.input_buf[0].X ),
    .GATE(\l_fifo.genblk1[20].entry.empty ),
    .RESET_B(net39),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[19].entry.input_buf[0].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[20].entry.latch[1]  (.D(\l_fifo.genblk1[20].entry.input_buf[1].X ),
    .GATE(\l_fifo.genblk1[20].entry.empty ),
    .RESET_B(net41),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[19].entry.input_buf[1].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[20].entry.latch[2]  (.D(\l_fifo.genblk1[20].entry.input_buf[2].X ),
    .GATE(\l_fifo.genblk1[20].entry.empty ),
    .RESET_B(net42),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[19].entry.input_buf[2].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[20].entry.latch[3]  (.D(\l_fifo.genblk1[20].entry.input_buf[3].X ),
    .GATE(\l_fifo.genblk1[20].entry.empty ),
    .RESET_B(net41),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[19].entry.input_buf[3].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[20].entry.latch[4]  (.D(\l_fifo.genblk1[20].entry.input_buf[4].X ),
    .GATE(\l_fifo.genblk1[20].entry.empty ),
    .RESET_B(net41),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[19].entry.input_buf[4].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[20].entry.latch[5]  (.D(\l_fifo.genblk1[20].entry.input_buf[5].X ),
    .GATE(\l_fifo.genblk1[20].entry.empty ),
    .RESET_B(net35),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[19].entry.input_buf[5].A ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[21].entry.input_buf[0].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[21].entry.input_buf[0].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[21].entry.input_buf[0].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[21].entry.input_buf[0].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[21].entry.input_buf[0].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[21].entry.input_buf[0].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[21].entry.input_buf[1].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[21].entry.input_buf[1].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[21].entry.input_buf[1].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[21].entry.input_buf[1].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[21].entry.input_buf[1].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[21].entry.input_buf[1].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[21].entry.input_buf[2].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[21].entry.input_buf[2].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[21].entry.input_buf[2].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[21].entry.input_buf[2].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[21].entry.input_buf[2].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[21].entry.input_buf[2].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[21].entry.input_buf[3].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[21].entry.input_buf[3].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[21].entry.input_buf[3].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[21].entry.input_buf[3].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[21].entry.input_buf[3].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[21].entry.input_buf[3].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[21].entry.input_buf[4].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[21].entry.input_buf[4].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[21].entry.input_buf[4].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[21].entry.input_buf[4].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[21].entry.input_buf[4].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[21].entry.input_buf[4].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[21].entry.input_buf[5].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[21].entry.input_buf[5].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[21].entry.input_buf[5].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[21].entry.input_buf[5].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[21].entry.input_buf[5].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[21].entry.input_buf[5].X ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[21].entry.latch[0]  (.D(\l_fifo.genblk1[21].entry.input_buf[0].X ),
    .GATE(\l_fifo.genblk1[21].entry.empty ),
    .RESET_B(net39),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[20].entry.input_buf[0].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[21].entry.latch[1]  (.D(\l_fifo.genblk1[21].entry.input_buf[1].X ),
    .GATE(\l_fifo.genblk1[21].entry.empty ),
    .RESET_B(net40),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[20].entry.input_buf[1].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[21].entry.latch[2]  (.D(\l_fifo.genblk1[21].entry.input_buf[2].X ),
    .GATE(\l_fifo.genblk1[21].entry.empty ),
    .RESET_B(net39),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[20].entry.input_buf[2].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[21].entry.latch[3]  (.D(\l_fifo.genblk1[21].entry.input_buf[3].X ),
    .GATE(\l_fifo.genblk1[21].entry.empty ),
    .RESET_B(net39),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[20].entry.input_buf[3].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[21].entry.latch[4]  (.D(\l_fifo.genblk1[21].entry.input_buf[4].X ),
    .GATE(\l_fifo.genblk1[21].entry.empty ),
    .RESET_B(net39),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[20].entry.input_buf[4].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[21].entry.latch[5]  (.D(\l_fifo.genblk1[21].entry.input_buf[5].X ),
    .GATE(\l_fifo.genblk1[21].entry.empty ),
    .RESET_B(net23),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[20].entry.input_buf[5].A ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[22].entry.input_buf[0].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[22].entry.input_buf[0].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[22].entry.input_buf[0].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[22].entry.input_buf[0].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[22].entry.input_buf[0].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[22].entry.input_buf[0].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[22].entry.input_buf[1].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[22].entry.input_buf[1].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[22].entry.input_buf[1].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[22].entry.input_buf[1].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[22].entry.input_buf[1].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[22].entry.input_buf[1].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[22].entry.input_buf[2].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[22].entry.input_buf[2].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[22].entry.input_buf[2].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[22].entry.input_buf[2].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[22].entry.input_buf[2].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[22].entry.input_buf[2].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[22].entry.input_buf[3].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[22].entry.input_buf[3].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[22].entry.input_buf[3].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[22].entry.input_buf[3].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[22].entry.input_buf[3].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[22].entry.input_buf[3].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[22].entry.input_buf[4].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[22].entry.input_buf[4].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[22].entry.input_buf[4].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[22].entry.input_buf[4].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[22].entry.input_buf[4].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[22].entry.input_buf[4].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[22].entry.input_buf[5].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[22].entry.input_buf[5].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[22].entry.input_buf[5].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[22].entry.input_buf[5].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[22].entry.input_buf[5].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[22].entry.input_buf[5].X ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[22].entry.latch[0]  (.D(\l_fifo.genblk1[22].entry.input_buf[0].X ),
    .GATE(\l_fifo.genblk1[22].entry.empty ),
    .RESET_B(net40),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[21].entry.input_buf[0].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[22].entry.latch[1]  (.D(\l_fifo.genblk1[22].entry.input_buf[1].X ),
    .GATE(\l_fifo.genblk1[22].entry.empty ),
    .RESET_B(net39),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[21].entry.input_buf[1].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[22].entry.latch[2]  (.D(\l_fifo.genblk1[22].entry.input_buf[2].X ),
    .GATE(\l_fifo.genblk1[22].entry.empty ),
    .RESET_B(net39),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[21].entry.input_buf[2].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[22].entry.latch[3]  (.D(\l_fifo.genblk1[22].entry.input_buf[3].X ),
    .GATE(\l_fifo.genblk1[22].entry.empty ),
    .RESET_B(net39),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[21].entry.input_buf[3].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[22].entry.latch[4]  (.D(\l_fifo.genblk1[22].entry.input_buf[4].X ),
    .GATE(\l_fifo.genblk1[22].entry.empty ),
    .RESET_B(net41),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[21].entry.input_buf[4].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[22].entry.latch[5]  (.D(\l_fifo.genblk1[22].entry.input_buf[5].X ),
    .GATE(\l_fifo.genblk1[22].entry.empty ),
    .RESET_B(net20),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[21].entry.input_buf[5].A ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[23].entry.input_buf[0].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[23].entry.input_buf[0].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[23].entry.input_buf[0].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[23].entry.input_buf[0].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[23].entry.input_buf[0].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[23].entry.input_buf[0].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[23].entry.input_buf[1].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[23].entry.input_buf[1].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[23].entry.input_buf[1].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[23].entry.input_buf[1].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[23].entry.input_buf[1].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[23].entry.input_buf[1].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[23].entry.input_buf[2].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[23].entry.input_buf[2].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[23].entry.input_buf[2].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[23].entry.input_buf[2].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[23].entry.input_buf[2].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[23].entry.input_buf[2].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[23].entry.input_buf[3].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[23].entry.input_buf[3].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[23].entry.input_buf[3].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[23].entry.input_buf[3].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[23].entry.input_buf[3].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[23].entry.input_buf[3].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[23].entry.input_buf[4].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[23].entry.input_buf[4].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[23].entry.input_buf[4].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[23].entry.input_buf[4].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[23].entry.input_buf[4].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[23].entry.input_buf[4].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[23].entry.input_buf[5].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[23].entry.input_buf[5].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[23].entry.input_buf[5].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[23].entry.input_buf[5].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[23].entry.input_buf[5].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[23].entry.input_buf[5].X ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[23].entry.latch[0]  (.D(\l_fifo.genblk1[23].entry.input_buf[0].X ),
    .GATE(\l_fifo.genblk1[23].entry.empty ),
    .RESET_B(net40),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[22].entry.input_buf[0].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[23].entry.latch[1]  (.D(\l_fifo.genblk1[23].entry.input_buf[1].X ),
    .GATE(\l_fifo.genblk1[23].entry.empty ),
    .RESET_B(net40),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[22].entry.input_buf[1].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[23].entry.latch[2]  (.D(\l_fifo.genblk1[23].entry.input_buf[2].X ),
    .GATE(\l_fifo.genblk1[23].entry.empty ),
    .RESET_B(net38),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[22].entry.input_buf[2].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[23].entry.latch[3]  (.D(\l_fifo.genblk1[23].entry.input_buf[3].X ),
    .GATE(\l_fifo.genblk1[23].entry.empty ),
    .RESET_B(net19),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[22].entry.input_buf[3].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[23].entry.latch[4]  (.D(\l_fifo.genblk1[23].entry.input_buf[4].X ),
    .GATE(\l_fifo.genblk1[23].entry.empty ),
    .RESET_B(net41),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[22].entry.input_buf[4].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[23].entry.latch[5]  (.D(\l_fifo.genblk1[23].entry.input_buf[5].X ),
    .GATE(\l_fifo.genblk1[23].entry.empty ),
    .RESET_B(net39),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[22].entry.input_buf[5].A ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[24].entry.input_buf[0].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[24].entry.input_buf[0].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[24].entry.input_buf[0].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[24].entry.input_buf[0].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[24].entry.input_buf[0].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[24].entry.input_buf[0].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[24].entry.input_buf[1].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[24].entry.input_buf[1].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[24].entry.input_buf[1].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[24].entry.input_buf[1].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[24].entry.input_buf[1].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[24].entry.input_buf[1].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[24].entry.input_buf[2].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[24].entry.input_buf[2].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[24].entry.input_buf[2].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[24].entry.input_buf[2].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[24].entry.input_buf[2].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[24].entry.input_buf[2].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[24].entry.input_buf[3].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[24].entry.input_buf[3].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[24].entry.input_buf[3].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[24].entry.input_buf[3].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[24].entry.input_buf[3].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[24].entry.input_buf[3].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[24].entry.input_buf[4].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[24].entry.input_buf[4].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[24].entry.input_buf[4].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[24].entry.input_buf[4].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[24].entry.input_buf[4].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[24].entry.input_buf[4].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[24].entry.input_buf[5].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[24].entry.input_buf[5].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[24].entry.input_buf[5].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[24].entry.input_buf[5].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[24].entry.input_buf[5].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[24].entry.input_buf[5].X ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[24].entry.latch[0]  (.D(\l_fifo.genblk1[24].entry.input_buf[0].X ),
    .GATE(\l_fifo.genblk1[24].entry.empty ),
    .RESET_B(net23),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[23].entry.input_buf[0].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[24].entry.latch[1]  (.D(\l_fifo.genblk1[24].entry.input_buf[1].X ),
    .GATE(\l_fifo.genblk1[24].entry.empty ),
    .RESET_B(net40),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[23].entry.input_buf[1].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[24].entry.latch[2]  (.D(\l_fifo.genblk1[24].entry.input_buf[2].X ),
    .GATE(\l_fifo.genblk1[24].entry.empty ),
    .RESET_B(net23),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[23].entry.input_buf[2].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[24].entry.latch[3]  (.D(\l_fifo.genblk1[24].entry.input_buf[3].X ),
    .GATE(\l_fifo.genblk1[24].entry.empty ),
    .RESET_B(net22),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[23].entry.input_buf[3].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[24].entry.latch[4]  (.D(\l_fifo.genblk1[24].entry.input_buf[4].X ),
    .GATE(\l_fifo.genblk1[24].entry.empty ),
    .RESET_B(net23),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[23].entry.input_buf[4].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[24].entry.latch[5]  (.D(\l_fifo.genblk1[24].entry.input_buf[5].X ),
    .GATE(\l_fifo.genblk1[24].entry.empty ),
    .RESET_B(net23),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[23].entry.input_buf[5].A ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[25].entry.input_buf[0].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[25].entry.input_buf[0].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[25].entry.input_buf[0].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[25].entry.input_buf[0].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[25].entry.input_buf[0].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[25].entry.input_buf[0].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[25].entry.input_buf[1].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[25].entry.input_buf[1].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[25].entry.input_buf[1].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[25].entry.input_buf[1].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[25].entry.input_buf[1].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[25].entry.input_buf[1].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[25].entry.input_buf[2].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[25].entry.input_buf[2].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[25].entry.input_buf[2].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[25].entry.input_buf[2].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[25].entry.input_buf[2].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[25].entry.input_buf[2].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[25].entry.input_buf[3].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[25].entry.input_buf[3].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[25].entry.input_buf[3].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[25].entry.input_buf[3].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[25].entry.input_buf[3].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[25].entry.input_buf[3].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[25].entry.input_buf[4].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[25].entry.input_buf[4].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[25].entry.input_buf[4].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[25].entry.input_buf[4].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[25].entry.input_buf[4].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[25].entry.input_buf[4].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[25].entry.input_buf[5].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[25].entry.input_buf[5].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[25].entry.input_buf[5].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[25].entry.input_buf[5].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[25].entry.input_buf[5].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[25].entry.input_buf[5].X ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[25].entry.latch[0]  (.D(\l_fifo.genblk1[25].entry.input_buf[0].X ),
    .GATE(\l_fifo.genblk1[25].entry.empty ),
    .RESET_B(net24),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[24].entry.input_buf[0].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[25].entry.latch[1]  (.D(\l_fifo.genblk1[25].entry.input_buf[1].X ),
    .GATE(\l_fifo.genblk1[25].entry.empty ),
    .RESET_B(net24),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[24].entry.input_buf[1].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[25].entry.latch[2]  (.D(\l_fifo.genblk1[25].entry.input_buf[2].X ),
    .GATE(\l_fifo.genblk1[25].entry.empty ),
    .RESET_B(net23),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[24].entry.input_buf[2].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[25].entry.latch[3]  (.D(\l_fifo.genblk1[25].entry.input_buf[3].X ),
    .GATE(\l_fifo.genblk1[25].entry.empty ),
    .RESET_B(net23),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[24].entry.input_buf[3].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[25].entry.latch[4]  (.D(\l_fifo.genblk1[25].entry.input_buf[4].X ),
    .GATE(\l_fifo.genblk1[25].entry.empty ),
    .RESET_B(net23),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[24].entry.input_buf[4].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[25].entry.latch[5]  (.D(\l_fifo.genblk1[25].entry.input_buf[5].X ),
    .GATE(\l_fifo.genblk1[25].entry.empty ),
    .RESET_B(net20),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[24].entry.input_buf[5].A ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[26].entry.input_buf[0].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[26].entry.input_buf[0].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[26].entry.input_buf[0].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[26].entry.input_buf[0].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[26].entry.input_buf[0].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[26].entry.input_buf[0].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[26].entry.input_buf[1].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[26].entry.input_buf[1].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[26].entry.input_buf[1].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[26].entry.input_buf[1].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[26].entry.input_buf[1].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[26].entry.input_buf[1].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[26].entry.input_buf[2].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[26].entry.input_buf[2].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[26].entry.input_buf[2].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[26].entry.input_buf[2].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[26].entry.input_buf[2].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[26].entry.input_buf[2].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[26].entry.input_buf[3].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[26].entry.input_buf[3].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[26].entry.input_buf[3].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[26].entry.input_buf[3].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[26].entry.input_buf[3].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[26].entry.input_buf[3].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[26].entry.input_buf[4].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[26].entry.input_buf[4].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[26].entry.input_buf[4].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[26].entry.input_buf[4].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[26].entry.input_buf[4].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[26].entry.input_buf[4].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[26].entry.input_buf[5].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[26].entry.input_buf[5].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[26].entry.input_buf[5].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[26].entry.input_buf[5].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[26].entry.input_buf[5].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[26].entry.input_buf[5].X ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[26].entry.latch[0]  (.D(\l_fifo.genblk1[26].entry.input_buf[0].X ),
    .GATE(\l_fifo.genblk1[26].entry.empty ),
    .RESET_B(net22),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[25].entry.input_buf[0].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[26].entry.latch[1]  (.D(\l_fifo.genblk1[26].entry.input_buf[1].X ),
    .GATE(\l_fifo.genblk1[26].entry.empty ),
    .RESET_B(net24),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[25].entry.input_buf[1].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[26].entry.latch[2]  (.D(\l_fifo.genblk1[26].entry.input_buf[2].X ),
    .GATE(\l_fifo.genblk1[26].entry.empty ),
    .RESET_B(net24),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[25].entry.input_buf[2].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[26].entry.latch[3]  (.D(\l_fifo.genblk1[26].entry.input_buf[3].X ),
    .GATE(\l_fifo.genblk1[26].entry.empty ),
    .RESET_B(net15),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[25].entry.input_buf[3].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[26].entry.latch[4]  (.D(\l_fifo.genblk1[26].entry.input_buf[4].X ),
    .GATE(\l_fifo.genblk1[26].entry.empty ),
    .RESET_B(net15),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[25].entry.input_buf[4].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[26].entry.latch[5]  (.D(\l_fifo.genblk1[26].entry.input_buf[5].X ),
    .GATE(\l_fifo.genblk1[26].entry.empty ),
    .RESET_B(net23),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[25].entry.input_buf[5].A ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[27].entry.input_buf[0].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[27].entry.input_buf[0].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[27].entry.input_buf[0].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[27].entry.input_buf[0].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[27].entry.input_buf[0].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[27].entry.input_buf[0].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[27].entry.input_buf[1].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[27].entry.input_buf[1].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[27].entry.input_buf[1].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[27].entry.input_buf[1].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[27].entry.input_buf[1].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[27].entry.input_buf[1].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[27].entry.input_buf[2].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[27].entry.input_buf[2].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[27].entry.input_buf[2].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[27].entry.input_buf[2].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[27].entry.input_buf[2].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[27].entry.input_buf[2].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[27].entry.input_buf[3].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[27].entry.input_buf[3].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[27].entry.input_buf[3].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[27].entry.input_buf[3].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[27].entry.input_buf[3].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[27].entry.input_buf[3].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[27].entry.input_buf[4].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[27].entry.input_buf[4].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[27].entry.input_buf[4].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[27].entry.input_buf[4].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[27].entry.input_buf[4].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[27].entry.input_buf[4].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[27].entry.input_buf[5].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[27].entry.input_buf[5].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[27].entry.input_buf[5].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[27].entry.input_buf[5].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[27].entry.input_buf[5].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[27].entry.input_buf[5].X ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[27].entry.latch[0]  (.D(\l_fifo.genblk1[27].entry.input_buf[0].X ),
    .GATE(\l_fifo.genblk1[27].entry.empty ),
    .RESET_B(net22),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[26].entry.input_buf[0].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[27].entry.latch[1]  (.D(\l_fifo.genblk1[27].entry.input_buf[1].X ),
    .GATE(\l_fifo.genblk1[27].entry.empty ),
    .RESET_B(net22),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[26].entry.input_buf[1].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[27].entry.latch[2]  (.D(\l_fifo.genblk1[27].entry.input_buf[2].X ),
    .GATE(\l_fifo.genblk1[27].entry.empty ),
    .RESET_B(net22),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[26].entry.input_buf[2].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[27].entry.latch[3]  (.D(\l_fifo.genblk1[27].entry.input_buf[3].X ),
    .GATE(\l_fifo.genblk1[27].entry.empty ),
    .RESET_B(net23),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[26].entry.input_buf[3].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[27].entry.latch[4]  (.D(\l_fifo.genblk1[27].entry.input_buf[4].X ),
    .GATE(\l_fifo.genblk1[27].entry.empty ),
    .RESET_B(net22),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[26].entry.input_buf[4].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[27].entry.latch[5]  (.D(\l_fifo.genblk1[27].entry.input_buf[5].X ),
    .GATE(\l_fifo.genblk1[27].entry.empty ),
    .RESET_B(net24),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[26].entry.input_buf[5].A ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[28].entry.input_buf[0].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[28].entry.input_buf[0].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[28].entry.input_buf[0].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[28].entry.input_buf[0].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[28].entry.input_buf[0].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[28].entry.input_buf[0].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[28].entry.input_buf[1].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[28].entry.input_buf[1].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[28].entry.input_buf[1].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[28].entry.input_buf[1].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[28].entry.input_buf[1].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[28].entry.input_buf[1].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[28].entry.input_buf[2].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[28].entry.input_buf[2].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[28].entry.input_buf[2].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[28].entry.input_buf[2].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[28].entry.input_buf[2].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[28].entry.input_buf[2].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[28].entry.input_buf[3].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[28].entry.input_buf[3].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[28].entry.input_buf[3].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[28].entry.input_buf[3].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[28].entry.input_buf[3].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[28].entry.input_buf[3].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[28].entry.input_buf[4].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[28].entry.input_buf[4].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[28].entry.input_buf[4].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[28].entry.input_buf[4].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[28].entry.input_buf[4].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[28].entry.input_buf[4].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[28].entry.input_buf[5].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[28].entry.input_buf[5].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[28].entry.input_buf[5].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[28].entry.input_buf[5].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[28].entry.input_buf[5].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[28].entry.input_buf[5].X ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[28].entry.latch[0]  (.D(\l_fifo.genblk1[28].entry.input_buf[0].X ),
    .GATE(\l_fifo.genblk1[28].entry.empty ),
    .RESET_B(net22),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[27].entry.input_buf[0].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[28].entry.latch[1]  (.D(\l_fifo.genblk1[28].entry.input_buf[1].X ),
    .GATE(\l_fifo.genblk1[28].entry.empty ),
    .RESET_B(net24),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[27].entry.input_buf[1].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[28].entry.latch[2]  (.D(\l_fifo.genblk1[28].entry.input_buf[2].X ),
    .GATE(\l_fifo.genblk1[28].entry.empty ),
    .RESET_B(net15),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[27].entry.input_buf[2].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[28].entry.latch[3]  (.D(\l_fifo.genblk1[28].entry.input_buf[3].X ),
    .GATE(\l_fifo.genblk1[28].entry.empty ),
    .RESET_B(net22),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[27].entry.input_buf[3].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[28].entry.latch[4]  (.D(\l_fifo.genblk1[28].entry.input_buf[4].X ),
    .GATE(\l_fifo.genblk1[28].entry.empty ),
    .RESET_B(net15),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[27].entry.input_buf[4].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[28].entry.latch[5]  (.D(\l_fifo.genblk1[28].entry.input_buf[5].X ),
    .GATE(\l_fifo.genblk1[28].entry.empty ),
    .RESET_B(net22),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[27].entry.input_buf[5].A ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[29].entry.input_buf[0].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[29].entry.input_buf[0].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[29].entry.input_buf[0].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[29].entry.input_buf[0].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[29].entry.input_buf[0].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[29].entry.input_buf[0].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[29].entry.input_buf[1].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[29].entry.input_buf[1].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[29].entry.input_buf[1].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[29].entry.input_buf[1].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[29].entry.input_buf[1].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[29].entry.input_buf[1].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[29].entry.input_buf[2].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[29].entry.input_buf[2].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[29].entry.input_buf[2].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[29].entry.input_buf[2].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[29].entry.input_buf[2].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[29].entry.input_buf[2].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[29].entry.input_buf[3].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[29].entry.input_buf[3].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[29].entry.input_buf[3].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[29].entry.input_buf[3].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[29].entry.input_buf[3].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[29].entry.input_buf[3].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[29].entry.input_buf[4].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[29].entry.input_buf[4].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[29].entry.input_buf[4].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[29].entry.input_buf[4].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[29].entry.input_buf[4].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[29].entry.input_buf[4].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[29].entry.input_buf[5].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[29].entry.input_buf[5].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[29].entry.input_buf[5].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[29].entry.input_buf[5].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[29].entry.input_buf[5].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[29].entry.input_buf[5].X ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[29].entry.latch[0]  (.D(\l_fifo.genblk1[29].entry.input_buf[0].X ),
    .GATE(\l_fifo.genblk1[29].entry.empty ),
    .RESET_B(net16),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[28].entry.input_buf[0].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[29].entry.latch[1]  (.D(\l_fifo.genblk1[29].entry.input_buf[1].X ),
    .GATE(\l_fifo.genblk1[29].entry.empty ),
    .RESET_B(net22),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[28].entry.input_buf[1].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[29].entry.latch[2]  (.D(\l_fifo.genblk1[29].entry.input_buf[2].X ),
    .GATE(\l_fifo.genblk1[29].entry.empty ),
    .RESET_B(net15),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[28].entry.input_buf[2].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[29].entry.latch[3]  (.D(\l_fifo.genblk1[29].entry.input_buf[3].X ),
    .GATE(\l_fifo.genblk1[29].entry.empty ),
    .RESET_B(net15),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[28].entry.input_buf[3].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[29].entry.latch[4]  (.D(\l_fifo.genblk1[29].entry.input_buf[4].X ),
    .GATE(\l_fifo.genblk1[29].entry.empty ),
    .RESET_B(net15),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[28].entry.input_buf[4].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[29].entry.latch[5]  (.D(\l_fifo.genblk1[29].entry.input_buf[5].X ),
    .GATE(\l_fifo.genblk1[29].entry.empty ),
    .RESET_B(net16),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[28].entry.input_buf[5].A ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[2].entry.input_buf[0].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[2].entry.input_buf[0].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[2].entry.input_buf[0].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[2].entry.input_buf[0].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[2].entry.input_buf[0].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[2].entry.input_buf[0].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[2].entry.input_buf[1].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[2].entry.input_buf[1].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[2].entry.input_buf[1].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[2].entry.input_buf[1].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[2].entry.input_buf[1].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[2].entry.input_buf[1].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[2].entry.input_buf[2].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[2].entry.input_buf[2].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[2].entry.input_buf[2].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[2].entry.input_buf[2].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[2].entry.input_buf[2].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[2].entry.input_buf[2].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[2].entry.input_buf[3].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[2].entry.input_buf[3].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[2].entry.input_buf[3].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[2].entry.input_buf[3].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[2].entry.input_buf[3].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[2].entry.input_buf[3].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[2].entry.input_buf[4].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[2].entry.input_buf[4].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[2].entry.input_buf[4].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[2].entry.input_buf[4].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[2].entry.input_buf[4].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[2].entry.input_buf[4].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[2].entry.input_buf[5].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[2].entry.input_buf[5].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[2].entry.input_buf[5].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[2].entry.input_buf[5].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[2].entry.input_buf[5].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[2].entry.input_buf[5].X ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[2].entry.latch[0]  (.D(\l_fifo.genblk1[2].entry.input_buf[0].X ),
    .GATE(\l_fifo.genblk1[2].entry.empty ),
    .RESET_B(net28),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[1].entry.input_buf[0].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[2].entry.latch[1]  (.D(\l_fifo.genblk1[2].entry.input_buf[1].X ),
    .GATE(\l_fifo.genblk1[2].entry.empty ),
    .RESET_B(net29),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[1].entry.input_buf[1].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[2].entry.latch[2]  (.D(\l_fifo.genblk1[2].entry.input_buf[2].X ),
    .GATE(\l_fifo.genblk1[2].entry.empty ),
    .RESET_B(net28),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[1].entry.input_buf[2].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[2].entry.latch[3]  (.D(\l_fifo.genblk1[2].entry.input_buf[3].X ),
    .GATE(\l_fifo.genblk1[2].entry.empty ),
    .RESET_B(net30),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[1].entry.input_buf[3].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[2].entry.latch[4]  (.D(\l_fifo.genblk1[2].entry.input_buf[4].X ),
    .GATE(\l_fifo.genblk1[2].entry.empty ),
    .RESET_B(net29),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[1].entry.input_buf[4].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[2].entry.latch[5]  (.D(\l_fifo.genblk1[2].entry.input_buf[5].X ),
    .GATE(\l_fifo.genblk1[2].entry.empty ),
    .RESET_B(net28),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[1].entry.input_buf[5].A ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[30].entry.input_buf[0].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[30].entry.input_buf[0].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[30].entry.input_buf[0].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[30].entry.input_buf[0].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[30].entry.input_buf[0].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[30].entry.input_buf[0].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[30].entry.input_buf[1].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[30].entry.input_buf[1].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[30].entry.input_buf[1].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[30].entry.input_buf[1].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[30].entry.input_buf[1].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[30].entry.input_buf[1].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[30].entry.input_buf[2].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[30].entry.input_buf[2].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[30].entry.input_buf[2].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[30].entry.input_buf[2].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[30].entry.input_buf[2].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[30].entry.input_buf[2].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[30].entry.input_buf[3].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[30].entry.input_buf[3].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[30].entry.input_buf[3].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[30].entry.input_buf[3].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[30].entry.input_buf[3].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[30].entry.input_buf[3].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[30].entry.input_buf[4].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[30].entry.input_buf[4].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[30].entry.input_buf[4].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[30].entry.input_buf[4].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[30].entry.input_buf[4].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[30].entry.input_buf[4].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[30].entry.input_buf[5].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[30].entry.input_buf[5].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[30].entry.input_buf[5].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[30].entry.input_buf[5].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[30].entry.input_buf[5].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[30].entry.input_buf[5].X ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[30].entry.latch[0]  (.D(\l_fifo.genblk1[30].entry.input_buf[0].X ),
    .GATE(\l_fifo.genblk1[30].entry.empty ),
    .RESET_B(net17),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[29].entry.input_buf[0].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[30].entry.latch[1]  (.D(\l_fifo.genblk1[30].entry.input_buf[1].X ),
    .GATE(\l_fifo.genblk1[30].entry.empty ),
    .RESET_B(net16),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[29].entry.input_buf[1].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[30].entry.latch[2]  (.D(\l_fifo.genblk1[30].entry.input_buf[2].X ),
    .GATE(\l_fifo.genblk1[30].entry.empty ),
    .RESET_B(net14),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[29].entry.input_buf[2].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[30].entry.latch[3]  (.D(\l_fifo.genblk1[30].entry.input_buf[3].X ),
    .GATE(\l_fifo.genblk1[30].entry.empty ),
    .RESET_B(net16),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[29].entry.input_buf[3].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[30].entry.latch[4]  (.D(\l_fifo.genblk1[30].entry.input_buf[4].X ),
    .GATE(\l_fifo.genblk1[30].entry.empty ),
    .RESET_B(net17),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[29].entry.input_buf[4].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[30].entry.latch[5]  (.D(\l_fifo.genblk1[30].entry.input_buf[5].X ),
    .GATE(\l_fifo.genblk1[30].entry.empty ),
    .RESET_B(net16),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[29].entry.input_buf[5].A ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[31].entry.input_buf[0].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[31].entry.input_buf[0].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[31].entry.input_buf[0].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[31].entry.input_buf[0].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[31].entry.input_buf[0].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[31].entry.input_buf[0].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[31].entry.input_buf[1].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[31].entry.input_buf[1].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[31].entry.input_buf[1].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[31].entry.input_buf[1].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[31].entry.input_buf[1].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[31].entry.input_buf[1].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[31].entry.input_buf[2].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[31].entry.input_buf[2].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[31].entry.input_buf[2].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[31].entry.input_buf[2].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[31].entry.input_buf[2].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[31].entry.input_buf[2].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[31].entry.input_buf[3].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[31].entry.input_buf[3].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[31].entry.input_buf[3].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[31].entry.input_buf[3].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[31].entry.input_buf[3].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[31].entry.input_buf[3].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[31].entry.input_buf[4].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[31].entry.input_buf[4].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[31].entry.input_buf[4].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[31].entry.input_buf[4].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[31].entry.input_buf[4].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[31].entry.input_buf[4].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[31].entry.input_buf[5].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[31].entry.input_buf[5].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[31].entry.input_buf[5].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[31].entry.input_buf[5].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[31].entry.input_buf[5].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[31].entry.input_buf[5].X ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[31].entry.latch[0]  (.D(\l_fifo.genblk1[31].entry.input_buf[0].X ),
    .GATE(\l_fifo.genblk1[31].entry.empty ),
    .RESET_B(net14),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[30].entry.input_buf[0].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[31].entry.latch[1]  (.D(\l_fifo.genblk1[31].entry.input_buf[1].X ),
    .GATE(\l_fifo.genblk1[31].entry.empty ),
    .RESET_B(net16),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[30].entry.input_buf[1].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[31].entry.latch[2]  (.D(\l_fifo.genblk1[31].entry.input_buf[2].X ),
    .GATE(\l_fifo.genblk1[31].entry.empty ),
    .RESET_B(net14),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[30].entry.input_buf[2].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[31].entry.latch[3]  (.D(\l_fifo.genblk1[31].entry.input_buf[3].X ),
    .GATE(\l_fifo.genblk1[31].entry.empty ),
    .RESET_B(net14),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[30].entry.input_buf[3].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[31].entry.latch[4]  (.D(\l_fifo.genblk1[31].entry.input_buf[4].X ),
    .GATE(\l_fifo.genblk1[31].entry.empty ),
    .RESET_B(net14),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[30].entry.input_buf[4].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[31].entry.latch[5]  (.D(\l_fifo.genblk1[31].entry.input_buf[5].X ),
    .GATE(\l_fifo.genblk1[31].entry.empty ),
    .RESET_B(net14),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[30].entry.input_buf[5].A ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[32].entry.input_buf[0].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[32].entry.input_buf[0].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[32].entry.input_buf[0].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[32].entry.input_buf[0].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[32].entry.input_buf[0].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[32].entry.input_buf[0].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[32].entry.input_buf[1].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[32].entry.input_buf[1].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[32].entry.input_buf[1].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[32].entry.input_buf[1].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[32].entry.input_buf[1].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[32].entry.input_buf[1].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[32].entry.input_buf[2].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[32].entry.input_buf[2].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[32].entry.input_buf[2].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[32].entry.input_buf[2].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[32].entry.input_buf[2].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[32].entry.input_buf[2].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[32].entry.input_buf[3].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[32].entry.input_buf[3].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[32].entry.input_buf[3].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[32].entry.input_buf[3].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[32].entry.input_buf[3].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[32].entry.input_buf[3].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[32].entry.input_buf[4].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[32].entry.input_buf[4].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[32].entry.input_buf[4].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[32].entry.input_buf[4].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[32].entry.input_buf[4].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[32].entry.input_buf[4].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[32].entry.input_buf[5].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[32].entry.input_buf[5].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[32].entry.input_buf[5].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[32].entry.input_buf[5].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[32].entry.input_buf[5].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[32].entry.input_buf[5].X ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[32].entry.latch[0]  (.D(\l_fifo.genblk1[32].entry.input_buf[0].X ),
    .GATE(\l_fifo.genblk1[32].entry.empty ),
    .RESET_B(net14),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[31].entry.input_buf[0].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[32].entry.latch[1]  (.D(\l_fifo.genblk1[32].entry.input_buf[1].X ),
    .GATE(\l_fifo.genblk1[32].entry.empty ),
    .RESET_B(net14),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[31].entry.input_buf[1].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[32].entry.latch[2]  (.D(\l_fifo.genblk1[32].entry.input_buf[2].X ),
    .GATE(\l_fifo.genblk1[32].entry.empty ),
    .RESET_B(net14),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[31].entry.input_buf[2].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[32].entry.latch[3]  (.D(\l_fifo.genblk1[32].entry.input_buf[3].X ),
    .GATE(\l_fifo.genblk1[32].entry.empty ),
    .RESET_B(net10),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[31].entry.input_buf[3].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[32].entry.latch[4]  (.D(\l_fifo.genblk1[32].entry.input_buf[4].X ),
    .GATE(\l_fifo.genblk1[32].entry.empty ),
    .RESET_B(net13),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[31].entry.input_buf[4].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[32].entry.latch[5]  (.D(\l_fifo.genblk1[32].entry.input_buf[5].X ),
    .GATE(\l_fifo.genblk1[32].entry.empty ),
    .RESET_B(net10),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[31].entry.input_buf[5].A ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[33].entry.input_buf[0].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[33].entry.input_buf[0].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[33].entry.input_buf[0].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[33].entry.input_buf[0].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[33].entry.input_buf[0].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[33].entry.input_buf[0].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[33].entry.input_buf[1].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[33].entry.input_buf[1].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[33].entry.input_buf[1].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[33].entry.input_buf[1].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[33].entry.input_buf[1].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[33].entry.input_buf[1].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[33].entry.input_buf[2].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[33].entry.input_buf[2].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[33].entry.input_buf[2].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[33].entry.input_buf[2].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[33].entry.input_buf[2].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[33].entry.input_buf[2].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[33].entry.input_buf[3].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[33].entry.input_buf[3].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[33].entry.input_buf[3].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[33].entry.input_buf[3].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[33].entry.input_buf[3].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[33].entry.input_buf[3].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[33].entry.input_buf[4].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[33].entry.input_buf[4].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[33].entry.input_buf[4].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[33].entry.input_buf[4].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[33].entry.input_buf[4].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[33].entry.input_buf[4].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[33].entry.input_buf[5].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[33].entry.input_buf[5].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[33].entry.input_buf[5].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[33].entry.input_buf[5].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[33].entry.input_buf[5].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[33].entry.input_buf[5].X ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[33].entry.latch[0]  (.D(\l_fifo.genblk1[33].entry.input_buf[0].X ),
    .GATE(\l_fifo.genblk1[33].entry.empty ),
    .RESET_B(net15),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[32].entry.input_buf[0].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[33].entry.latch[1]  (.D(\l_fifo.genblk1[33].entry.input_buf[1].X ),
    .GATE(\l_fifo.genblk1[33].entry.empty ),
    .RESET_B(net15),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[32].entry.input_buf[1].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[33].entry.latch[2]  (.D(\l_fifo.genblk1[33].entry.input_buf[2].X ),
    .GATE(\l_fifo.genblk1[33].entry.empty ),
    .RESET_B(net14),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[32].entry.input_buf[2].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[33].entry.latch[3]  (.D(\l_fifo.genblk1[33].entry.input_buf[3].X ),
    .GATE(\l_fifo.genblk1[33].entry.empty ),
    .RESET_B(net11),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[32].entry.input_buf[3].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[33].entry.latch[4]  (.D(\l_fifo.genblk1[33].entry.input_buf[4].X ),
    .GATE(\l_fifo.genblk1[33].entry.empty ),
    .RESET_B(net11),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[32].entry.input_buf[4].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[33].entry.latch[5]  (.D(\l_fifo.genblk1[33].entry.input_buf[5].X ),
    .GATE(\l_fifo.genblk1[33].entry.empty ),
    .RESET_B(net12),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[32].entry.input_buf[5].A ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[34].entry.input_buf[0].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[34].entry.input_buf[0].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[34].entry.input_buf[0].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[34].entry.input_buf[0].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[34].entry.input_buf[0].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[34].entry.input_buf[0].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[34].entry.input_buf[1].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[34].entry.input_buf[1].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[34].entry.input_buf[1].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[34].entry.input_buf[1].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[34].entry.input_buf[1].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[34].entry.input_buf[1].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[34].entry.input_buf[2].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[34].entry.input_buf[2].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[34].entry.input_buf[2].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[34].entry.input_buf[2].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[34].entry.input_buf[2].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[34].entry.input_buf[2].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[34].entry.input_buf[3].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[34].entry.input_buf[3].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[34].entry.input_buf[3].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[34].entry.input_buf[3].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[34].entry.input_buf[3].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[34].entry.input_buf[3].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[34].entry.input_buf[4].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[34].entry.input_buf[4].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[34].entry.input_buf[4].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[34].entry.input_buf[4].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[34].entry.input_buf[4].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[34].entry.input_buf[4].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[34].entry.input_buf[5].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[34].entry.input_buf[5].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[34].entry.input_buf[5].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[34].entry.input_buf[5].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[34].entry.input_buf[5].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[34].entry.input_buf[5].X ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[34].entry.latch[0]  (.D(\l_fifo.genblk1[34].entry.input_buf[0].X ),
    .GATE(\l_fifo.genblk1[34].entry.empty ),
    .RESET_B(net13),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[33].entry.input_buf[0].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[34].entry.latch[1]  (.D(\l_fifo.genblk1[34].entry.input_buf[1].X ),
    .GATE(\l_fifo.genblk1[34].entry.empty ),
    .RESET_B(net10),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[33].entry.input_buf[1].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[34].entry.latch[2]  (.D(\l_fifo.genblk1[34].entry.input_buf[2].X ),
    .GATE(\l_fifo.genblk1[34].entry.empty ),
    .RESET_B(net15),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[33].entry.input_buf[2].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[34].entry.latch[3]  (.D(\l_fifo.genblk1[34].entry.input_buf[3].X ),
    .GATE(\l_fifo.genblk1[34].entry.empty ),
    .RESET_B(net18),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[33].entry.input_buf[3].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[34].entry.latch[4]  (.D(\l_fifo.genblk1[34].entry.input_buf[4].X ),
    .GATE(\l_fifo.genblk1[34].entry.empty ),
    .RESET_B(net12),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[33].entry.input_buf[4].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[34].entry.latch[5]  (.D(\l_fifo.genblk1[34].entry.input_buf[5].X ),
    .GATE(\l_fifo.genblk1[34].entry.empty ),
    .RESET_B(net11),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[33].entry.input_buf[5].A ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[35].entry.input_buf[0].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[35].entry.input_buf[0].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[35].entry.input_buf[0].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[35].entry.input_buf[0].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[35].entry.input_buf[0].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[35].entry.input_buf[0].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[35].entry.input_buf[1].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[35].entry.input_buf[1].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[35].entry.input_buf[1].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[35].entry.input_buf[1].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[35].entry.input_buf[1].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[35].entry.input_buf[1].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[35].entry.input_buf[2].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[35].entry.input_buf[2].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[35].entry.input_buf[2].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[35].entry.input_buf[2].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[35].entry.input_buf[2].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[35].entry.input_buf[2].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[35].entry.input_buf[3].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[35].entry.input_buf[3].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[35].entry.input_buf[3].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[35].entry.input_buf[3].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[35].entry.input_buf[3].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[35].entry.input_buf[3].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[35].entry.input_buf[4].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[35].entry.input_buf[4].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[35].entry.input_buf[4].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[35].entry.input_buf[4].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[35].entry.input_buf[4].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[35].entry.input_buf[4].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[35].entry.input_buf[5].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[35].entry.input_buf[5].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[35].entry.input_buf[5].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[35].entry.input_buf[5].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[35].entry.input_buf[5].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[35].entry.input_buf[5].X ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[35].entry.latch[0]  (.D(\l_fifo.genblk1[35].entry.input_buf[0].X ),
    .GATE(\l_fifo.genblk1[35].entry.empty ),
    .RESET_B(net10),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[34].entry.input_buf[0].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[35].entry.latch[1]  (.D(\l_fifo.genblk1[35].entry.input_buf[1].X ),
    .GATE(\l_fifo.genblk1[35].entry.empty ),
    .RESET_B(net10),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[34].entry.input_buf[1].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[35].entry.latch[2]  (.D(\l_fifo.genblk1[35].entry.input_buf[2].X ),
    .GATE(\l_fifo.genblk1[35].entry.empty ),
    .RESET_B(net12),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[34].entry.input_buf[2].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[35].entry.latch[3]  (.D(\l_fifo.genblk1[35].entry.input_buf[3].X ),
    .GATE(\l_fifo.genblk1[35].entry.empty ),
    .RESET_B(net21),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[34].entry.input_buf[3].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[35].entry.latch[4]  (.D(\l_fifo.genblk1[35].entry.input_buf[4].X ),
    .GATE(\l_fifo.genblk1[35].entry.empty ),
    .RESET_B(net10),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[34].entry.input_buf[4].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[35].entry.latch[5]  (.D(\l_fifo.genblk1[35].entry.input_buf[5].X ),
    .GATE(\l_fifo.genblk1[35].entry.empty ),
    .RESET_B(net11),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[34].entry.input_buf[5].A ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[36].entry.input_buf[0].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[36].entry.input_buf[0].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[36].entry.input_buf[0].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[36].entry.input_buf[0].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[36].entry.input_buf[0].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[36].entry.input_buf[0].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[36].entry.input_buf[1].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[36].entry.input_buf[1].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[36].entry.input_buf[1].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[36].entry.input_buf[1].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[36].entry.input_buf[1].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[36].entry.input_buf[1].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[36].entry.input_buf[2].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[36].entry.input_buf[2].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[36].entry.input_buf[2].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[36].entry.input_buf[2].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[36].entry.input_buf[2].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[36].entry.input_buf[2].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[36].entry.input_buf[3].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[36].entry.input_buf[3].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[36].entry.input_buf[3].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[36].entry.input_buf[3].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[36].entry.input_buf[3].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[36].entry.input_buf[3].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[36].entry.input_buf[4].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[36].entry.input_buf[4].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[36].entry.input_buf[4].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[36].entry.input_buf[4].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[36].entry.input_buf[4].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[36].entry.input_buf[4].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[36].entry.input_buf[5].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[36].entry.input_buf[5].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[36].entry.input_buf[5].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[36].entry.input_buf[5].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[36].entry.input_buf[5].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[36].entry.input_buf[5].X ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[36].entry.latch[0]  (.D(\l_fifo.genblk1[36].entry.input_buf[0].X ),
    .GATE(\l_fifo.genblk1[36].entry.empty ),
    .RESET_B(net10),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[35].entry.input_buf[0].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[36].entry.latch[1]  (.D(\l_fifo.genblk1[36].entry.input_buf[1].X ),
    .GATE(\l_fifo.genblk1[36].entry.empty ),
    .RESET_B(net8),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[35].entry.input_buf[1].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[36].entry.latch[2]  (.D(\l_fifo.genblk1[36].entry.input_buf[2].X ),
    .GATE(\l_fifo.genblk1[36].entry.empty ),
    .RESET_B(net11),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[35].entry.input_buf[2].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[36].entry.latch[3]  (.D(\l_fifo.genblk1[36].entry.input_buf[3].X ),
    .GATE(\l_fifo.genblk1[36].entry.empty ),
    .RESET_B(net18),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[35].entry.input_buf[3].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[36].entry.latch[4]  (.D(\l_fifo.genblk1[36].entry.input_buf[4].X ),
    .GATE(\l_fifo.genblk1[36].entry.empty ),
    .RESET_B(net12),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[35].entry.input_buf[4].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[36].entry.latch[5]  (.D(\l_fifo.genblk1[36].entry.input_buf[5].X ),
    .GATE(\l_fifo.genblk1[36].entry.empty ),
    .RESET_B(net10),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[35].entry.input_buf[5].A ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[37].entry.input_buf[0].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[37].entry.input_buf[0].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[37].entry.input_buf[0].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[37].entry.input_buf[0].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[37].entry.input_buf[0].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[37].entry.input_buf[0].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[37].entry.input_buf[1].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[37].entry.input_buf[1].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[37].entry.input_buf[1].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[37].entry.input_buf[1].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[37].entry.input_buf[1].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[37].entry.input_buf[1].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[37].entry.input_buf[2].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[37].entry.input_buf[2].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[37].entry.input_buf[2].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[37].entry.input_buf[2].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[37].entry.input_buf[2].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[37].entry.input_buf[2].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[37].entry.input_buf[3].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[37].entry.input_buf[3].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[37].entry.input_buf[3].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[37].entry.input_buf[3].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[37].entry.input_buf[3].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[37].entry.input_buf[3].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[37].entry.input_buf[4].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[37].entry.input_buf[4].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[37].entry.input_buf[4].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[37].entry.input_buf[4].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[37].entry.input_buf[4].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[37].entry.input_buf[4].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[37].entry.input_buf[5].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[37].entry.input_buf[5].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[37].entry.input_buf[5].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[37].entry.input_buf[5].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[37].entry.input_buf[5].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[37].entry.input_buf[5].X ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[37].entry.latch[0]  (.D(\l_fifo.genblk1[37].entry.input_buf[0].X ),
    .GATE(\l_fifo.genblk1[37].entry.empty ),
    .RESET_B(net11),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[36].entry.input_buf[0].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[37].entry.latch[1]  (.D(\l_fifo.genblk1[37].entry.input_buf[1].X ),
    .GATE(\l_fifo.genblk1[37].entry.empty ),
    .RESET_B(net10),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[36].entry.input_buf[1].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[37].entry.latch[2]  (.D(\l_fifo.genblk1[37].entry.input_buf[2].X ),
    .GATE(\l_fifo.genblk1[37].entry.empty ),
    .RESET_B(net11),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[36].entry.input_buf[2].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[37].entry.latch[3]  (.D(\l_fifo.genblk1[37].entry.input_buf[3].X ),
    .GATE(\l_fifo.genblk1[37].entry.empty ),
    .RESET_B(net8),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[36].entry.input_buf[3].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[37].entry.latch[4]  (.D(\l_fifo.genblk1[37].entry.input_buf[4].X ),
    .GATE(\l_fifo.genblk1[37].entry.empty ),
    .RESET_B(net10),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[36].entry.input_buf[4].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[37].entry.latch[5]  (.D(\l_fifo.genblk1[37].entry.input_buf[5].X ),
    .GATE(\l_fifo.genblk1[37].entry.empty ),
    .RESET_B(net11),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[36].entry.input_buf[5].A ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[38].entry.input_buf[0].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[38].entry.input_buf[0].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[38].entry.input_buf[0].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[38].entry.input_buf[0].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[38].entry.input_buf[0].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[38].entry.input_buf[0].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[38].entry.input_buf[1].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[38].entry.input_buf[1].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[38].entry.input_buf[1].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[38].entry.input_buf[1].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[38].entry.input_buf[1].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[38].entry.input_buf[1].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[38].entry.input_buf[2].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[38].entry.input_buf[2].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[38].entry.input_buf[2].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[38].entry.input_buf[2].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[38].entry.input_buf[2].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[38].entry.input_buf[2].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[38].entry.input_buf[3].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[38].entry.input_buf[3].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[38].entry.input_buf[3].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[38].entry.input_buf[3].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[38].entry.input_buf[3].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[38].entry.input_buf[3].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[38].entry.input_buf[4].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[38].entry.input_buf[4].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[38].entry.input_buf[4].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[38].entry.input_buf[4].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[38].entry.input_buf[4].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[38].entry.input_buf[4].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[38].entry.input_buf[5].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[38].entry.input_buf[5].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[38].entry.input_buf[5].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[38].entry.input_buf[5].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[38].entry.input_buf[5].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[38].entry.input_buf[5].X ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[38].entry.latch[0]  (.D(\l_fifo.genblk1[38].entry.input_buf[0].X ),
    .GATE(\l_fifo.genblk1[38].entry.empty ),
    .RESET_B(net18),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[37].entry.input_buf[0].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[38].entry.latch[1]  (.D(\l_fifo.genblk1[38].entry.input_buf[1].X ),
    .GATE(\l_fifo.genblk1[38].entry.empty ),
    .RESET_B(net18),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[37].entry.input_buf[1].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[38].entry.latch[2]  (.D(\l_fifo.genblk1[38].entry.input_buf[2].X ),
    .GATE(\l_fifo.genblk1[38].entry.empty ),
    .RESET_B(net18),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[37].entry.input_buf[2].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[38].entry.latch[3]  (.D(\l_fifo.genblk1[38].entry.input_buf[3].X ),
    .GATE(\l_fifo.genblk1[38].entry.empty ),
    .RESET_B(net11),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[37].entry.input_buf[3].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[38].entry.latch[4]  (.D(\l_fifo.genblk1[38].entry.input_buf[4].X ),
    .GATE(\l_fifo.genblk1[38].entry.empty ),
    .RESET_B(net21),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[37].entry.input_buf[4].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[38].entry.latch[5]  (.D(\l_fifo.genblk1[38].entry.input_buf[5].X ),
    .GATE(\l_fifo.genblk1[38].entry.empty ),
    .RESET_B(net11),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[37].entry.input_buf[5].A ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[39].entry.input_buf[0].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[39].entry.input_buf[0].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[39].entry.input_buf[0].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[39].entry.input_buf[0].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[39].entry.input_buf[0].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[39].entry.input_buf[0].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[39].entry.input_buf[1].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[39].entry.input_buf[1].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[39].entry.input_buf[1].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[39].entry.input_buf[1].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[39].entry.input_buf[1].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[39].entry.input_buf[1].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[39].entry.input_buf[2].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[39].entry.input_buf[2].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[39].entry.input_buf[2].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[39].entry.input_buf[2].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[39].entry.input_buf[2].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[39].entry.input_buf[2].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[39].entry.input_buf[3].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[39].entry.input_buf[3].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[39].entry.input_buf[3].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[39].entry.input_buf[3].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[39].entry.input_buf[3].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[39].entry.input_buf[3].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[39].entry.input_buf[4].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[39].entry.input_buf[4].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[39].entry.input_buf[4].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[39].entry.input_buf[4].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[39].entry.input_buf[4].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[39].entry.input_buf[4].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[39].entry.input_buf[5].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[39].entry.input_buf[5].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[39].entry.input_buf[5].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[39].entry.input_buf[5].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[39].entry.input_buf[5].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[39].entry.input_buf[5].X ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[39].entry.latch[0]  (.D(\l_fifo.genblk1[39].entry.input_buf[0].X ),
    .GATE(\l_fifo.genblk1[39].entry.empty ),
    .RESET_B(net18),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[38].entry.input_buf[0].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[39].entry.latch[1]  (.D(\l_fifo.genblk1[39].entry.input_buf[1].X ),
    .GATE(\l_fifo.genblk1[39].entry.empty ),
    .RESET_B(net18),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[38].entry.input_buf[1].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[39].entry.latch[2]  (.D(\l_fifo.genblk1[39].entry.input_buf[2].X ),
    .GATE(\l_fifo.genblk1[39].entry.empty ),
    .RESET_B(net21),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[38].entry.input_buf[2].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[39].entry.latch[3]  (.D(\l_fifo.genblk1[39].entry.input_buf[3].X ),
    .GATE(\l_fifo.genblk1[39].entry.empty ),
    .RESET_B(net18),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[38].entry.input_buf[3].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[39].entry.latch[4]  (.D(\l_fifo.genblk1[39].entry.input_buf[4].X ),
    .GATE(\l_fifo.genblk1[39].entry.empty ),
    .RESET_B(net20),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[38].entry.input_buf[4].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[39].entry.latch[5]  (.D(\l_fifo.genblk1[39].entry.input_buf[5].X ),
    .GATE(\l_fifo.genblk1[39].entry.empty ),
    .RESET_B(net18),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[38].entry.input_buf[5].A ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[3].entry.input_buf[0].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[3].entry.input_buf[0].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[3].entry.input_buf[0].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[3].entry.input_buf[0].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[3].entry.input_buf[0].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[3].entry.input_buf[0].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[3].entry.input_buf[1].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[3].entry.input_buf[1].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[3].entry.input_buf[1].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[3].entry.input_buf[1].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[3].entry.input_buf[1].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[3].entry.input_buf[1].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[3].entry.input_buf[2].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[3].entry.input_buf[2].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[3].entry.input_buf[2].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[3].entry.input_buf[2].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[3].entry.input_buf[2].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[3].entry.input_buf[2].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[3].entry.input_buf[3].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[3].entry.input_buf[3].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[3].entry.input_buf[3].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[3].entry.input_buf[3].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[3].entry.input_buf[3].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[3].entry.input_buf[3].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[3].entry.input_buf[4].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[3].entry.input_buf[4].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[3].entry.input_buf[4].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[3].entry.input_buf[4].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[3].entry.input_buf[4].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[3].entry.input_buf[4].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[3].entry.input_buf[5].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[3].entry.input_buf[5].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[3].entry.input_buf[5].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[3].entry.input_buf[5].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[3].entry.input_buf[5].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[3].entry.input_buf[5].X ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[3].entry.latch[0]  (.D(\l_fifo.genblk1[3].entry.input_buf[0].X ),
    .GATE(\l_fifo.genblk1[3].entry.empty ),
    .RESET_B(net32),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[2].entry.input_buf[0].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[3].entry.latch[1]  (.D(\l_fifo.genblk1[3].entry.input_buf[1].X ),
    .GATE(\l_fifo.genblk1[3].entry.empty ),
    .RESET_B(net32),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[2].entry.input_buf[1].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[3].entry.latch[2]  (.D(\l_fifo.genblk1[3].entry.input_buf[2].X ),
    .GATE(\l_fifo.genblk1[3].entry.empty ),
    .RESET_B(net28),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[2].entry.input_buf[2].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[3].entry.latch[3]  (.D(\l_fifo.genblk1[3].entry.input_buf[3].X ),
    .GATE(\l_fifo.genblk1[3].entry.empty ),
    .RESET_B(net32),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[2].entry.input_buf[3].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[3].entry.latch[4]  (.D(\l_fifo.genblk1[3].entry.input_buf[4].X ),
    .GATE(\l_fifo.genblk1[3].entry.empty ),
    .RESET_B(net29),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[2].entry.input_buf[4].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[3].entry.latch[5]  (.D(\l_fifo.genblk1[3].entry.input_buf[5].X ),
    .GATE(\l_fifo.genblk1[3].entry.empty ),
    .RESET_B(net32),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[2].entry.input_buf[5].A ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[40].entry.input_buf[0].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[40].entry.input_buf[0].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[40].entry.input_buf[0].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[40].entry.input_buf[0].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[40].entry.input_buf[0].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[40].entry.input_buf[0].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[40].entry.input_buf[1].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[40].entry.input_buf[1].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[40].entry.input_buf[1].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[40].entry.input_buf[1].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[40].entry.input_buf[1].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[40].entry.input_buf[1].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[40].entry.input_buf[2].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[40].entry.input_buf[2].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[40].entry.input_buf[2].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[40].entry.input_buf[2].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[40].entry.input_buf[2].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[40].entry.input_buf[2].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[40].entry.input_buf[3].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[40].entry.input_buf[3].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[40].entry.input_buf[3].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[40].entry.input_buf[3].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[40].entry.input_buf[3].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[40].entry.input_buf[3].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[40].entry.input_buf[4].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[40].entry.input_buf[4].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[40].entry.input_buf[4].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[40].entry.input_buf[4].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[40].entry.input_buf[4].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[40].entry.input_buf[4].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[40].entry.input_buf[5].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[40].entry.input_buf[5].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[40].entry.input_buf[5].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[40].entry.input_buf[5].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[40].entry.input_buf[5].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[40].entry.input_buf[5].X ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[40].entry.latch[0]  (.D(\l_fifo.genblk1[40].entry.input_buf[0].X ),
    .GATE(\l_fifo.genblk1[40].entry.empty ),
    .RESET_B(net19),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[39].entry.input_buf[0].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[40].entry.latch[1]  (.D(\l_fifo.genblk1[40].entry.input_buf[1].X ),
    .GATE(\l_fifo.genblk1[40].entry.empty ),
    .RESET_B(net19),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[39].entry.input_buf[1].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[40].entry.latch[2]  (.D(\l_fifo.genblk1[40].entry.input_buf[2].X ),
    .GATE(\l_fifo.genblk1[40].entry.empty ),
    .RESET_B(net20),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[39].entry.input_buf[2].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[40].entry.latch[3]  (.D(\l_fifo.genblk1[40].entry.input_buf[3].X ),
    .GATE(\l_fifo.genblk1[40].entry.empty ),
    .RESET_B(net18),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[39].entry.input_buf[3].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[40].entry.latch[4]  (.D(\l_fifo.genblk1[40].entry.input_buf[4].X ),
    .GATE(\l_fifo.genblk1[40].entry.empty ),
    .RESET_B(net20),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[39].entry.input_buf[4].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[40].entry.latch[5]  (.D(\l_fifo.genblk1[40].entry.input_buf[5].X ),
    .GATE(\l_fifo.genblk1[40].entry.empty ),
    .RESET_B(net20),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[39].entry.input_buf[5].A ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[41].entry.input_buf[0].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[41].entry.input_buf[0].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[41].entry.input_buf[0].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[41].entry.input_buf[0].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[41].entry.input_buf[0].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[41].entry.input_buf[0].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[41].entry.input_buf[1].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[41].entry.input_buf[1].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[41].entry.input_buf[1].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[41].entry.input_buf[1].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[41].entry.input_buf[1].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[41].entry.input_buf[1].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[41].entry.input_buf[2].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[41].entry.input_buf[2].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[41].entry.input_buf[2].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[41].entry.input_buf[2].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[41].entry.input_buf[2].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[41].entry.input_buf[2].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[41].entry.input_buf[3].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[41].entry.input_buf[3].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[41].entry.input_buf[3].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[41].entry.input_buf[3].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[41].entry.input_buf[3].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[41].entry.input_buf[3].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[41].entry.input_buf[4].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[41].entry.input_buf[4].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[41].entry.input_buf[4].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[41].entry.input_buf[4].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[41].entry.input_buf[4].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[41].entry.input_buf[4].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[41].entry.input_buf[5].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[41].entry.input_buf[5].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[41].entry.input_buf[5].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[41].entry.input_buf[5].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[41].entry.input_buf[5].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[41].entry.input_buf[5].X ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[41].entry.latch[0]  (.D(\l_fifo.genblk1[41].entry.input_buf[0].X ),
    .GATE(\l_fifo.genblk1[41].entry.empty ),
    .RESET_B(net19),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[40].entry.input_buf[0].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[41].entry.latch[1]  (.D(\l_fifo.genblk1[41].entry.input_buf[1].X ),
    .GATE(\l_fifo.genblk1[41].entry.empty ),
    .RESET_B(net19),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[40].entry.input_buf[1].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[41].entry.latch[2]  (.D(\l_fifo.genblk1[41].entry.input_buf[2].X ),
    .GATE(\l_fifo.genblk1[41].entry.empty ),
    .RESET_B(net38),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[40].entry.input_buf[2].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[41].entry.latch[3]  (.D(\l_fifo.genblk1[41].entry.input_buf[3].X ),
    .GATE(\l_fifo.genblk1[41].entry.empty ),
    .RESET_B(net19),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[40].entry.input_buf[3].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[41].entry.latch[4]  (.D(\l_fifo.genblk1[41].entry.input_buf[4].X ),
    .GATE(\l_fifo.genblk1[41].entry.empty ),
    .RESET_B(net35),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[40].entry.input_buf[4].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[41].entry.latch[5]  (.D(\l_fifo.genblk1[41].entry.input_buf[5].X ),
    .GATE(\l_fifo.genblk1[41].entry.empty ),
    .RESET_B(net19),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[40].entry.input_buf[5].A ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[42].entry.input_buf[0].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[42].entry.input_buf[0].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[42].entry.input_buf[0].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[42].entry.input_buf[0].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[42].entry.input_buf[0].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[42].entry.input_buf[0].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[42].entry.input_buf[1].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[42].entry.input_buf[1].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[42].entry.input_buf[1].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[42].entry.input_buf[1].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[42].entry.input_buf[1].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[42].entry.input_buf[1].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[42].entry.input_buf[2].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[42].entry.input_buf[2].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[42].entry.input_buf[2].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[42].entry.input_buf[2].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[42].entry.input_buf[2].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[42].entry.input_buf[2].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[42].entry.input_buf[3].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[42].entry.input_buf[3].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[42].entry.input_buf[3].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[42].entry.input_buf[3].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[42].entry.input_buf[3].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[42].entry.input_buf[3].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[42].entry.input_buf[4].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[42].entry.input_buf[4].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[42].entry.input_buf[4].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[42].entry.input_buf[4].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[42].entry.input_buf[4].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[42].entry.input_buf[4].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[42].entry.input_buf[5].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[42].entry.input_buf[5].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[42].entry.input_buf[5].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[42].entry.input_buf[5].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[42].entry.input_buf[5].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[42].entry.input_buf[5].X ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[42].entry.latch[0]  (.D(\l_fifo.genblk1[42].entry.input_buf[0].X ),
    .GATE(\l_fifo.genblk1[42].entry.empty ),
    .RESET_B(net26),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[41].entry.input_buf[0].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[42].entry.latch[1]  (.D(\l_fifo.genblk1[42].entry.input_buf[1].X ),
    .GATE(\l_fifo.genblk1[42].entry.empty ),
    .RESET_B(net9),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[41].entry.input_buf[1].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[42].entry.latch[2]  (.D(\l_fifo.genblk1[42].entry.input_buf[2].X ),
    .GATE(\l_fifo.genblk1[42].entry.empty ),
    .RESET_B(net35),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[41].entry.input_buf[2].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[42].entry.latch[3]  (.D(\l_fifo.genblk1[42].entry.input_buf[3].X ),
    .GATE(\l_fifo.genblk1[42].entry.empty ),
    .RESET_B(net27),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[41].entry.input_buf[3].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[42].entry.latch[4]  (.D(\l_fifo.genblk1[42].entry.input_buf[4].X ),
    .GATE(\l_fifo.genblk1[42].entry.empty ),
    .RESET_B(net35),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[41].entry.input_buf[4].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[42].entry.latch[5]  (.D(\l_fifo.genblk1[42].entry.input_buf[5].X ),
    .GATE(\l_fifo.genblk1[42].entry.empty ),
    .RESET_B(net19),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[41].entry.input_buf[5].A ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[43].entry.input_buf[0].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[43].entry.input_buf[0].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[43].entry.input_buf[0].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[43].entry.input_buf[0].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[43].entry.input_buf[0].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[43].entry.input_buf[0].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[43].entry.input_buf[1].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[43].entry.input_buf[1].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[43].entry.input_buf[1].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[43].entry.input_buf[1].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[43].entry.input_buf[1].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[43].entry.input_buf[1].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[43].entry.input_buf[2].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[43].entry.input_buf[2].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[43].entry.input_buf[2].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[43].entry.input_buf[2].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[43].entry.input_buf[2].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[43].entry.input_buf[2].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[43].entry.input_buf[3].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[43].entry.input_buf[3].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[43].entry.input_buf[3].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[43].entry.input_buf[3].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[43].entry.input_buf[3].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[43].entry.input_buf[3].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[43].entry.input_buf[4].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[43].entry.input_buf[4].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[43].entry.input_buf[4].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[43].entry.input_buf[4].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[43].entry.input_buf[4].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[43].entry.input_buf[4].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[43].entry.input_buf[5].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[43].entry.input_buf[5].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[43].entry.input_buf[5].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[43].entry.input_buf[5].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[43].entry.input_buf[5].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[43].entry.input_buf[5].X ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[43].entry.latch[0]  (.D(\l_fifo.genblk1[43].entry.input_buf[0].X ),
    .GATE(\l_fifo.genblk1[43].entry.empty ),
    .RESET_B(net9),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[42].entry.input_buf[0].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[43].entry.latch[1]  (.D(\l_fifo.genblk1[43].entry.input_buf[1].X ),
    .GATE(\l_fifo.genblk1[43].entry.empty ),
    .RESET_B(net27),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[42].entry.input_buf[1].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[43].entry.latch[2]  (.D(\l_fifo.genblk1[43].entry.input_buf[2].X ),
    .GATE(\l_fifo.genblk1[43].entry.empty ),
    .RESET_B(net35),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[42].entry.input_buf[2].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[43].entry.latch[3]  (.D(\l_fifo.genblk1[43].entry.input_buf[3].X ),
    .GATE(\l_fifo.genblk1[43].entry.empty ),
    .RESET_B(net26),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[42].entry.input_buf[3].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[43].entry.latch[4]  (.D(\l_fifo.genblk1[43].entry.input_buf[4].X ),
    .GATE(\l_fifo.genblk1[43].entry.empty ),
    .RESET_B(net35),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[42].entry.input_buf[4].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[43].entry.latch[5]  (.D(\l_fifo.genblk1[43].entry.input_buf[5].X ),
    .GATE(\l_fifo.genblk1[43].entry.empty ),
    .RESET_B(net19),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[42].entry.input_buf[5].A ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[44].entry.input_buf[0].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[44].entry.input_buf[0].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[44].entry.input_buf[0].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[44].entry.input_buf[0].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[44].entry.input_buf[0].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[44].entry.input_buf[0].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[44].entry.input_buf[1].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[44].entry.input_buf[1].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[44].entry.input_buf[1].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[44].entry.input_buf[1].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[44].entry.input_buf[1].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[44].entry.input_buf[1].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[44].entry.input_buf[2].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[44].entry.input_buf[2].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[44].entry.input_buf[2].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[44].entry.input_buf[2].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[44].entry.input_buf[2].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[44].entry.input_buf[2].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[44].entry.input_buf[3].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[44].entry.input_buf[3].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[44].entry.input_buf[3].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[44].entry.input_buf[3].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[44].entry.input_buf[3].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[44].entry.input_buf[3].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[44].entry.input_buf[4].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[44].entry.input_buf[4].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[44].entry.input_buf[4].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[44].entry.input_buf[4].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[44].entry.input_buf[4].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[44].entry.input_buf[4].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[44].entry.input_buf[5].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[44].entry.input_buf[5].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[44].entry.input_buf[5].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[44].entry.input_buf[5].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[44].entry.input_buf[5].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[44].entry.input_buf[5].X ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[44].entry.latch[0]  (.D(\l_fifo.genblk1[44].entry.input_buf[0].X ),
    .GATE(\l_fifo.genblk1[44].entry.empty ),
    .RESET_B(net8),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[43].entry.input_buf[0].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[44].entry.latch[1]  (.D(\l_fifo.genblk1[44].entry.input_buf[1].X ),
    .GATE(\l_fifo.genblk1[44].entry.empty ),
    .RESET_B(net27),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[43].entry.input_buf[1].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[44].entry.latch[2]  (.D(\l_fifo.genblk1[44].entry.input_buf[2].X ),
    .GATE(\l_fifo.genblk1[44].entry.empty ),
    .RESET_B(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[43].entry.input_buf[2].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[44].entry.latch[3]  (.D(\l_fifo.genblk1[44].entry.input_buf[3].X ),
    .GATE(\l_fifo.genblk1[44].entry.empty ),
    .RESET_B(net26),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[43].entry.input_buf[3].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[44].entry.latch[4]  (.D(\l_fifo.genblk1[44].entry.input_buf[4].X ),
    .GATE(\l_fifo.genblk1[44].entry.empty ),
    .RESET_B(net27),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[43].entry.input_buf[4].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[44].entry.latch[5]  (.D(\l_fifo.genblk1[44].entry.input_buf[5].X ),
    .GATE(\l_fifo.genblk1[44].entry.empty ),
    .RESET_B(net26),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[43].entry.input_buf[5].A ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[45].entry.input_buf[0].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[45].entry.input_buf[0].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[45].entry.input_buf[0].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[45].entry.input_buf[0].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[45].entry.input_buf[0].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[45].entry.input_buf[0].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[45].entry.input_buf[1].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[45].entry.input_buf[1].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[45].entry.input_buf[1].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[45].entry.input_buf[1].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[45].entry.input_buf[1].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[45].entry.input_buf[1].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[45].entry.input_buf[2].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[45].entry.input_buf[2].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[45].entry.input_buf[2].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[45].entry.input_buf[2].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[45].entry.input_buf[2].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[45].entry.input_buf[2].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[45].entry.input_buf[3].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[45].entry.input_buf[3].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[45].entry.input_buf[3].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[45].entry.input_buf[3].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[45].entry.input_buf[3].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[45].entry.input_buf[3].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[45].entry.input_buf[4].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[45].entry.input_buf[4].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[45].entry.input_buf[4].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[45].entry.input_buf[4].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[45].entry.input_buf[4].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[45].entry.input_buf[4].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[45].entry.input_buf[5].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[45].entry.input_buf[5].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[45].entry.input_buf[5].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[45].entry.input_buf[5].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[45].entry.input_buf[5].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[45].entry.input_buf[5].X ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[45].entry.latch[0]  (.D(\l_fifo.genblk1[45].entry.input_buf[0].X ),
    .GATE(\l_fifo.genblk1[45].entry.empty ),
    .RESET_B(net8),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[44].entry.input_buf[0].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[45].entry.latch[1]  (.D(\l_fifo.genblk1[45].entry.input_buf[1].X ),
    .GATE(\l_fifo.genblk1[45].entry.empty ),
    .RESET_B(net26),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[44].entry.input_buf[1].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[45].entry.latch[2]  (.D(\l_fifo.genblk1[45].entry.input_buf[2].X ),
    .GATE(\l_fifo.genblk1[45].entry.empty ),
    .RESET_B(net27),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[44].entry.input_buf[2].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[45].entry.latch[3]  (.D(\l_fifo.genblk1[45].entry.input_buf[3].X ),
    .GATE(\l_fifo.genblk1[45].entry.empty ),
    .RESET_B(net26),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[44].entry.input_buf[3].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[45].entry.latch[4]  (.D(\l_fifo.genblk1[45].entry.input_buf[4].X ),
    .GATE(\l_fifo.genblk1[45].entry.empty ),
    .RESET_B(net31),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[44].entry.input_buf[4].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[45].entry.latch[5]  (.D(\l_fifo.genblk1[45].entry.input_buf[5].X ),
    .GATE(\l_fifo.genblk1[45].entry.empty ),
    .RESET_B(net31),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[44].entry.input_buf[5].A ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[46].entry.input_buf[0].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[46].entry.input_buf[0].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[46].entry.input_buf[0].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[46].entry.input_buf[0].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[46].entry.input_buf[0].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[46].entry.input_buf[0].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[46].entry.input_buf[1].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[46].entry.input_buf[1].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[46].entry.input_buf[1].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[46].entry.input_buf[1].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[46].entry.input_buf[1].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[46].entry.input_buf[1].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[46].entry.input_buf[2].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[46].entry.input_buf[2].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[46].entry.input_buf[2].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[46].entry.input_buf[2].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[46].entry.input_buf[2].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[46].entry.input_buf[2].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[46].entry.input_buf[3].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[46].entry.input_buf[3].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[46].entry.input_buf[3].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[46].entry.input_buf[3].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[46].entry.input_buf[3].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[46].entry.input_buf[3].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[46].entry.input_buf[4].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[46].entry.input_buf[4].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[46].entry.input_buf[4].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[46].entry.input_buf[4].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[46].entry.input_buf[4].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[46].entry.input_buf[4].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[46].entry.input_buf[5].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[46].entry.input_buf[5].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[46].entry.input_buf[5].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[46].entry.input_buf[5].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[46].entry.input_buf[5].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[46].entry.input_buf[5].X ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[46].entry.latch[0]  (.D(\l_fifo.genblk1[46].entry.input_buf[0].X ),
    .GATE(\l_fifo.genblk1[46].entry.empty ),
    .RESET_B(net26),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[45].entry.input_buf[0].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[46].entry.latch[1]  (.D(\l_fifo.genblk1[46].entry.input_buf[1].X ),
    .GATE(\l_fifo.genblk1[46].entry.empty ),
    .RESET_B(net31),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[45].entry.input_buf[1].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[46].entry.latch[2]  (.D(\l_fifo.genblk1[46].entry.input_buf[2].X ),
    .GATE(\l_fifo.genblk1[46].entry.empty ),
    .RESET_B(net31),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[45].entry.input_buf[2].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[46].entry.latch[3]  (.D(\l_fifo.genblk1[46].entry.input_buf[3].X ),
    .GATE(\l_fifo.genblk1[46].entry.empty ),
    .RESET_B(net30),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[45].entry.input_buf[3].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[46].entry.latch[4]  (.D(\l_fifo.genblk1[46].entry.input_buf[4].X ),
    .GATE(\l_fifo.genblk1[46].entry.empty ),
    .RESET_B(net32),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[45].entry.input_buf[4].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[46].entry.latch[5]  (.D(\l_fifo.genblk1[46].entry.input_buf[5].X ),
    .GATE(\l_fifo.genblk1[46].entry.empty ),
    .RESET_B(net30),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[45].entry.input_buf[5].A ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[47].entry.input_buf[0].genblk1[0].genblk1.buf_first  (.A(\data_in_buffer[0].X ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[47].entry.input_buf[0].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[47].entry.input_buf[0].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[47].entry.input_buf[0].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[47].entry.input_buf[0].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[47].entry.input_buf[1].genblk1[0].genblk1.buf_first  (.A(\data_in_buffer[1].X ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[47].entry.input_buf[1].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[47].entry.input_buf[1].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[47].entry.input_buf[1].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[47].entry.input_buf[1].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[47].entry.input_buf[2].genblk1[0].genblk1.buf_first  (.A(\data_in_buffer[2].X ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[47].entry.input_buf[2].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[47].entry.input_buf[2].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[47].entry.input_buf[2].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[47].entry.input_buf[2].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[47].entry.input_buf[3].genblk1[0].genblk1.buf_first  (.A(\data_in_buffer[3].X ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[47].entry.input_buf[3].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[47].entry.input_buf[3].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[47].entry.input_buf[3].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[47].entry.input_buf[3].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[47].entry.input_buf[4].genblk1[0].genblk1.buf_first  (.A(\data_in_buffer[4].X ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[47].entry.input_buf[4].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[47].entry.input_buf[4].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[47].entry.input_buf[4].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[47].entry.input_buf[4].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[47].entry.input_buf[5].genblk1[0].genblk1.buf_first  (.A(\data_in_buffer[5].X ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[47].entry.input_buf[5].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[47].entry.input_buf[5].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[47].entry.input_buf[5].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[47].entry.input_buf[5].X ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[47].entry.latch[0]  (.D(\l_fifo.genblk1[47].entry.input_buf[0].X ),
    .GATE(\l_fifo.genblk1[47].entry.empty ),
    .RESET_B(net26),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[46].entry.input_buf[0].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[47].entry.latch[1]  (.D(\l_fifo.genblk1[47].entry.input_buf[1].X ),
    .GATE(\l_fifo.genblk1[47].entry.empty ),
    .RESET_B(net30),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[46].entry.input_buf[1].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[47].entry.latch[2]  (.D(\l_fifo.genblk1[47].entry.input_buf[2].X ),
    .GATE(\l_fifo.genblk1[47].entry.empty ),
    .RESET_B(net49),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[46].entry.input_buf[2].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[47].entry.latch[3]  (.D(\l_fifo.genblk1[47].entry.input_buf[3].X ),
    .GATE(\l_fifo.genblk1[47].entry.empty ),
    .RESET_B(net28),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[46].entry.input_buf[3].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[47].entry.latch[4]  (.D(\l_fifo.genblk1[47].entry.input_buf[4].X ),
    .GATE(\l_fifo.genblk1[47].entry.empty ),
    .RESET_B(net28),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[46].entry.input_buf[4].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[47].entry.latch[5]  (.D(\l_fifo.genblk1[47].entry.input_buf[5].X ),
    .GATE(\l_fifo.genblk1[47].entry.empty ),
    .RESET_B(net28),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[46].entry.input_buf[5].A ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[4].entry.input_buf[0].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[4].entry.input_buf[0].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[4].entry.input_buf[0].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[4].entry.input_buf[0].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[4].entry.input_buf[0].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[4].entry.input_buf[0].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[4].entry.input_buf[1].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[4].entry.input_buf[1].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[4].entry.input_buf[1].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[4].entry.input_buf[1].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[4].entry.input_buf[1].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[4].entry.input_buf[1].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[4].entry.input_buf[2].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[4].entry.input_buf[2].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[4].entry.input_buf[2].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[4].entry.input_buf[2].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[4].entry.input_buf[2].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[4].entry.input_buf[2].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[4].entry.input_buf[3].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[4].entry.input_buf[3].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[4].entry.input_buf[3].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[4].entry.input_buf[3].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[4].entry.input_buf[3].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[4].entry.input_buf[3].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[4].entry.input_buf[4].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[4].entry.input_buf[4].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[4].entry.input_buf[4].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[4].entry.input_buf[4].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[4].entry.input_buf[4].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[4].entry.input_buf[4].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[4].entry.input_buf[5].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[4].entry.input_buf[5].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[4].entry.input_buf[5].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[4].entry.input_buf[5].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[4].entry.input_buf[5].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[4].entry.input_buf[5].X ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[4].entry.latch[0]  (.D(\l_fifo.genblk1[4].entry.input_buf[0].X ),
    .GATE(\l_fifo.genblk1[4].entry.empty ),
    .RESET_B(net32),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[3].entry.input_buf[0].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[4].entry.latch[1]  (.D(\l_fifo.genblk1[4].entry.input_buf[1].X ),
    .GATE(\l_fifo.genblk1[4].entry.empty ),
    .RESET_B(net30),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[3].entry.input_buf[1].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[4].entry.latch[2]  (.D(\l_fifo.genblk1[4].entry.input_buf[2].X ),
    .GATE(\l_fifo.genblk1[4].entry.empty ),
    .RESET_B(net32),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[3].entry.input_buf[2].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[4].entry.latch[3]  (.D(\l_fifo.genblk1[4].entry.input_buf[3].X ),
    .GATE(\l_fifo.genblk1[4].entry.empty ),
    .RESET_B(net33),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[3].entry.input_buf[3].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[4].entry.latch[4]  (.D(\l_fifo.genblk1[4].entry.input_buf[4].X ),
    .GATE(\l_fifo.genblk1[4].entry.empty ),
    .RESET_B(net30),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[3].entry.input_buf[4].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[4].entry.latch[5]  (.D(\l_fifo.genblk1[4].entry.input_buf[5].X ),
    .GATE(\l_fifo.genblk1[4].entry.empty ),
    .RESET_B(net32),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[3].entry.input_buf[5].A ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[5].entry.input_buf[0].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[5].entry.input_buf[0].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[5].entry.input_buf[0].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[5].entry.input_buf[0].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[5].entry.input_buf[0].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[5].entry.input_buf[0].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[5].entry.input_buf[1].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[5].entry.input_buf[1].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[5].entry.input_buf[1].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[5].entry.input_buf[1].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[5].entry.input_buf[1].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[5].entry.input_buf[1].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[5].entry.input_buf[2].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[5].entry.input_buf[2].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[5].entry.input_buf[2].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[5].entry.input_buf[2].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[5].entry.input_buf[2].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[5].entry.input_buf[2].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[5].entry.input_buf[3].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[5].entry.input_buf[3].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[5].entry.input_buf[3].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[5].entry.input_buf[3].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[5].entry.input_buf[3].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[5].entry.input_buf[3].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[5].entry.input_buf[4].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[5].entry.input_buf[4].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[5].entry.input_buf[4].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[5].entry.input_buf[4].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[5].entry.input_buf[4].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[5].entry.input_buf[4].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[5].entry.input_buf[5].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[5].entry.input_buf[5].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[5].entry.input_buf[5].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[5].entry.input_buf[5].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[5].entry.input_buf[5].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[5].entry.input_buf[5].X ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[5].entry.latch[0]  (.D(\l_fifo.genblk1[5].entry.input_buf[0].X ),
    .GATE(\l_fifo.genblk1[5].entry.empty ),
    .RESET_B(net30),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[4].entry.input_buf[0].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[5].entry.latch[1]  (.D(\l_fifo.genblk1[5].entry.input_buf[1].X ),
    .GATE(\l_fifo.genblk1[5].entry.empty ),
    .RESET_B(net32),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[4].entry.input_buf[1].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[5].entry.latch[2]  (.D(\l_fifo.genblk1[5].entry.input_buf[2].X ),
    .GATE(\l_fifo.genblk1[5].entry.empty ),
    .RESET_B(net30),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[4].entry.input_buf[2].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[5].entry.latch[3]  (.D(\l_fifo.genblk1[5].entry.input_buf[3].X ),
    .GATE(\l_fifo.genblk1[5].entry.empty ),
    .RESET_B(net32),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[4].entry.input_buf[3].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[5].entry.latch[4]  (.D(\l_fifo.genblk1[5].entry.input_buf[4].X ),
    .GATE(\l_fifo.genblk1[5].entry.empty ),
    .RESET_B(net43),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[4].entry.input_buf[4].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[5].entry.latch[5]  (.D(\l_fifo.genblk1[5].entry.input_buf[5].X ),
    .GATE(\l_fifo.genblk1[5].entry.empty ),
    .RESET_B(net33),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[4].entry.input_buf[5].A ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[6].entry.input_buf[0].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[6].entry.input_buf[0].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[6].entry.input_buf[0].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[6].entry.input_buf[0].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[6].entry.input_buf[0].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[6].entry.input_buf[0].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[6].entry.input_buf[1].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[6].entry.input_buf[1].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[6].entry.input_buf[1].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[6].entry.input_buf[1].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[6].entry.input_buf[1].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[6].entry.input_buf[1].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[6].entry.input_buf[2].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[6].entry.input_buf[2].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[6].entry.input_buf[2].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[6].entry.input_buf[2].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[6].entry.input_buf[2].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[6].entry.input_buf[2].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[6].entry.input_buf[3].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[6].entry.input_buf[3].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[6].entry.input_buf[3].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[6].entry.input_buf[3].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[6].entry.input_buf[3].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[6].entry.input_buf[3].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[6].entry.input_buf[4].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[6].entry.input_buf[4].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[6].entry.input_buf[4].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[6].entry.input_buf[4].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[6].entry.input_buf[4].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[6].entry.input_buf[4].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[6].entry.input_buf[5].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[6].entry.input_buf[5].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[6].entry.input_buf[5].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[6].entry.input_buf[5].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[6].entry.input_buf[5].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[6].entry.input_buf[5].X ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[6].entry.latch[0]  (.D(\l_fifo.genblk1[6].entry.input_buf[0].X ),
    .GATE(\l_fifo.genblk1[6].entry.empty ),
    .RESET_B(net27),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[5].entry.input_buf[0].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[6].entry.latch[1]  (.D(\l_fifo.genblk1[6].entry.input_buf[1].X ),
    .GATE(\l_fifo.genblk1[6].entry.empty ),
    .RESET_B(net31),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[5].entry.input_buf[1].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[6].entry.latch[2]  (.D(\l_fifo.genblk1[6].entry.input_buf[2].X ),
    .GATE(\l_fifo.genblk1[6].entry.empty ),
    .RESET_B(net31),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[5].entry.input_buf[2].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[6].entry.latch[3]  (.D(\l_fifo.genblk1[6].entry.input_buf[3].X ),
    .GATE(\l_fifo.genblk1[6].entry.empty ),
    .RESET_B(net31),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[5].entry.input_buf[3].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[6].entry.latch[4]  (.D(\l_fifo.genblk1[6].entry.input_buf[4].X ),
    .GATE(\l_fifo.genblk1[6].entry.empty ),
    .RESET_B(net30),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[5].entry.input_buf[4].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[6].entry.latch[5]  (.D(\l_fifo.genblk1[6].entry.input_buf[5].X ),
    .GATE(\l_fifo.genblk1[6].entry.empty ),
    .RESET_B(net43),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[5].entry.input_buf[5].A ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[7].entry.input_buf[0].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[7].entry.input_buf[0].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[7].entry.input_buf[0].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[7].entry.input_buf[0].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[7].entry.input_buf[0].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[7].entry.input_buf[0].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[7].entry.input_buf[1].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[7].entry.input_buf[1].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[7].entry.input_buf[1].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[7].entry.input_buf[1].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[7].entry.input_buf[1].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[7].entry.input_buf[1].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[7].entry.input_buf[2].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[7].entry.input_buf[2].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[7].entry.input_buf[2].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[7].entry.input_buf[2].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[7].entry.input_buf[2].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[7].entry.input_buf[2].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[7].entry.input_buf[3].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[7].entry.input_buf[3].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[7].entry.input_buf[3].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[7].entry.input_buf[3].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[7].entry.input_buf[3].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[7].entry.input_buf[3].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[7].entry.input_buf[4].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[7].entry.input_buf[4].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[7].entry.input_buf[4].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[7].entry.input_buf[4].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[7].entry.input_buf[4].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[7].entry.input_buf[4].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[7].entry.input_buf[5].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[7].entry.input_buf[5].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[7].entry.input_buf[5].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[7].entry.input_buf[5].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[7].entry.input_buf[5].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[7].entry.input_buf[5].X ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[7].entry.latch[0]  (.D(\l_fifo.genblk1[7].entry.input_buf[0].X ),
    .GATE(\l_fifo.genblk1[7].entry.empty ),
    .RESET_B(net38),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[6].entry.input_buf[0].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[7].entry.latch[1]  (.D(\l_fifo.genblk1[7].entry.input_buf[1].X ),
    .GATE(\l_fifo.genblk1[7].entry.empty ),
    .RESET_B(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[6].entry.input_buf[1].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[7].entry.latch[2]  (.D(\l_fifo.genblk1[7].entry.input_buf[2].X ),
    .GATE(\l_fifo.genblk1[7].entry.empty ),
    .RESET_B(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[6].entry.input_buf[2].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[7].entry.latch[3]  (.D(\l_fifo.genblk1[7].entry.input_buf[3].X ),
    .GATE(\l_fifo.genblk1[7].entry.empty ),
    .RESET_B(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[6].entry.input_buf[3].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[7].entry.latch[4]  (.D(\l_fifo.genblk1[7].entry.input_buf[4].X ),
    .GATE(\l_fifo.genblk1[7].entry.empty ),
    .RESET_B(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[6].entry.input_buf[4].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[7].entry.latch[5]  (.D(\l_fifo.genblk1[7].entry.input_buf[5].X ),
    .GATE(\l_fifo.genblk1[7].entry.empty ),
    .RESET_B(net37),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[6].entry.input_buf[5].A ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[8].entry.input_buf[0].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[8].entry.input_buf[0].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[8].entry.input_buf[0].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[8].entry.input_buf[0].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[8].entry.input_buf[0].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[8].entry.input_buf[0].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[8].entry.input_buf[1].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[8].entry.input_buf[1].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[8].entry.input_buf[1].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[8].entry.input_buf[1].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[8].entry.input_buf[1].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[8].entry.input_buf[1].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[8].entry.input_buf[2].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[8].entry.input_buf[2].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[8].entry.input_buf[2].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[8].entry.input_buf[2].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[8].entry.input_buf[2].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[8].entry.input_buf[2].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[8].entry.input_buf[3].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[8].entry.input_buf[3].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[8].entry.input_buf[3].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[8].entry.input_buf[3].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[8].entry.input_buf[3].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[8].entry.input_buf[3].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[8].entry.input_buf[4].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[8].entry.input_buf[4].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[8].entry.input_buf[4].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[8].entry.input_buf[4].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[8].entry.input_buf[4].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[8].entry.input_buf[4].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[8].entry.input_buf[5].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[8].entry.input_buf[5].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[8].entry.input_buf[5].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[8].entry.input_buf[5].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[8].entry.input_buf[5].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[8].entry.input_buf[5].X ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[8].entry.latch[0]  (.D(\l_fifo.genblk1[8].entry.input_buf[0].X ),
    .GATE(\l_fifo.genblk1[8].entry.empty ),
    .RESET_B(net35),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[7].entry.input_buf[0].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[8].entry.latch[1]  (.D(\l_fifo.genblk1[8].entry.input_buf[1].X ),
    .GATE(\l_fifo.genblk1[8].entry.empty ),
    .RESET_B(net35),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[7].entry.input_buf[1].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[8].entry.latch[2]  (.D(\l_fifo.genblk1[8].entry.input_buf[2].X ),
    .GATE(\l_fifo.genblk1[8].entry.empty ),
    .RESET_B(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[7].entry.input_buf[2].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[8].entry.latch[3]  (.D(\l_fifo.genblk1[8].entry.input_buf[3].X ),
    .GATE(\l_fifo.genblk1[8].entry.empty ),
    .RESET_B(net35),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[7].entry.input_buf[3].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[8].entry.latch[4]  (.D(\l_fifo.genblk1[8].entry.input_buf[4].X ),
    .GATE(\l_fifo.genblk1[8].entry.empty ),
    .RESET_B(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[7].entry.input_buf[4].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[8].entry.latch[5]  (.D(\l_fifo.genblk1[8].entry.input_buf[5].X ),
    .GATE(\l_fifo.genblk1[8].entry.empty ),
    .RESET_B(net38),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[7].entry.input_buf[5].A ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[9].entry.input_buf[0].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[9].entry.input_buf[0].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[9].entry.input_buf[0].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[9].entry.input_buf[0].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[9].entry.input_buf[0].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[9].entry.input_buf[0].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[9].entry.input_buf[1].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[9].entry.input_buf[1].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[9].entry.input_buf[1].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[9].entry.input_buf[1].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[9].entry.input_buf[1].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[9].entry.input_buf[1].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[9].entry.input_buf[2].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[9].entry.input_buf[2].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[9].entry.input_buf[2].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[9].entry.input_buf[2].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[9].entry.input_buf[2].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[9].entry.input_buf[2].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[9].entry.input_buf[3].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[9].entry.input_buf[3].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[9].entry.input_buf[3].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[9].entry.input_buf[3].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[9].entry.input_buf[3].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[9].entry.input_buf[3].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[9].entry.input_buf[4].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[9].entry.input_buf[4].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[9].entry.input_buf[4].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[9].entry.input_buf[4].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[9].entry.input_buf[4].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[9].entry.input_buf[4].X ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[9].entry.input_buf[5].genblk1[0].genblk1.buf_first  (.A(\l_fifo.genblk1[9].entry.input_buf[5].A ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[9].entry.input_buf[5].genblk1[0].mid ));
 sky130_fd_sc_hd__clkbuf_1 \l_fifo.genblk1[9].entry.input_buf[5].genblk1[0].genblk2.buf_last  (.A(\l_fifo.genblk1[9].entry.input_buf[5].genblk1[0].mid ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\l_fifo.genblk1[9].entry.input_buf[5].X ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[9].entry.latch[0]  (.D(\l_fifo.genblk1[9].entry.input_buf[0].X ),
    .GATE(\l_fifo.genblk1[10].entry.next_is_empty ),
    .RESET_B(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[8].entry.input_buf[0].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[9].entry.latch[1]  (.D(\l_fifo.genblk1[9].entry.input_buf[1].X ),
    .GATE(\l_fifo.genblk1[10].entry.next_is_empty ),
    .RESET_B(net37),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[8].entry.input_buf[1].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[9].entry.latch[2]  (.D(\l_fifo.genblk1[9].entry.input_buf[2].X ),
    .GATE(\l_fifo.genblk1[10].entry.next_is_empty ),
    .RESET_B(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[8].entry.input_buf[2].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[9].entry.latch[3]  (.D(\l_fifo.genblk1[9].entry.input_buf[3].X ),
    .GATE(\l_fifo.genblk1[10].entry.next_is_empty ),
    .RESET_B(net37),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[8].entry.input_buf[3].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[9].entry.latch[4]  (.D(\l_fifo.genblk1[9].entry.input_buf[4].X ),
    .GATE(\l_fifo.genblk1[10].entry.next_is_empty ),
    .RESET_B(net44),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[8].entry.input_buf[4].A ));
 sky130_fd_sc_hd__dlrtp_1 \l_fifo.genblk1[9].entry.latch[5]  (.D(\l_fifo.genblk1[9].entry.input_buf[5].X ),
    .GATE(\l_fifo.genblk1[10].entry.next_is_empty ),
    .RESET_B(net37),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\l_fifo.genblk1[8].entry.input_buf[5].A ));
endmodule
