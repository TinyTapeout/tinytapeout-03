// This is the unpowered netlist.
module scan_controller (clk,
    la_scan_clk_in,
    la_scan_data_in,
    la_scan_data_out,
    la_scan_latch_en,
    la_scan_select,
    ready,
    reset,
    scan_clk_in,
    scan_clk_out,
    scan_data_in,
    scan_data_out,
    scan_latch_en,
    scan_select,
    set_clk_div,
    slow_clk,
    active_select,
    driver_sel,
    inputs,
    oeb,
    outputs);
 input clk;
 input la_scan_clk_in;
 input la_scan_data_in;
 output la_scan_data_out;
 input la_scan_latch_en;
 input la_scan_select;
 output ready;
 input reset;
 input scan_clk_in;
 output scan_clk_out;
 input scan_data_in;
 output scan_data_out;
 output scan_latch_en;
 output scan_select;
 input set_clk_div;
 output slow_clk;
 input [8:0] active_select;
 input [1:0] driver_sel;
 input [7:0] inputs;
 output [37:0] oeb;
 output [7:0] outputs;

 wire net43;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net44;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net45;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire active;
 wire \aio_input_reg[0] ;
 wire \aio_input_reg[1] ;
 wire \aio_input_reg[2] ;
 wire \aio_input_reg[3] ;
 wire \aio_input_reg[4] ;
 wire \aio_input_reg[5] ;
 wire \aio_input_reg[6] ;
 wire \aio_input_reg[7] ;
 wire aio_input_sh;
 wire \aio_input_shift[0] ;
 wire \aio_input_shift[1] ;
 wire \aio_input_shift[2] ;
 wire \aio_input_shift[3] ;
 wire \aio_input_shift[4] ;
 wire \aio_input_shift[5] ;
 wire \aio_input_shift[6] ;
 wire \aio_input_shift[7] ;
 wire \aio_input_sync[0] ;
 wire \aio_input_sync[1] ;
 wire \aio_input_sync[2] ;
 wire \aio_input_sync[3] ;
 wire \aio_input_sync[4] ;
 wire \aio_input_sync[5] ;
 wire \aio_input_sync[6] ;
 wire \aio_input_sync[7] ;
 wire aio_output_cap;
 wire \aio_output_reg[0] ;
 wire \aio_output_reg[1] ;
 wire \aio_output_reg[2] ;
 wire \aio_output_reg[3] ;
 wire \aio_output_reg[4] ;
 wire \aio_output_reg[5] ;
 wire \aio_output_reg[6] ;
 wire \aio_output_reg[7] ;
 wire \aio_output_shift[0] ;
 wire \aio_output_shift[1] ;
 wire \aio_output_shift[2] ;
 wire \aio_output_shift[3] ;
 wire \aio_output_shift[4] ;
 wire \aio_output_shift[5] ;
 wire \aio_output_shift[6] ;
 wire \aio_output_shift[7] ;
 wire \bit_cnt[0] ;
 wire \bit_cnt[1] ;
 wire \bit_cnt[2] ;
 wire \bit_cnt[3] ;
 wire \clk_divider_I.active ;
 wire \clk_divider_I.ce ;
 wire \clk_divider_I.compare[0] ;
 wire \clk_divider_I.compare[1] ;
 wire \clk_divider_I.compare[2] ;
 wire \clk_divider_I.compare[3] ;
 wire \clk_divider_I.compare[4] ;
 wire \clk_divider_I.compare[5] ;
 wire \clk_divider_I.compare[6] ;
 wire \clk_divider_I.compare[7] ;
 wire \clk_divider_I.counter[0] ;
 wire \clk_divider_I.counter[1] ;
 wire \clk_divider_I.counter[2] ;
 wire \clk_divider_I.counter[3] ;
 wire \clk_divider_I.counter[4] ;
 wire \clk_divider_I.counter[5] ;
 wire \clk_divider_I.counter[6] ;
 wire \clk_divider_I.counter[7] ;
 wire \clk_divider_I.reset ;
 wire \clk_divider_I.set_now ;
 wire \clk_divider_I.set_sync[0] ;
 wire \clk_divider_I.set_sync[1] ;
 wire clknet_0_clk;
 wire clknet_0_scan_clk_in;
 wire clknet_1_0__leaf_scan_clk_in;
 wire clknet_1_1__leaf_scan_clk_in;
 wire clknet_3_0__leaf_clk;
 wire clknet_3_1__leaf_clk;
 wire clknet_3_2__leaf_clk;
 wire clknet_3_3__leaf_clk;
 wire clknet_3_4__leaf_clk;
 wire clknet_3_5__leaf_clk;
 wire clknet_3_6__leaf_clk;
 wire clknet_3_7__leaf_clk;
 wire int_scan_clk_out;
 wire int_scan_data_out;
 wire int_scan_latch_en;
 wire int_scan_select;
 wire net1;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net2;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net3;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net4;
 wire net40;
 wire net41;
 wire net42;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net9;
 wire net90;
 wire net91;
 wire \proj_cnt[0] ;
 wire \proj_cnt[1] ;
 wire \proj_cnt[2] ;
 wire \proj_cnt[3] ;
 wire \proj_cnt[4] ;
 wire \proj_cnt[5] ;
 wire \proj_cnt[6] ;
 wire \proj_cnt[7] ;
 wire \proj_cnt[8] ;
 wire \rst_shift[0] ;
 wire \rst_shift[1] ;
 wire \state[0] ;
 wire \state[12] ;
 wire \state[13] ;
 wire \state[1] ;
 wire \state[2] ;
 wire \state[3] ;
 wire \state[4] ;
 wire \state[5] ;
 wire \state[6] ;
 wire \state[8] ;
 wire \state[9] ;
 wire \ws_cfg[0] ;
 wire \ws_cfg[1] ;
 wire \ws_cfg[2] ;
 wire \ws_cfg[3] ;
 wire \ws_cfg[4] ;
 wire \ws_cfg[5] ;
 wire \ws_cfg[6] ;
 wire \ws_cfg[7] ;
 wire \ws_cnt[0] ;
 wire \ws_cnt[1] ;
 wire \ws_cnt[2] ;
 wire \ws_cnt[3] ;
 wire \ws_cnt[4] ;
 wire \ws_cnt[5] ;
 wire \ws_cnt[6] ;
 wire \ws_cnt[7] ;
 wire ws_set_now;
 wire \ws_set_sync[0] ;
 wire \ws_set_sync[1] ;
 wire \ws_set_sync[2] ;

 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(_0247_));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(net15));
 sky130_fd_sc_hd__fill_2 FILLER_0_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_158 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_202 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_210 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_216 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_258 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_398 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_471 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_13 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_227 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_238 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_40 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_452 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_78 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_124 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_148 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_180 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_192 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_43 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_66 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_122 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_172 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_298 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_39 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_396 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_471 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_63 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_78 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_124 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_131 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_185 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_242 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_263 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_319 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_376 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_409 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_454 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_87 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_9 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_105 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_201 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_214 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_276 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_329 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_58 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_13 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_135 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_142 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_191 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_267 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_286 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_13 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_204 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_299 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_319 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_341 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_371 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_387 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_455 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_462 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_196 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_208 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_295 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_375 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_402 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_420 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_454 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_87 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_182 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_215 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_264 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_350 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_443 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_467 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_70 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_126 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_144 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_372 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_46 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_64 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_71 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_79 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_117 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_122 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_182 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_32 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_44 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_472 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_91 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_115 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_124 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_182 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_217 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_280 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_320 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_35 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_400 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_42 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_16 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_174 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_182 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_213 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_22 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_28 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_341 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_380 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_66 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_8 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_112 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_208 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_229 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_284 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_36 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_388 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_406 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_56 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_67 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_187 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_196 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_243 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_292 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_344 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_368 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_422 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_92 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_127 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_202 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_214 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_226 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_401 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_471 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_32 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_44 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_471 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_204 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_441 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_17 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_21 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_266 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_272 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_314 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_322 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_398 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_406 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_471 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_62 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_70 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_76 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_155 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_20 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_457 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_471 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_255 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_310 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_368 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_120 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_322 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_471 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_230 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_375 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_402 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_420 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_425 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_471 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_183 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_282 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_385 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_471 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_56 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_118 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_180 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_192 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_204 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_270 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_28 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_347 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_364 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_435 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_458 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_465 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_120 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_242 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_291 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_427 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_431 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_124 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_179 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_266 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_322 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_376 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_454 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_79 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_95 ();
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_56 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_57 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_58 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_59 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_60 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_61 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_62 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_63 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_64 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_65 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_66 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_67 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_68 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_69 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_70 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_71 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_72 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_73 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_74 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_75 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_76 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_77 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_78 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_79 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_80 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_81 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_82 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_83 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_84 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_85 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_86 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_87 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_88 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_89 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_90 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_91 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_92 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_93 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_94 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_95 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_96 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_97 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_98 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_99 ();
 sky130_fd_sc_hd__inv_2 _0421_ (.A(\clk_divider_I.counter[7] ),
    .Y(_0127_));
 sky130_fd_sc_hd__inv_2 _0422_ (.A(\clk_divider_I.counter[5] ),
    .Y(_0128_));
 sky130_fd_sc_hd__inv_2 _0423_ (.A(\clk_divider_I.counter[6] ),
    .Y(_0129_));
 sky130_fd_sc_hd__a22o_1 _0424_ (.A1(_0128_),
    .A2(\clk_divider_I.compare[5] ),
    .B1(\clk_divider_I.compare[6] ),
    .B2(_0129_),
    .X(_0130_));
 sky130_fd_sc_hd__inv_2 _0425_ (.A(\clk_divider_I.counter[1] ),
    .Y(_0131_));
 sky130_fd_sc_hd__inv_2 _0426_ (.A(\clk_divider_I.counter[2] ),
    .Y(_0132_));
 sky130_fd_sc_hd__xor2_1 _0427_ (.A(\clk_divider_I.counter[0] ),
    .B(\clk_divider_I.compare[0] ),
    .X(_0133_));
 sky130_fd_sc_hd__a221o_1 _0428_ (.A1(_0131_),
    .A2(\clk_divider_I.compare[1] ),
    .B1(\clk_divider_I.compare[2] ),
    .B2(_0132_),
    .C1(_0133_),
    .X(_0134_));
 sky130_fd_sc_hd__xnor2_1 _0429_ (.A(\clk_divider_I.counter[3] ),
    .B(\clk_divider_I.compare[3] ),
    .Y(_0135_));
 sky130_fd_sc_hd__o221a_1 _0430_ (.A1(_0131_),
    .A2(\clk_divider_I.compare[1] ),
    .B1(\clk_divider_I.compare[2] ),
    .B2(_0132_),
    .C1(_0135_),
    .X(_0136_));
 sky130_fd_sc_hd__inv_2 _0431_ (.A(\clk_divider_I.compare[4] ),
    .Y(_0137_));
 sky130_fd_sc_hd__o22a_1 _0432_ (.A1(\clk_divider_I.counter[4] ),
    .A2(_0137_),
    .B1(\clk_divider_I.compare[7] ),
    .B2(_0127_),
    .X(_0138_));
 sky130_fd_sc_hd__o2bb2a_1 _0433_ (.A1_N(\clk_divider_I.counter[4] ),
    .A2_N(_0137_),
    .B1(\clk_divider_I.compare[5] ),
    .B2(_0128_),
    .X(_0139_));
 sky130_fd_sc_hd__o211a_1 _0434_ (.A1(_0129_),
    .A2(\clk_divider_I.compare[6] ),
    .B1(_0138_),
    .C1(_0139_),
    .X(_0140_));
 sky130_fd_sc_hd__nand3b_1 _0435_ (.A_N(_0134_),
    .B(_0136_),
    .C(_0140_),
    .Y(_0141_));
 sky130_fd_sc_hd__a211oi_1 _0436_ (.A1(_0127_),
    .A2(\clk_divider_I.compare[7] ),
    .B1(_0130_),
    .C1(_0141_),
    .Y(_0142_));
 sky130_fd_sc_hd__nand2_2 _0437_ (.A(\clk_divider_I.ce ),
    .B(_0142_),
    .Y(_0143_));
 sky130_fd_sc_hd__xnor2_1 _0438_ (.A(net41),
    .B(_0143_),
    .Y(_0144_));
 sky130_fd_sc_hd__clkbuf_1 _0439_ (.A(_0144_),
    .X(_0125_));
 sky130_fd_sc_hd__and3_1 _0440_ (.A(\clk_divider_I.ce ),
    .B(\clk_divider_I.counter[1] ),
    .C(\clk_divider_I.counter[0] ),
    .X(_0145_));
 sky130_fd_sc_hd__inv_2 _0441_ (.A(_0145_),
    .Y(_0146_));
 sky130_fd_sc_hd__nor2_1 _0442_ (.A(_0132_),
    .B(_0146_),
    .Y(_0147_));
 sky130_fd_sc_hd__and3_1 _0443_ (.A(\clk_divider_I.counter[4] ),
    .B(\clk_divider_I.counter[3] ),
    .C(_0147_),
    .X(_0148_));
 sky130_fd_sc_hd__nand2_1 _0444_ (.A(\clk_divider_I.counter[5] ),
    .B(_0148_),
    .Y(_0149_));
 sky130_fd_sc_hd__nor2_1 _0445_ (.A(_0129_),
    .B(_0149_),
    .Y(_0150_));
 sky130_fd_sc_hd__a21boi_1 _0446_ (.A1(\clk_divider_I.counter[7] ),
    .A2(_0150_),
    .B1_N(_0143_),
    .Y(_0151_));
 sky130_fd_sc_hd__o21a_1 _0447_ (.A1(\clk_divider_I.counter[7] ),
    .A2(_0150_),
    .B1(_0151_),
    .X(_0152_));
 sky130_fd_sc_hd__clkbuf_1 _0448_ (.A(_0152_),
    .X(_0124_));
 sky130_fd_sc_hd__a221oi_1 _0449_ (.A1(\clk_divider_I.ce ),
    .A2(_0142_),
    .B1(_0149_),
    .B2(_0129_),
    .C1(_0150_),
    .Y(_0153_));
 sky130_fd_sc_hd__clkbuf_1 _0450_ (.A(_0153_),
    .X(_0123_));
 sky130_fd_sc_hd__or2_1 _0451_ (.A(\clk_divider_I.counter[5] ),
    .B(_0148_),
    .X(_0154_));
 sky130_fd_sc_hd__and3_1 _0452_ (.A(_0143_),
    .B(_0149_),
    .C(_0154_),
    .X(_0155_));
 sky130_fd_sc_hd__clkbuf_1 _0453_ (.A(_0155_),
    .X(_0122_));
 sky130_fd_sc_hd__clkinv_2 _0454_ (.A(_0148_),
    .Y(_0156_));
 sky130_fd_sc_hd__a31o_1 _0455_ (.A1(\clk_divider_I.counter[3] ),
    .A2(\clk_divider_I.counter[2] ),
    .A3(_0145_),
    .B1(\clk_divider_I.counter[4] ),
    .X(_0157_));
 sky130_fd_sc_hd__and3_1 _0456_ (.A(_0143_),
    .B(_0156_),
    .C(_0157_),
    .X(_0158_));
 sky130_fd_sc_hd__clkbuf_1 _0457_ (.A(_0158_),
    .X(_0121_));
 sky130_fd_sc_hd__o21ai_1 _0458_ (.A1(\clk_divider_I.counter[3] ),
    .A2(_0147_),
    .B1(_0143_),
    .Y(_0159_));
 sky130_fd_sc_hd__a21oi_1 _0459_ (.A1(\clk_divider_I.counter[3] ),
    .A2(_0147_),
    .B1(_0159_),
    .Y(_0160_));
 sky130_fd_sc_hd__clkbuf_1 _0460_ (.A(_0160_),
    .X(_0120_));
 sky130_fd_sc_hd__o21ai_1 _0461_ (.A1(\clk_divider_I.counter[2] ),
    .A2(_0145_),
    .B1(_0143_),
    .Y(_0161_));
 sky130_fd_sc_hd__nor2_1 _0462_ (.A(_0147_),
    .B(_0161_),
    .Y(_0162_));
 sky130_fd_sc_hd__clkbuf_1 _0463_ (.A(_0162_),
    .X(_0119_));
 sky130_fd_sc_hd__a21o_1 _0464_ (.A1(\clk_divider_I.ce ),
    .A2(\clk_divider_I.counter[0] ),
    .B1(\clk_divider_I.counter[1] ),
    .X(_0163_));
 sky130_fd_sc_hd__and3_1 _0465_ (.A(_0143_),
    .B(_0146_),
    .C(_0163_),
    .X(_0164_));
 sky130_fd_sc_hd__clkbuf_1 _0466_ (.A(_0164_),
    .X(_0118_));
 sky130_fd_sc_hd__o21ai_1 _0467_ (.A1(\clk_divider_I.ce ),
    .A2(\clk_divider_I.counter[0] ),
    .B1(_0143_),
    .Y(_0165_));
 sky130_fd_sc_hd__a21oi_1 _0468_ (.A1(\clk_divider_I.ce ),
    .A2(\clk_divider_I.counter[0] ),
    .B1(_0165_),
    .Y(_0166_));
 sky130_fd_sc_hd__clkbuf_1 _0469_ (.A(_0166_),
    .X(_0117_));
 sky130_fd_sc_hd__mux2_1 _0470_ (.A0(\ws_cfg[7] ),
    .A1(net19),
    .S(ws_set_now),
    .X(_0167_));
 sky130_fd_sc_hd__clkbuf_1 _0471_ (.A(_0167_),
    .X(_0072_));
 sky130_fd_sc_hd__mux2_1 _0472_ (.A0(\ws_cfg[6] ),
    .A1(net18),
    .S(ws_set_now),
    .X(_0168_));
 sky130_fd_sc_hd__clkbuf_1 _0473_ (.A(_0168_),
    .X(_0071_));
 sky130_fd_sc_hd__mux2_1 _0474_ (.A0(\ws_cfg[5] ),
    .A1(net17),
    .S(ws_set_now),
    .X(_0169_));
 sky130_fd_sc_hd__clkbuf_1 _0475_ (.A(_0169_),
    .X(_0070_));
 sky130_fd_sc_hd__mux2_1 _0476_ (.A0(\ws_cfg[4] ),
    .A1(net16),
    .S(ws_set_now),
    .X(_0170_));
 sky130_fd_sc_hd__clkbuf_1 _0477_ (.A(_0170_),
    .X(_0069_));
 sky130_fd_sc_hd__mux2_1 _0478_ (.A0(\ws_cfg[3] ),
    .A1(net15),
    .S(ws_set_now),
    .X(_0171_));
 sky130_fd_sc_hd__clkbuf_1 _0479_ (.A(_0171_),
    .X(_0068_));
 sky130_fd_sc_hd__mux2_1 _0480_ (.A0(\ws_cfg[2] ),
    .A1(net14),
    .S(ws_set_now),
    .X(_0172_));
 sky130_fd_sc_hd__clkbuf_1 _0481_ (.A(_0172_),
    .X(_0067_));
 sky130_fd_sc_hd__mux2_1 _0482_ (.A0(\ws_cfg[1] ),
    .A1(net13),
    .S(ws_set_now),
    .X(_0173_));
 sky130_fd_sc_hd__clkbuf_1 _0483_ (.A(_0173_),
    .X(_0066_));
 sky130_fd_sc_hd__mux2_1 _0484_ (.A0(\ws_cfg[0] ),
    .A1(net12),
    .S(ws_set_now),
    .X(_0174_));
 sky130_fd_sc_hd__clkbuf_1 _0485_ (.A(_0174_),
    .X(_0065_));
 sky130_fd_sc_hd__clkinv_2 _0486_ (.A(net24),
    .Y(_0175_));
 sky130_fd_sc_hd__clkbuf_1 _0487_ (.A(_0175_),
    .X(_0021_));
 sky130_fd_sc_hd__clkinv_2 _0488_ (.A(net24),
    .Y(_0176_));
 sky130_fd_sc_hd__clkbuf_1 _0489_ (.A(_0176_),
    .X(_0019_));
 sky130_fd_sc_hd__inv_2 _0490_ (.A(net24),
    .Y(_0177_));
 sky130_fd_sc_hd__clkbuf_1 _0491_ (.A(_0177_),
    .X(_0017_));
 sky130_fd_sc_hd__inv_2 _0492_ (.A(\ws_cnt[2] ),
    .Y(_0178_));
 sky130_fd_sc_hd__clkbuf_4 _0493_ (.A(\state[3] ),
    .X(_0179_));
 sky130_fd_sc_hd__mux2_1 _0494_ (.A0(\ws_cfg[3] ),
    .A1(\ws_cfg[2] ),
    .S(_0179_),
    .X(_0180_));
 sky130_fd_sc_hd__nor2_1 _0495_ (.A(_0178_),
    .B(_0180_),
    .Y(_0181_));
 sky130_fd_sc_hd__inv_2 _0496_ (.A(\ws_cnt[3] ),
    .Y(_0182_));
 sky130_fd_sc_hd__mux2_1 _0497_ (.A0(\ws_cfg[4] ),
    .A1(\ws_cfg[3] ),
    .S(_0179_),
    .X(_0183_));
 sky130_fd_sc_hd__mux2_1 _0498_ (.A0(\ws_cfg[6] ),
    .A1(\ws_cfg[5] ),
    .S(_0179_),
    .X(_0184_));
 sky130_fd_sc_hd__inv_2 _0499_ (.A(\ws_cnt[5] ),
    .Y(_0185_));
 sky130_fd_sc_hd__inv_2 _0500_ (.A(\ws_cnt[0] ),
    .Y(_0186_));
 sky130_fd_sc_hd__mux2_1 _0501_ (.A0(\ws_cfg[1] ),
    .A1(\ws_cfg[0] ),
    .S(\state[3] ),
    .X(_0187_));
 sky130_fd_sc_hd__mux2_1 _0502_ (.A0(\ws_cfg[7] ),
    .A1(\ws_cfg[6] ),
    .S(_0179_),
    .X(_0188_));
 sky130_fd_sc_hd__inv_2 _0503_ (.A(\ws_cnt[6] ),
    .Y(_0189_));
 sky130_fd_sc_hd__a22o_1 _0504_ (.A1(_0186_),
    .A2(_0187_),
    .B1(_0188_),
    .B2(_0189_),
    .X(_0190_));
 sky130_fd_sc_hd__a221o_1 _0505_ (.A1(_0182_),
    .A2(_0183_),
    .B1(_0184_),
    .B2(_0185_),
    .C1(_0190_),
    .X(_0191_));
 sky130_fd_sc_hd__nand2_1 _0506_ (.A(\ws_cfg[7] ),
    .B(_0179_),
    .Y(_0192_));
 sky130_fd_sc_hd__nor2_1 _0507_ (.A(\ws_cnt[7] ),
    .B(_0192_),
    .Y(_0193_));
 sky130_fd_sc_hd__a2bb2o_1 _0508_ (.A1_N(_0185_),
    .A2_N(_0184_),
    .B1(_0192_),
    .B2(\ws_cnt[7] ),
    .X(_0194_));
 sky130_fd_sc_hd__mux2_1 _0509_ (.A0(\ws_cfg[2] ),
    .A1(\ws_cfg[1] ),
    .S(_0179_),
    .X(_0195_));
 sky130_fd_sc_hd__inv_2 _0510_ (.A(\ws_cnt[1] ),
    .Y(_0196_));
 sky130_fd_sc_hd__a2bb2o_1 _0511_ (.A1_N(_0186_),
    .A2_N(_0187_),
    .B1(_0195_),
    .B2(_0196_),
    .X(_0197_));
 sky130_fd_sc_hd__or4_1 _0512_ (.A(_0191_),
    .B(_0193_),
    .C(_0194_),
    .D(_0197_),
    .X(_0198_));
 sky130_fd_sc_hd__mux2_1 _0513_ (.A0(\ws_cfg[5] ),
    .A1(\ws_cfg[4] ),
    .S(_0179_),
    .X(_0199_));
 sky130_fd_sc_hd__xor2_1 _0514_ (.A(\ws_cnt[4] ),
    .B(_0199_),
    .X(_0200_));
 sky130_fd_sc_hd__o2bb2a_1 _0515_ (.A1_N(_0178_),
    .A2_N(_0180_),
    .B1(_0195_),
    .B2(_0196_),
    .X(_0201_));
 sky130_fd_sc_hd__o221a_1 _0516_ (.A1(_0182_),
    .A2(_0183_),
    .B1(_0188_),
    .B2(_0189_),
    .C1(_0201_),
    .X(_0202_));
 sky130_fd_sc_hd__or4b_4 _0517_ (.A(_0181_),
    .B(_0198_),
    .C(_0200_),
    .D_N(_0202_),
    .X(_0203_));
 sky130_fd_sc_hd__mux2_1 _0518_ (.A0(\state[1] ),
    .A1(\state[8] ),
    .S(_0203_),
    .X(_0204_));
 sky130_fd_sc_hd__clkbuf_1 _0519_ (.A(_0204_),
    .X(_0056_));
 sky130_fd_sc_hd__a21o_1 _0520_ (.A1(\state[1] ),
    .A2(_0203_),
    .B1(\state[13] ),
    .X(_0205_));
 sky130_fd_sc_hd__clkbuf_1 _0521_ (.A(_0205_),
    .X(_0008_));
 sky130_fd_sc_hd__inv_2 _0522_ (.A(_0203_),
    .Y(_0206_));
 sky130_fd_sc_hd__inv_2 _0523_ (.A(\proj_cnt[2] ),
    .Y(_0207_));
 sky130_fd_sc_hd__clkinv_2 _0524_ (.A(\proj_cnt[0] ),
    .Y(_0208_));
 sky130_fd_sc_hd__and4b_1 _0525_ (.A_N(\proj_cnt[8] ),
    .B(\proj_cnt[7] ),
    .C(\proj_cnt[6] ),
    .D(\proj_cnt[3] ),
    .X(_0209_));
 sky130_fd_sc_hd__and4_1 _0526_ (.A(_0207_),
    .B(\proj_cnt[1] ),
    .C(_0208_),
    .D(_0209_),
    .X(_0210_));
 sky130_fd_sc_hd__and3_1 _0527_ (.A(\proj_cnt[5] ),
    .B(\proj_cnt[4] ),
    .C(_0210_),
    .X(_0211_));
 sky130_fd_sc_hd__nand2_1 _0528_ (.A(net1),
    .B(_0211_),
    .Y(_0212_));
 sky130_fd_sc_hd__xnor2_1 _0529_ (.A(\proj_cnt[4] ),
    .B(net5),
    .Y(_0213_));
 sky130_fd_sc_hd__xnor2_1 _0530_ (.A(\proj_cnt[7] ),
    .B(net8),
    .Y(_0214_));
 sky130_fd_sc_hd__xnor2_1 _0531_ (.A(\proj_cnt[8] ),
    .B(net9),
    .Y(_0215_));
 sky130_fd_sc_hd__inv_2 _0532_ (.A(\proj_cnt[1] ),
    .Y(_0216_));
 sky130_fd_sc_hd__xor2_1 _0533_ (.A(\proj_cnt[3] ),
    .B(net4),
    .X(_0217_));
 sky130_fd_sc_hd__a221o_1 _0534_ (.A1(_0208_),
    .A2(net1),
    .B1(net2),
    .B2(_0216_),
    .C1(_0217_),
    .X(_0218_));
 sky130_fd_sc_hd__xnor2_1 _0535_ (.A(\proj_cnt[2] ),
    .B(net3),
    .Y(_0219_));
 sky130_fd_sc_hd__xnor2_1 _0536_ (.A(\proj_cnt[5] ),
    .B(net6),
    .Y(_0220_));
 sky130_fd_sc_hd__xnor2_1 _0537_ (.A(\proj_cnt[6] ),
    .B(net7),
    .Y(_0221_));
 sky130_fd_sc_hd__o221a_1 _0538_ (.A1(_0208_),
    .A2(net1),
    .B1(net2),
    .B2(_0216_),
    .C1(_0221_),
    .X(_0222_));
 sky130_fd_sc_hd__and4b_1 _0539_ (.A_N(_0218_),
    .B(_0219_),
    .C(_0220_),
    .D(_0222_),
    .X(_0223_));
 sky130_fd_sc_hd__a41o_1 _0540_ (.A1(_0213_),
    .A2(_0214_),
    .A3(_0215_),
    .A4(_0223_),
    .B1(_0208_),
    .X(_0224_));
 sky130_fd_sc_hd__nand2_1 _0541_ (.A(_0212_),
    .B(_0224_),
    .Y(_0225_));
 sky130_fd_sc_hd__and4b_1 _0542_ (.A_N(\bit_cnt[3] ),
    .B(\bit_cnt[2] ),
    .C(\bit_cnt[1] ),
    .D(\bit_cnt[0] ),
    .X(_0226_));
 sky130_fd_sc_hd__or4b_1 _0543_ (.A(\bit_cnt[2] ),
    .B(\bit_cnt[1] ),
    .C(\bit_cnt[0] ),
    .D_N(\bit_cnt[3] ),
    .X(_0227_));
 sky130_fd_sc_hd__a21bo_1 _0544_ (.A1(_0212_),
    .A2(_0224_),
    .B1_N(_0227_),
    .X(_0228_));
 sky130_fd_sc_hd__o21a_2 _0545_ (.A1(_0225_),
    .A2(_0226_),
    .B1(_0228_),
    .X(_0229_));
 sky130_fd_sc_hd__nand2_1 _0546_ (.A(_0211_),
    .B(_0229_),
    .Y(_0230_));
 sky130_fd_sc_hd__a22o_1 _0547_ (.A1(\state[8] ),
    .A2(_0206_),
    .B1(_0230_),
    .B2(\state[12] ),
    .X(_0231_));
 sky130_fd_sc_hd__clkbuf_1 _0548_ (.A(_0231_),
    .X(_0012_));
 sky130_fd_sc_hd__a21o_1 _0549_ (.A1(\state[6] ),
    .A2(_0203_),
    .B1(\state[9] ),
    .X(_0232_));
 sky130_fd_sc_hd__clkbuf_1 _0550_ (.A(_0232_),
    .X(_0013_));
 sky130_fd_sc_hd__inv_2 _0551_ (.A(\clk_divider_I.ce ),
    .Y(_0233_));
 sky130_fd_sc_hd__nand4_1 _0552_ (.A(_0213_),
    .B(_0214_),
    .C(_0215_),
    .D(_0223_),
    .Y(_0234_));
 sky130_fd_sc_hd__inv_2 _0553_ (.A(_0234_),
    .Y(_0235_));
 sky130_fd_sc_hd__nor2_1 _0554_ (.A(\clk_divider_I.ce ),
    .B(aio_input_sh),
    .Y(_0236_));
 sky130_fd_sc_hd__a31oi_1 _0555_ (.A1(_0233_),
    .A2(_0235_),
    .A3(_0229_),
    .B1(_0236_),
    .Y(_0237_));
 sky130_fd_sc_hd__clkbuf_1 _0556_ (.A(_0237_),
    .X(_0011_));
 sky130_fd_sc_hd__a32o_1 _0557_ (.A1(aio_input_sh),
    .A2(_0235_),
    .A3(_0229_),
    .B1(\state[2] ),
    .B2(_0203_),
    .X(_0238_));
 sky130_fd_sc_hd__clkbuf_1 _0558_ (.A(_0238_),
    .X(_0009_));
 sky130_fd_sc_hd__inv_2 _0559_ (.A(active),
    .Y(_0239_));
 sky130_fd_sc_hd__a21o_1 _0560_ (.A1(\state[0] ),
    .A2(_0239_),
    .B1(aio_output_cap),
    .X(_0240_));
 sky130_fd_sc_hd__clkbuf_1 _0561_ (.A(_0240_),
    .X(_0007_));
 sky130_fd_sc_hd__a32o_1 _0562_ (.A1(\state[12] ),
    .A2(_0211_),
    .A3(_0229_),
    .B1(_0203_),
    .B2(_0179_),
    .X(_0241_));
 sky130_fd_sc_hd__clkbuf_1 _0563_ (.A(_0241_),
    .X(_0010_));
 sky130_fd_sc_hd__buf_2 _0564_ (.A(net11),
    .X(_0242_));
 sky130_fd_sc_hd__and2_1 _0565_ (.A(_0242_),
    .B(net10),
    .X(_0243_));
 sky130_fd_sc_hd__clkbuf_1 _0566_ (.A(_0243_),
    .X(_0003_));
 sky130_fd_sc_hd__clkbuf_4 _0567_ (.A(net11),
    .X(_0244_));
 sky130_fd_sc_hd__mux2_2 _0568_ (.A0(clknet_1_1__leaf_scan_clk_in),
    .A1(\aio_output_reg[0] ),
    .S(_0244_),
    .X(_0245_));
 sky130_fd_sc_hd__buf_2 _0569_ (.A(_0245_),
    .X(net28));
 sky130_fd_sc_hd__mux2_1 _0570_ (.A0(net25),
    .A1(\aio_output_reg[1] ),
    .S(_0244_),
    .X(_0246_));
 sky130_fd_sc_hd__clkbuf_1 _0571_ (.A(_0246_),
    .X(net29));
 sky130_fd_sc_hd__and2_1 _0572_ (.A(_0242_),
    .B(\aio_output_reg[2] ),
    .X(_0247_));
 sky130_fd_sc_hd__clkbuf_1 _0573_ (.A(_0247_),
    .X(net30));
 sky130_fd_sc_hd__and2_1 _0574_ (.A(_0242_),
    .B(\aio_output_reg[3] ),
    .X(_0248_));
 sky130_fd_sc_hd__clkbuf_1 _0575_ (.A(_0248_),
    .X(net31));
 sky130_fd_sc_hd__and2_1 _0576_ (.A(_0242_),
    .B(\aio_output_reg[4] ),
    .X(_0249_));
 sky130_fd_sc_hd__clkbuf_1 _0577_ (.A(_0249_),
    .X(net32));
 sky130_fd_sc_hd__and2_1 _0578_ (.A(_0242_),
    .B(\aio_output_reg[5] ),
    .X(_0250_));
 sky130_fd_sc_hd__clkbuf_1 _0579_ (.A(_0250_),
    .X(net33));
 sky130_fd_sc_hd__and2_1 _0580_ (.A(_0242_),
    .B(\aio_output_reg[6] ),
    .X(_0251_));
 sky130_fd_sc_hd__clkbuf_1 _0581_ (.A(_0251_),
    .X(net34));
 sky130_fd_sc_hd__and2_1 _0582_ (.A(_0242_),
    .B(\aio_output_reg[7] ),
    .X(_0252_));
 sky130_fd_sc_hd__clkbuf_1 _0583_ (.A(_0252_),
    .X(net35));
 sky130_fd_sc_hd__mux2_1 _0584_ (.A0(net12),
    .A1(net20),
    .S(net10),
    .X(_0253_));
 sky130_fd_sc_hd__mux2_1 _0585_ (.A0(_0253_),
    .A1(int_scan_clk_out),
    .S(_0244_),
    .X(_0254_));
 sky130_fd_sc_hd__clkbuf_1 _0586_ (.A(_0254_),
    .X(net37));
 sky130_fd_sc_hd__mux2_1 _0587_ (.A0(net13),
    .A1(net21),
    .S(net10),
    .X(_0255_));
 sky130_fd_sc_hd__mux2_1 _0588_ (.A0(_0255_),
    .A1(int_scan_data_out),
    .S(_0244_),
    .X(_0256_));
 sky130_fd_sc_hd__clkbuf_1 _0589_ (.A(_0256_),
    .X(net38));
 sky130_fd_sc_hd__mux2_1 _0590_ (.A0(net14),
    .A1(net23),
    .S(net10),
    .X(_0257_));
 sky130_fd_sc_hd__mux2_1 _0591_ (.A0(_0257_),
    .A1(int_scan_select),
    .S(_0244_),
    .X(_0258_));
 sky130_fd_sc_hd__clkbuf_1 _0592_ (.A(_0258_),
    .X(net40));
 sky130_fd_sc_hd__mux2_1 _0593_ (.A0(net15),
    .A1(net22),
    .S(net10),
    .X(_0259_));
 sky130_fd_sc_hd__mux2_1 _0594_ (.A0(_0259_),
    .A1(int_scan_latch_en),
    .S(net11),
    .X(_0260_));
 sky130_fd_sc_hd__clkbuf_1 _0595_ (.A(_0260_),
    .X(net39));
 sky130_fd_sc_hd__and2_1 _0596_ (.A(\state[6] ),
    .B(_0206_),
    .X(_0261_));
 sky130_fd_sc_hd__clkbuf_1 _0597_ (.A(_0261_),
    .X(_0006_));
 sky130_fd_sc_hd__inv_2 _0598_ (.A(\state[0] ),
    .Y(_0262_));
 sky130_fd_sc_hd__nor2_1 _0599_ (.A(_0262_),
    .B(_0239_),
    .Y(_0263_));
 sky130_fd_sc_hd__clkbuf_2 _0600_ (.A(_0263_),
    .X(net36));
 sky130_fd_sc_hd__and2_1 _0601_ (.A(_0179_),
    .B(_0206_),
    .X(_0264_));
 sky130_fd_sc_hd__clkbuf_1 _0602_ (.A(_0264_),
    .X(_0005_));
 sky130_fd_sc_hd__and2_1 _0603_ (.A(\state[2] ),
    .B(_0206_),
    .X(_0265_));
 sky130_fd_sc_hd__clkbuf_1 _0604_ (.A(_0265_),
    .X(_0004_));
 sky130_fd_sc_hd__or2_1 _0605_ (.A(\state[12] ),
    .B(aio_input_sh),
    .X(_0266_));
 sky130_fd_sc_hd__buf_2 _0606_ (.A(_0266_),
    .X(_0267_));
 sky130_fd_sc_hd__or2_1 _0607_ (.A(\state[13] ),
    .B(_0267_),
    .X(_0268_));
 sky130_fd_sc_hd__clkbuf_1 _0608_ (.A(_0268_),
    .X(_0000_));
 sky130_fd_sc_hd__or3_1 _0609_ (.A(\state[1] ),
    .B(\state[13] ),
    .C(\state[6] ),
    .X(_0269_));
 sky130_fd_sc_hd__clkbuf_1 _0610_ (.A(_0269_),
    .X(_0001_));
 sky130_fd_sc_hd__and2b_1 _0611_ (.A_N(\ws_set_sync[2] ),
    .B(\ws_set_sync[1] ),
    .X(_0270_));
 sky130_fd_sc_hd__clkbuf_1 _0612_ (.A(_0270_),
    .X(_0002_));
 sky130_fd_sc_hd__and2b_1 _0613_ (.A_N(\clk_divider_I.active ),
    .B(\clk_divider_I.set_sync[1] ),
    .X(_0271_));
 sky130_fd_sc_hd__clkbuf_1 _0614_ (.A(_0271_),
    .X(_0014_));
 sky130_fd_sc_hd__buf_4 _0615_ (.A(\clk_divider_I.reset ),
    .X(_0272_));
 sky130_fd_sc_hd__inv_2 _0616_ (.A(_0272_),
    .Y(_0273_));
 sky130_fd_sc_hd__clkbuf_1 _0617_ (.A(_0273_),
    .X(_0015_));
 sky130_fd_sc_hd__clkinv_2 _0618_ (.A(_0272_),
    .Y(_0274_));
 sky130_fd_sc_hd__clkbuf_1 _0619_ (.A(_0274_),
    .X(_0016_));
 sky130_fd_sc_hd__mux2_1 _0620_ (.A0(\clk_divider_I.compare[0] ),
    .A1(net12),
    .S(\clk_divider_I.set_now ),
    .X(_0275_));
 sky130_fd_sc_hd__clkbuf_1 _0621_ (.A(_0275_),
    .X(_0057_));
 sky130_fd_sc_hd__mux2_1 _0622_ (.A0(\clk_divider_I.compare[1] ),
    .A1(net13),
    .S(\clk_divider_I.set_now ),
    .X(_0276_));
 sky130_fd_sc_hd__clkbuf_1 _0623_ (.A(_0276_),
    .X(_0058_));
 sky130_fd_sc_hd__mux2_1 _0624_ (.A0(\clk_divider_I.compare[2] ),
    .A1(net14),
    .S(\clk_divider_I.set_now ),
    .X(_0277_));
 sky130_fd_sc_hd__clkbuf_1 _0625_ (.A(_0277_),
    .X(_0059_));
 sky130_fd_sc_hd__mux2_1 _0626_ (.A0(\clk_divider_I.compare[3] ),
    .A1(net15),
    .S(\clk_divider_I.set_now ),
    .X(_0278_));
 sky130_fd_sc_hd__clkbuf_1 _0627_ (.A(_0278_),
    .X(_0060_));
 sky130_fd_sc_hd__mux2_1 _0628_ (.A0(\clk_divider_I.compare[4] ),
    .A1(net16),
    .S(\clk_divider_I.set_now ),
    .X(_0279_));
 sky130_fd_sc_hd__clkbuf_1 _0629_ (.A(_0279_),
    .X(_0061_));
 sky130_fd_sc_hd__mux2_1 _0630_ (.A0(\clk_divider_I.compare[5] ),
    .A1(net17),
    .S(\clk_divider_I.set_now ),
    .X(_0280_));
 sky130_fd_sc_hd__clkbuf_1 _0631_ (.A(_0280_),
    .X(_0062_));
 sky130_fd_sc_hd__mux2_1 _0632_ (.A0(\clk_divider_I.compare[6] ),
    .A1(net18),
    .S(\clk_divider_I.set_now ),
    .X(_0281_));
 sky130_fd_sc_hd__clkbuf_1 _0633_ (.A(_0281_),
    .X(_0063_));
 sky130_fd_sc_hd__mux2_1 _0634_ (.A0(\clk_divider_I.compare[7] ),
    .A1(net19),
    .S(\clk_divider_I.set_now ),
    .X(_0282_));
 sky130_fd_sc_hd__clkbuf_1 _0635_ (.A(_0282_),
    .X(_0064_));
 sky130_fd_sc_hd__inv_2 _0636__1 (.A(clknet_3_0__leaf_clk),
    .Y(net81));
 sky130_fd_sc_hd__buf_2 _0637_ (.A(net81),
    .X(_0018_));
 sky130_fd_sc_hd__inv_2 _0638__2 (.A(clknet_3_1__leaf_clk),
    .Y(net82));
 sky130_fd_sc_hd__buf_2 _0639_ (.A(net82),
    .X(_0020_));
 sky130_fd_sc_hd__inv_2 _0640__3 (.A(clknet_3_1__leaf_clk),
    .Y(net83));
 sky130_fd_sc_hd__buf_2 _0641_ (.A(net83),
    .X(_0022_));
 sky130_fd_sc_hd__clkinv_2 _0642_ (.A(_0272_),
    .Y(_0286_));
 sky130_fd_sc_hd__clkbuf_1 _0643_ (.A(_0286_),
    .X(_0023_));
 sky130_fd_sc_hd__inv_2 _0644_ (.A(_0272_),
    .Y(_0287_));
 sky130_fd_sc_hd__clkbuf_1 _0645_ (.A(_0287_),
    .X(_0024_));
 sky130_fd_sc_hd__clkinv_2 _0646_ (.A(_0272_),
    .Y(_0288_));
 sky130_fd_sc_hd__clkbuf_1 _0647_ (.A(_0288_),
    .X(_0025_));
 sky130_fd_sc_hd__inv_2 _0648_ (.A(_0272_),
    .Y(_0289_));
 sky130_fd_sc_hd__clkbuf_1 _0649_ (.A(_0289_),
    .X(_0026_));
 sky130_fd_sc_hd__clkinv_2 _0650_ (.A(_0272_),
    .Y(_0290_));
 sky130_fd_sc_hd__clkbuf_1 _0651_ (.A(_0290_),
    .X(_0027_));
 sky130_fd_sc_hd__clkinv_2 _0652_ (.A(_0272_),
    .Y(_0291_));
 sky130_fd_sc_hd__clkbuf_1 _0653_ (.A(_0291_),
    .X(_0028_));
 sky130_fd_sc_hd__inv_2 _0654_ (.A(_0272_),
    .Y(_0292_));
 sky130_fd_sc_hd__clkbuf_1 _0655_ (.A(_0292_),
    .X(_0029_));
 sky130_fd_sc_hd__inv_2 _0656_ (.A(_0272_),
    .Y(_0293_));
 sky130_fd_sc_hd__clkbuf_1 _0657_ (.A(_0293_),
    .X(_0030_));
 sky130_fd_sc_hd__clkbuf_8 _0658_ (.A(\clk_divider_I.reset ),
    .X(_0294_));
 sky130_fd_sc_hd__inv_2 _0659_ (.A(_0294_),
    .Y(_0295_));
 sky130_fd_sc_hd__clkbuf_1 _0660_ (.A(_0295_),
    .X(_0031_));
 sky130_fd_sc_hd__clkinv_2 _0661_ (.A(_0294_),
    .Y(_0296_));
 sky130_fd_sc_hd__clkbuf_1 _0662_ (.A(_0296_),
    .X(_0032_));
 sky130_fd_sc_hd__clkinv_2 _0663_ (.A(_0294_),
    .Y(_0297_));
 sky130_fd_sc_hd__clkbuf_1 _0664_ (.A(_0297_),
    .X(_0033_));
 sky130_fd_sc_hd__inv_2 _0665_ (.A(_0294_),
    .Y(_0298_));
 sky130_fd_sc_hd__clkbuf_1 _0666_ (.A(_0298_),
    .X(_0034_));
 sky130_fd_sc_hd__inv_2 _0667_ (.A(_0294_),
    .Y(_0299_));
 sky130_fd_sc_hd__clkbuf_1 _0668_ (.A(_0299_),
    .X(_0035_));
 sky130_fd_sc_hd__clkinv_2 _0669_ (.A(_0294_),
    .Y(_0300_));
 sky130_fd_sc_hd__clkbuf_1 _0670_ (.A(_0300_),
    .X(_0036_));
 sky130_fd_sc_hd__clkinv_2 _0671_ (.A(_0294_),
    .Y(_0301_));
 sky130_fd_sc_hd__clkbuf_1 _0672_ (.A(_0301_),
    .X(_0037_));
 sky130_fd_sc_hd__inv_2 _0673_ (.A(_0294_),
    .Y(_0302_));
 sky130_fd_sc_hd__clkbuf_1 _0674_ (.A(_0302_),
    .X(_0038_));
 sky130_fd_sc_hd__inv_2 _0675_ (.A(_0294_),
    .Y(_0303_));
 sky130_fd_sc_hd__clkbuf_1 _0676_ (.A(_0303_),
    .X(_0039_));
 sky130_fd_sc_hd__inv_2 _0677_ (.A(_0294_),
    .Y(_0304_));
 sky130_fd_sc_hd__clkbuf_1 _0678_ (.A(_0304_),
    .X(_0040_));
 sky130_fd_sc_hd__buf_4 _0679_ (.A(\clk_divider_I.reset ),
    .X(_0305_));
 sky130_fd_sc_hd__inv_2 _0680_ (.A(_0305_),
    .Y(_0306_));
 sky130_fd_sc_hd__clkbuf_1 _0681_ (.A(_0306_),
    .X(_0041_));
 sky130_fd_sc_hd__clkinv_2 _0682_ (.A(_0305_),
    .Y(_0307_));
 sky130_fd_sc_hd__clkbuf_1 _0683_ (.A(_0307_),
    .X(_0042_));
 sky130_fd_sc_hd__inv_2 _0684_ (.A(_0305_),
    .Y(_0308_));
 sky130_fd_sc_hd__clkbuf_1 _0685_ (.A(_0308_),
    .X(_0043_));
 sky130_fd_sc_hd__mux2_1 _0686_ (.A0(\aio_input_shift[1] ),
    .A1(\aio_input_shift[0] ),
    .S(aio_input_sh),
    .X(_0309_));
 sky130_fd_sc_hd__mux2_1 _0687_ (.A0(\aio_input_reg[1] ),
    .A1(_0309_),
    .S(_0233_),
    .X(_0310_));
 sky130_fd_sc_hd__clkbuf_1 _0688_ (.A(_0310_),
    .X(_0073_));
 sky130_fd_sc_hd__mux2_1 _0689_ (.A0(\aio_input_shift[2] ),
    .A1(\aio_input_shift[1] ),
    .S(aio_input_sh),
    .X(_0311_));
 sky130_fd_sc_hd__mux2_1 _0690_ (.A0(\aio_input_reg[2] ),
    .A1(_0311_),
    .S(_0233_),
    .X(_0312_));
 sky130_fd_sc_hd__clkbuf_1 _0691_ (.A(_0312_),
    .X(_0074_));
 sky130_fd_sc_hd__mux2_1 _0692_ (.A0(\aio_input_shift[3] ),
    .A1(\aio_input_shift[2] ),
    .S(aio_input_sh),
    .X(_0313_));
 sky130_fd_sc_hd__mux2_1 _0693_ (.A0(\aio_input_reg[3] ),
    .A1(_0313_),
    .S(_0233_),
    .X(_0314_));
 sky130_fd_sc_hd__clkbuf_1 _0694_ (.A(_0314_),
    .X(_0075_));
 sky130_fd_sc_hd__mux2_1 _0695_ (.A0(\aio_input_shift[4] ),
    .A1(\aio_input_shift[3] ),
    .S(aio_input_sh),
    .X(_0315_));
 sky130_fd_sc_hd__mux2_1 _0696_ (.A0(\aio_input_reg[4] ),
    .A1(_0315_),
    .S(_0233_),
    .X(_0316_));
 sky130_fd_sc_hd__clkbuf_1 _0697_ (.A(_0316_),
    .X(_0076_));
 sky130_fd_sc_hd__mux2_1 _0698_ (.A0(\aio_input_shift[5] ),
    .A1(\aio_input_shift[4] ),
    .S(aio_input_sh),
    .X(_0317_));
 sky130_fd_sc_hd__mux2_1 _0699_ (.A0(\aio_input_reg[5] ),
    .A1(_0317_),
    .S(_0233_),
    .X(_0318_));
 sky130_fd_sc_hd__clkbuf_1 _0700_ (.A(_0318_),
    .X(_0077_));
 sky130_fd_sc_hd__mux2_1 _0701_ (.A0(\aio_input_shift[6] ),
    .A1(\aio_input_shift[5] ),
    .S(aio_input_sh),
    .X(_0319_));
 sky130_fd_sc_hd__mux2_1 _0702_ (.A0(\aio_input_reg[6] ),
    .A1(_0319_),
    .S(_0233_),
    .X(_0320_));
 sky130_fd_sc_hd__clkbuf_1 _0703_ (.A(_0320_),
    .X(_0078_));
 sky130_fd_sc_hd__mux2_1 _0704_ (.A0(\aio_input_shift[7] ),
    .A1(\aio_input_shift[6] ),
    .S(aio_input_sh),
    .X(_0321_));
 sky130_fd_sc_hd__mux2_1 _0705_ (.A0(\aio_input_reg[7] ),
    .A1(_0321_),
    .S(_0233_),
    .X(_0322_));
 sky130_fd_sc_hd__clkbuf_1 _0706_ (.A(_0322_),
    .X(_0079_));
 sky130_fd_sc_hd__o211ai_1 _0707_ (.A1(_0225_),
    .A2(_0226_),
    .B1(_0228_),
    .C1(_0266_),
    .Y(_0323_));
 sky130_fd_sc_hd__buf_2 _0708_ (.A(_0323_),
    .X(_0324_));
 sky130_fd_sc_hd__a21oi_1 _0709_ (.A1(\bit_cnt[0] ),
    .A2(_0267_),
    .B1(\state[0] ),
    .Y(_0325_));
 sky130_fd_sc_hd__o211a_1 _0710_ (.A1(\bit_cnt[0] ),
    .A2(_0267_),
    .B1(_0324_),
    .C1(_0325_),
    .X(_0326_));
 sky130_fd_sc_hd__clkbuf_1 _0711_ (.A(_0326_),
    .X(_0080_));
 sky130_fd_sc_hd__a21oi_1 _0712_ (.A1(\bit_cnt[0] ),
    .A2(_0267_),
    .B1(\bit_cnt[1] ),
    .Y(_0327_));
 sky130_fd_sc_hd__and3_1 _0713_ (.A(\bit_cnt[1] ),
    .B(\bit_cnt[0] ),
    .C(_0266_),
    .X(_0328_));
 sky130_fd_sc_hd__nor3_1 _0714_ (.A(\state[0] ),
    .B(_0327_),
    .C(_0328_),
    .Y(_0329_));
 sky130_fd_sc_hd__clkbuf_1 _0715_ (.A(_0329_),
    .X(_0081_));
 sky130_fd_sc_hd__and2_1 _0716_ (.A(\bit_cnt[2] ),
    .B(_0328_),
    .X(_0330_));
 sky130_fd_sc_hd__nor2_1 _0717_ (.A(\state[0] ),
    .B(_0330_),
    .Y(_0331_));
 sky130_fd_sc_hd__o21a_1 _0718_ (.A1(\bit_cnt[2] ),
    .A2(_0328_),
    .B1(_0331_),
    .X(_0332_));
 sky130_fd_sc_hd__clkbuf_1 _0719_ (.A(_0332_),
    .X(_0082_));
 sky130_fd_sc_hd__nand2_1 _0720_ (.A(\bit_cnt[3] ),
    .B(_0330_),
    .Y(_0333_));
 sky130_fd_sc_hd__or2_1 _0721_ (.A(\bit_cnt[3] ),
    .B(_0330_),
    .X(_0334_));
 sky130_fd_sc_hd__and4_1 _0722_ (.A(_0262_),
    .B(_0324_),
    .C(_0333_),
    .D(_0334_),
    .X(_0335_));
 sky130_fd_sc_hd__clkbuf_1 _0723_ (.A(_0335_),
    .X(_0083_));
 sky130_fd_sc_hd__o21ai_1 _0724_ (.A1(_0208_),
    .A2(_0324_),
    .B1(_0262_),
    .Y(_0336_));
 sky130_fd_sc_hd__a21oi_1 _0725_ (.A1(_0208_),
    .A2(_0324_),
    .B1(_0336_),
    .Y(_0337_));
 sky130_fd_sc_hd__clkbuf_1 _0726_ (.A(_0337_),
    .X(_0084_));
 sky130_fd_sc_hd__and2_1 _0727_ (.A(_0229_),
    .B(_0267_),
    .X(_0338_));
 sky130_fd_sc_hd__nor2_1 _0728_ (.A(_0216_),
    .B(_0208_),
    .Y(_0339_));
 sky130_fd_sc_hd__o21a_1 _0729_ (.A1(_0208_),
    .A2(_0324_),
    .B1(_0216_),
    .X(_0340_));
 sky130_fd_sc_hd__a211oi_1 _0730_ (.A1(_0338_),
    .A2(_0339_),
    .B1(_0340_),
    .C1(\state[0] ),
    .Y(_0341_));
 sky130_fd_sc_hd__clkbuf_1 _0731_ (.A(_0341_),
    .X(_0085_));
 sky130_fd_sc_hd__o31a_1 _0732_ (.A1(_0216_),
    .A2(_0208_),
    .A3(_0324_),
    .B1(_0207_),
    .X(_0342_));
 sky130_fd_sc_hd__or3b_1 _0733_ (.A(_0207_),
    .B(_0323_),
    .C_N(_0339_),
    .X(_0343_));
 sky130_fd_sc_hd__nor3b_1 _0734_ (.A(\state[0] ),
    .B(_0342_),
    .C_N(_0343_),
    .Y(_0344_));
 sky130_fd_sc_hd__clkbuf_1 _0735_ (.A(_0344_),
    .X(_0086_));
 sky130_fd_sc_hd__inv_2 _0736_ (.A(\proj_cnt[3] ),
    .Y(_0345_));
 sky130_fd_sc_hd__and3_1 _0737_ (.A(\proj_cnt[3] ),
    .B(\proj_cnt[2] ),
    .C(_0339_),
    .X(_0346_));
 sky130_fd_sc_hd__a221oi_1 _0738_ (.A1(_0345_),
    .A2(_0343_),
    .B1(_0346_),
    .B2(_0338_),
    .C1(\state[0] ),
    .Y(_0347_));
 sky130_fd_sc_hd__clkbuf_1 _0739_ (.A(_0347_),
    .X(_0087_));
 sky130_fd_sc_hd__a31oi_1 _0740_ (.A1(_0229_),
    .A2(_0267_),
    .A3(_0346_),
    .B1(\proj_cnt[4] ),
    .Y(_0348_));
 sky130_fd_sc_hd__a41o_1 _0741_ (.A1(\proj_cnt[4] ),
    .A2(_0229_),
    .A3(_0267_),
    .A4(_0346_),
    .B1(\state[0] ),
    .X(_0349_));
 sky130_fd_sc_hd__nor2_1 _0742_ (.A(_0348_),
    .B(_0349_),
    .Y(_0350_));
 sky130_fd_sc_hd__clkbuf_1 _0743_ (.A(_0350_),
    .X(_0088_));
 sky130_fd_sc_hd__and3_1 _0744_ (.A(\proj_cnt[5] ),
    .B(\proj_cnt[4] ),
    .C(_0346_),
    .X(_0351_));
 sky130_fd_sc_hd__inv_2 _0745_ (.A(_0351_),
    .Y(_0352_));
 sky130_fd_sc_hd__a41o_1 _0746_ (.A1(\proj_cnt[4] ),
    .A2(_0229_),
    .A3(_0267_),
    .A4(_0346_),
    .B1(\proj_cnt[5] ),
    .X(_0353_));
 sky130_fd_sc_hd__o211a_1 _0747_ (.A1(_0324_),
    .A2(_0352_),
    .B1(_0353_),
    .C1(_0262_),
    .X(_0354_));
 sky130_fd_sc_hd__clkbuf_1 _0748_ (.A(_0354_),
    .X(_0089_));
 sky130_fd_sc_hd__o21ba_1 _0749_ (.A1(_0324_),
    .A2(_0352_),
    .B1_N(\proj_cnt[6] ),
    .X(_0355_));
 sky130_fd_sc_hd__a41o_1 _0750_ (.A1(\proj_cnt[6] ),
    .A2(_0229_),
    .A3(_0267_),
    .A4(_0351_),
    .B1(\state[0] ),
    .X(_0356_));
 sky130_fd_sc_hd__nor2_1 _0751_ (.A(_0355_),
    .B(_0356_),
    .Y(_0357_));
 sky130_fd_sc_hd__clkbuf_1 _0752_ (.A(_0357_),
    .X(_0090_));
 sky130_fd_sc_hd__and3_1 _0753_ (.A(\proj_cnt[7] ),
    .B(\proj_cnt[6] ),
    .C(_0351_),
    .X(_0358_));
 sky130_fd_sc_hd__inv_2 _0754_ (.A(_0358_),
    .Y(_0359_));
 sky130_fd_sc_hd__a41o_1 _0755_ (.A1(\proj_cnt[6] ),
    .A2(_0229_),
    .A3(_0267_),
    .A4(_0351_),
    .B1(\proj_cnt[7] ),
    .X(_0360_));
 sky130_fd_sc_hd__o211a_1 _0756_ (.A1(_0324_),
    .A2(_0359_),
    .B1(_0360_),
    .C1(_0262_),
    .X(_0361_));
 sky130_fd_sc_hd__clkbuf_1 _0757_ (.A(_0361_),
    .X(_0091_));
 sky130_fd_sc_hd__inv_2 _0758_ (.A(\proj_cnt[8] ),
    .Y(_0362_));
 sky130_fd_sc_hd__o21ai_1 _0759_ (.A1(_0324_),
    .A2(_0359_),
    .B1(_0362_),
    .Y(_0363_));
 sky130_fd_sc_hd__or3_1 _0760_ (.A(_0362_),
    .B(_0323_),
    .C(_0359_),
    .X(_0364_));
 sky130_fd_sc_hd__and3_1 _0761_ (.A(_0262_),
    .B(_0363_),
    .C(_0364_),
    .X(_0365_));
 sky130_fd_sc_hd__clkbuf_1 _0762_ (.A(_0365_),
    .X(_0092_));
 sky130_fd_sc_hd__and2_1 _0763_ (.A(_0242_),
    .B(\aio_input_sync[0] ),
    .X(_0366_));
 sky130_fd_sc_hd__clkbuf_1 _0764_ (.A(_0366_),
    .X(_0093_));
 sky130_fd_sc_hd__and2_1 _0765_ (.A(_0242_),
    .B(\aio_input_sync[1] ),
    .X(_0367_));
 sky130_fd_sc_hd__clkbuf_1 _0766_ (.A(_0367_),
    .X(_0094_));
 sky130_fd_sc_hd__and2_1 _0767_ (.A(_0242_),
    .B(\aio_input_sync[2] ),
    .X(_0368_));
 sky130_fd_sc_hd__clkbuf_1 _0768_ (.A(_0368_),
    .X(_0095_));
 sky130_fd_sc_hd__and2_1 _0769_ (.A(_0244_),
    .B(\aio_input_sync[3] ),
    .X(_0369_));
 sky130_fd_sc_hd__clkbuf_1 _0770_ (.A(_0369_),
    .X(_0096_));
 sky130_fd_sc_hd__and2_1 _0771_ (.A(_0244_),
    .B(\aio_input_sync[4] ),
    .X(_0370_));
 sky130_fd_sc_hd__clkbuf_1 _0772_ (.A(_0370_),
    .X(_0097_));
 sky130_fd_sc_hd__and2_1 _0773_ (.A(_0244_),
    .B(\aio_input_sync[5] ),
    .X(_0371_));
 sky130_fd_sc_hd__clkbuf_1 _0774_ (.A(_0371_),
    .X(_0098_));
 sky130_fd_sc_hd__and2_1 _0775_ (.A(_0244_),
    .B(\aio_input_sync[6] ),
    .X(_0372_));
 sky130_fd_sc_hd__clkbuf_1 _0776_ (.A(_0372_),
    .X(_0099_));
 sky130_fd_sc_hd__and2_1 _0777_ (.A(_0244_),
    .B(\aio_input_sync[7] ),
    .X(_0373_));
 sky130_fd_sc_hd__clkbuf_1 _0778_ (.A(_0373_),
    .X(_0100_));
 sky130_fd_sc_hd__mux2_1 _0779_ (.A0(\aio_output_reg[0] ),
    .A1(net87),
    .S(aio_output_cap),
    .X(_0374_));
 sky130_fd_sc_hd__clkbuf_1 _0780_ (.A(_0374_),
    .X(_0101_));
 sky130_fd_sc_hd__mux2_1 _0781_ (.A0(\aio_output_reg[1] ),
    .A1(net90),
    .S(aio_output_cap),
    .X(_0375_));
 sky130_fd_sc_hd__clkbuf_1 _0782_ (.A(_0375_),
    .X(_0102_));
 sky130_fd_sc_hd__mux2_1 _0783_ (.A0(\aio_output_reg[2] ),
    .A1(net91),
    .S(aio_output_cap),
    .X(_0376_));
 sky130_fd_sc_hd__clkbuf_1 _0784_ (.A(_0376_),
    .X(_0103_));
 sky130_fd_sc_hd__mux2_1 _0785_ (.A0(\aio_output_reg[3] ),
    .A1(net86),
    .S(aio_output_cap),
    .X(_0377_));
 sky130_fd_sc_hd__clkbuf_1 _0786_ (.A(_0377_),
    .X(_0104_));
 sky130_fd_sc_hd__mux2_1 _0787_ (.A0(\aio_output_reg[4] ),
    .A1(net89),
    .S(aio_output_cap),
    .X(_0378_));
 sky130_fd_sc_hd__clkbuf_1 _0788_ (.A(_0378_),
    .X(_0105_));
 sky130_fd_sc_hd__mux2_1 _0789_ (.A0(\aio_output_reg[5] ),
    .A1(net85),
    .S(aio_output_cap),
    .X(_0379_));
 sky130_fd_sc_hd__clkbuf_1 _0790_ (.A(_0379_),
    .X(_0106_));
 sky130_fd_sc_hd__mux2_1 _0791_ (.A0(\aio_output_reg[6] ),
    .A1(net88),
    .S(aio_output_cap),
    .X(_0380_));
 sky130_fd_sc_hd__clkbuf_1 _0792_ (.A(_0380_),
    .X(_0107_));
 sky130_fd_sc_hd__mux2_1 _0793_ (.A0(\aio_output_reg[7] ),
    .A1(net84),
    .S(aio_output_cap),
    .X(_0381_));
 sky130_fd_sc_hd__clkbuf_1 _0794_ (.A(_0381_),
    .X(_0108_));
 sky130_fd_sc_hd__inv_2 _0795_ (.A(_0305_),
    .Y(_0382_));
 sky130_fd_sc_hd__clkbuf_1 _0796_ (.A(_0382_),
    .X(_0044_));
 sky130_fd_sc_hd__clkinv_2 _0797_ (.A(_0305_),
    .Y(_0383_));
 sky130_fd_sc_hd__clkbuf_1 _0798_ (.A(_0383_),
    .X(_0045_));
 sky130_fd_sc_hd__clkinv_2 _0799_ (.A(_0305_),
    .Y(_0384_));
 sky130_fd_sc_hd__clkbuf_1 _0800_ (.A(_0384_),
    .X(_0046_));
 sky130_fd_sc_hd__or4_1 _0801_ (.A(\state[1] ),
    .B(_0179_),
    .C(\state[6] ),
    .D(\state[2] ),
    .X(_0385_));
 sky130_fd_sc_hd__o21a_2 _0802_ (.A1(\state[8] ),
    .A2(_0385_),
    .B1(_0203_),
    .X(_0386_));
 sky130_fd_sc_hd__and2_1 _0803_ (.A(_0186_),
    .B(_0386_),
    .X(_0387_));
 sky130_fd_sc_hd__clkbuf_1 _0804_ (.A(_0387_),
    .X(_0109_));
 sky130_fd_sc_hd__or2_1 _0805_ (.A(\ws_cnt[0] ),
    .B(\ws_cnt[1] ),
    .X(_0388_));
 sky130_fd_sc_hd__nand2_1 _0806_ (.A(\ws_cnt[0] ),
    .B(\ws_cnt[1] ),
    .Y(_0389_));
 sky130_fd_sc_hd__and3_1 _0807_ (.A(_0386_),
    .B(_0388_),
    .C(_0389_),
    .X(_0390_));
 sky130_fd_sc_hd__clkbuf_1 _0808_ (.A(_0390_),
    .X(_0110_));
 sky130_fd_sc_hd__nor2_1 _0809_ (.A(_0178_),
    .B(_0389_),
    .Y(_0391_));
 sky130_fd_sc_hd__nand2_1 _0810_ (.A(_0178_),
    .B(_0389_),
    .Y(_0392_));
 sky130_fd_sc_hd__and3b_1 _0811_ (.A_N(_0391_),
    .B(_0392_),
    .C(_0386_),
    .X(_0393_));
 sky130_fd_sc_hd__clkbuf_1 _0812_ (.A(_0393_),
    .X(_0111_));
 sky130_fd_sc_hd__and2_1 _0813_ (.A(\ws_cnt[3] ),
    .B(_0391_),
    .X(_0394_));
 sky130_fd_sc_hd__or2_1 _0814_ (.A(\ws_cnt[3] ),
    .B(_0391_),
    .X(_0395_));
 sky130_fd_sc_hd__and3b_1 _0815_ (.A_N(_0394_),
    .B(_0395_),
    .C(_0386_),
    .X(_0396_));
 sky130_fd_sc_hd__clkbuf_1 _0816_ (.A(_0396_),
    .X(_0112_));
 sky130_fd_sc_hd__and3_1 _0817_ (.A(\ws_cnt[3] ),
    .B(\ws_cnt[4] ),
    .C(_0391_),
    .X(_0397_));
 sky130_fd_sc_hd__o21ai_1 _0818_ (.A1(\ws_cnt[4] ),
    .A2(_0394_),
    .B1(_0386_),
    .Y(_0398_));
 sky130_fd_sc_hd__nor2_1 _0819_ (.A(_0397_),
    .B(_0398_),
    .Y(_0399_));
 sky130_fd_sc_hd__clkbuf_1 _0820_ (.A(_0399_),
    .X(_0113_));
 sky130_fd_sc_hd__and3_1 _0821_ (.A(\ws_cnt[4] ),
    .B(\ws_cnt[5] ),
    .C(_0394_),
    .X(_0400_));
 sky130_fd_sc_hd__o21ai_1 _0822_ (.A1(\ws_cnt[5] ),
    .A2(_0397_),
    .B1(_0386_),
    .Y(_0401_));
 sky130_fd_sc_hd__nor2_1 _0823_ (.A(_0400_),
    .B(_0401_),
    .Y(_0402_));
 sky130_fd_sc_hd__clkbuf_1 _0824_ (.A(_0402_),
    .X(_0114_));
 sky130_fd_sc_hd__nand2_1 _0825_ (.A(\ws_cnt[6] ),
    .B(_0400_),
    .Y(_0403_));
 sky130_fd_sc_hd__or2_1 _0826_ (.A(\ws_cnt[6] ),
    .B(_0400_),
    .X(_0404_));
 sky130_fd_sc_hd__and3_1 _0827_ (.A(_0386_),
    .B(_0403_),
    .C(_0404_),
    .X(_0405_));
 sky130_fd_sc_hd__clkbuf_1 _0828_ (.A(_0405_),
    .X(_0115_));
 sky130_fd_sc_hd__nor2_1 _0829_ (.A(\ws_cnt[7] ),
    .B(_0403_),
    .Y(_0406_));
 sky130_fd_sc_hd__and2_1 _0830_ (.A(\ws_cnt[7] ),
    .B(_0403_),
    .X(_0407_));
 sky130_fd_sc_hd__o21a_1 _0831_ (.A1(_0406_),
    .A2(_0407_),
    .B1(_0386_),
    .X(_0408_));
 sky130_fd_sc_hd__clkbuf_1 _0832_ (.A(_0408_),
    .X(_0116_));
 sky130_fd_sc_hd__clkinv_2 _0833_ (.A(_0305_),
    .Y(_0409_));
 sky130_fd_sc_hd__clkbuf_1 _0834_ (.A(_0409_),
    .X(_0047_));
 sky130_fd_sc_hd__clkinv_2 _0835_ (.A(_0305_),
    .Y(_0410_));
 sky130_fd_sc_hd__clkbuf_1 _0836_ (.A(_0410_),
    .X(_0048_));
 sky130_fd_sc_hd__clkinv_2 _0837_ (.A(_0305_),
    .Y(_0411_));
 sky130_fd_sc_hd__clkbuf_1 _0838_ (.A(_0411_),
    .X(_0049_));
 sky130_fd_sc_hd__inv_2 _0839_ (.A(_0305_),
    .Y(_0412_));
 sky130_fd_sc_hd__clkbuf_1 _0840_ (.A(_0412_),
    .X(_0050_));
 sky130_fd_sc_hd__clkinv_2 _0841_ (.A(\clk_divider_I.reset ),
    .Y(_0413_));
 sky130_fd_sc_hd__clkbuf_1 _0842_ (.A(_0413_),
    .X(_0051_));
 sky130_fd_sc_hd__clkinv_2 _0843_ (.A(\clk_divider_I.reset ),
    .Y(_0414_));
 sky130_fd_sc_hd__clkbuf_1 _0844_ (.A(_0414_),
    .X(_0052_));
 sky130_fd_sc_hd__clkinv_2 _0845_ (.A(\clk_divider_I.reset ),
    .Y(_0415_));
 sky130_fd_sc_hd__clkbuf_1 _0846_ (.A(_0415_),
    .X(_0053_));
 sky130_fd_sc_hd__clkinv_2 _0847_ (.A(\clk_divider_I.reset ),
    .Y(_0416_));
 sky130_fd_sc_hd__clkbuf_1 _0848_ (.A(_0416_),
    .X(_0054_));
 sky130_fd_sc_hd__inv_2 _0849_ (.A(\clk_divider_I.reset ),
    .Y(_0417_));
 sky130_fd_sc_hd__clkbuf_1 _0850_ (.A(_0417_),
    .X(_0055_));
 sky130_fd_sc_hd__mux2_1 _0851_ (.A0(\aio_input_reg[0] ),
    .A1(net41),
    .S(\clk_divider_I.active ),
    .X(_0418_));
 sky130_fd_sc_hd__a22o_1 _0852_ (.A1(\aio_input_shift[0] ),
    .A2(_0236_),
    .B1(_0418_),
    .B2(\clk_divider_I.ce ),
    .X(_0419_));
 sky130_fd_sc_hd__clkbuf_1 _0853_ (.A(_0419_),
    .X(_0126_));
 sky130_fd_sc_hd__dfrtp_1 _0854_ (.CLK(clknet_3_7__leaf_clk),
    .D(_0056_),
    .RESET_B(_0015_),
    .Q(\state[8] ));
 sky130_fd_sc_hd__dfrtp_1 _0855_ (.CLK(clknet_3_4__leaf_clk),
    .D(net11),
    .RESET_B(_0016_),
    .Q(active));
 sky130_fd_sc_hd__dfxtp_1 _0856_ (.CLK(clknet_3_1__leaf_clk),
    .D(_0057_),
    .Q(\clk_divider_I.compare[0] ));
 sky130_fd_sc_hd__dfxtp_1 _0857_ (.CLK(clknet_3_1__leaf_clk),
    .D(_0058_),
    .Q(\clk_divider_I.compare[1] ));
 sky130_fd_sc_hd__dfxtp_1 _0858_ (.CLK(clknet_3_1__leaf_clk),
    .D(_0059_),
    .Q(\clk_divider_I.compare[2] ));
 sky130_fd_sc_hd__dfxtp_1 _0859_ (.CLK(clknet_3_3__leaf_clk),
    .D(_0060_),
    .Q(\clk_divider_I.compare[3] ));
 sky130_fd_sc_hd__dfxtp_1 _0860_ (.CLK(clknet_3_1__leaf_clk),
    .D(_0061_),
    .Q(\clk_divider_I.compare[4] ));
 sky130_fd_sc_hd__dfxtp_1 _0861_ (.CLK(clknet_3_0__leaf_clk),
    .D(_0062_),
    .Q(\clk_divider_I.compare[5] ));
 sky130_fd_sc_hd__dfxtp_1 _0862_ (.CLK(clknet_3_0__leaf_clk),
    .D(_0063_),
    .Q(\clk_divider_I.compare[6] ));
 sky130_fd_sc_hd__dfxtp_1 _0863_ (.CLK(clknet_3_1__leaf_clk),
    .D(_0064_),
    .Q(\clk_divider_I.compare[7] ));
 sky130_fd_sc_hd__dfxtp_1 _0864_ (.CLK(clknet_3_4__leaf_clk),
    .D(net12),
    .Q(\aio_input_sync[0] ));
 sky130_fd_sc_hd__dfxtp_1 _0865_ (.CLK(clknet_3_3__leaf_clk),
    .D(net13),
    .Q(\aio_input_sync[1] ));
 sky130_fd_sc_hd__dfxtp_1 _0866_ (.CLK(clknet_3_6__leaf_clk),
    .D(net14),
    .Q(\aio_input_sync[2] ));
 sky130_fd_sc_hd__dfxtp_1 _0867_ (.CLK(clknet_3_7__leaf_clk),
    .D(net15),
    .Q(\aio_input_sync[3] ));
 sky130_fd_sc_hd__dfxtp_1 _0868_ (.CLK(clknet_3_3__leaf_clk),
    .D(net16),
    .Q(\aio_input_sync[4] ));
 sky130_fd_sc_hd__dfxtp_1 _0869_ (.CLK(clknet_3_3__leaf_clk),
    .D(net17),
    .Q(\aio_input_sync[5] ));
 sky130_fd_sc_hd__dfxtp_1 _0870_ (.CLK(clknet_3_2__leaf_clk),
    .D(net18),
    .Q(\aio_input_sync[6] ));
 sky130_fd_sc_hd__dfxtp_1 _0871_ (.CLK(clknet_3_6__leaf_clk),
    .D(net19),
    .Q(\aio_input_sync[7] ));
 sky130_fd_sc_hd__dfstp_1 _0872_ (.CLK(_0018_),
    .D(net42),
    .SET_B(_0017_),
    .Q(\rst_shift[0] ));
 sky130_fd_sc_hd__conb_1 _0872__42 (.LO(net42));
 sky130_fd_sc_hd__dfstp_1 _0873_ (.CLK(_0020_),
    .D(\rst_shift[0] ),
    .SET_B(_0019_),
    .Q(\rst_shift[1] ));
 sky130_fd_sc_hd__dfstp_4 _0874_ (.CLK(_0022_),
    .D(\rst_shift[1] ),
    .SET_B(_0021_),
    .Q(\clk_divider_I.reset ));
 sky130_fd_sc_hd__dfstp_2 _0875_ (.CLK(clknet_3_4__leaf_clk),
    .D(_0007_),
    .SET_B(_0023_),
    .Q(\state[0] ));
 sky130_fd_sc_hd__dfrtp_1 _0876_ (.CLK(clknet_3_7__leaf_clk),
    .D(_0008_),
    .RESET_B(_0024_),
    .Q(\state[1] ));
 sky130_fd_sc_hd__dfrtp_1 _0877_ (.CLK(clknet_3_7__leaf_clk),
    .D(_0009_),
    .RESET_B(_0025_),
    .Q(\state[2] ));
 sky130_fd_sc_hd__dfrtp_1 _0878_ (.CLK(clknet_3_6__leaf_clk),
    .D(_0010_),
    .RESET_B(_0026_),
    .Q(\state[3] ));
 sky130_fd_sc_hd__dfrtp_1 _0879_ (.CLK(clknet_3_6__leaf_clk),
    .D(_0011_),
    .RESET_B(_0027_),
    .Q(\state[4] ));
 sky130_fd_sc_hd__dfrtp_1 _0880_ (.CLK(clknet_3_7__leaf_clk),
    .D(_0012_),
    .RESET_B(_0028_),
    .Q(\state[5] ));
 sky130_fd_sc_hd__dfrtp_1 _0881_ (.CLK(clknet_3_7__leaf_clk),
    .D(_0013_),
    .RESET_B(_0029_),
    .Q(\state[6] ));
 sky130_fd_sc_hd__dfrtp_4 _0882_ (.CLK(clknet_3_4__leaf_clk),
    .D(net36),
    .RESET_B(_0030_),
    .Q(\clk_divider_I.ce ));
 sky130_fd_sc_hd__dfrtp_1 _0883_ (.CLK(clknet_3_7__leaf_clk),
    .D(_0004_),
    .RESET_B(_0031_),
    .Q(\state[9] ));
 sky130_fd_sc_hd__dfrtp_4 _0884_ (.CLK(clknet_3_6__leaf_clk),
    .D(_0005_),
    .RESET_B(_0032_),
    .Q(aio_output_cap));
 sky130_fd_sc_hd__dfrtp_4 _0885_ (.CLK(clknet_3_5__leaf_clk),
    .D(\state[4] ),
    .RESET_B(_0033_),
    .Q(aio_input_sh));
 sky130_fd_sc_hd__dfrtp_1 _0886_ (.CLK(clknet_3_7__leaf_clk),
    .D(\state[5] ),
    .RESET_B(_0034_),
    .Q(\state[12] ));
 sky130_fd_sc_hd__dfrtp_1 _0887_ (.CLK(clknet_3_7__leaf_clk),
    .D(_0006_),
    .RESET_B(_0035_),
    .Q(\state[13] ));
 sky130_fd_sc_hd__dfrtp_1 _0888_ (.CLK(clknet_3_3__leaf_clk),
    .D(_0065_),
    .RESET_B(_0036_),
    .Q(\ws_cfg[0] ));
 sky130_fd_sc_hd__dfrtp_1 _0889_ (.CLK(clknet_3_3__leaf_clk),
    .D(_0066_),
    .RESET_B(_0037_),
    .Q(\ws_cfg[1] ));
 sky130_fd_sc_hd__dfstp_1 _0890_ (.CLK(clknet_3_3__leaf_clk),
    .D(_0067_),
    .SET_B(_0038_),
    .Q(\ws_cfg[2] ));
 sky130_fd_sc_hd__dfrtp_1 _0891_ (.CLK(clknet_3_3__leaf_clk),
    .D(_0068_),
    .RESET_B(_0039_),
    .Q(\ws_cfg[3] ));
 sky130_fd_sc_hd__dfstp_1 _0892_ (.CLK(clknet_3_2__leaf_clk),
    .D(_0069_),
    .SET_B(_0040_),
    .Q(\ws_cfg[4] ));
 sky130_fd_sc_hd__dfrtp_1 _0893_ (.CLK(clknet_3_0__leaf_clk),
    .D(_0070_),
    .RESET_B(_0041_),
    .Q(\ws_cfg[5] ));
 sky130_fd_sc_hd__dfrtp_1 _0894_ (.CLK(clknet_3_0__leaf_clk),
    .D(_0071_),
    .RESET_B(_0042_),
    .Q(\ws_cfg[6] ));
 sky130_fd_sc_hd__dfrtp_1 _0895_ (.CLK(clknet_3_1__leaf_clk),
    .D(_0072_),
    .RESET_B(_0043_),
    .Q(\ws_cfg[7] ));
 sky130_fd_sc_hd__dfxtp_1 _0896_ (.CLK(clknet_3_6__leaf_clk),
    .D(_0073_),
    .Q(\aio_input_shift[1] ));
 sky130_fd_sc_hd__dfxtp_1 _0897_ (.CLK(clknet_3_6__leaf_clk),
    .D(_0074_),
    .Q(\aio_input_shift[2] ));
 sky130_fd_sc_hd__dfxtp_1 _0898_ (.CLK(clknet_3_7__leaf_clk),
    .D(_0075_),
    .Q(\aio_input_shift[3] ));
 sky130_fd_sc_hd__dfxtp_1 _0899_ (.CLK(clknet_3_3__leaf_clk),
    .D(_0076_),
    .Q(\aio_input_shift[4] ));
 sky130_fd_sc_hd__dfxtp_1 _0900_ (.CLK(clknet_3_3__leaf_clk),
    .D(_0077_),
    .Q(\aio_input_shift[5] ));
 sky130_fd_sc_hd__dfxtp_1 _0901_ (.CLK(clknet_3_6__leaf_clk),
    .D(_0078_),
    .Q(\aio_input_shift[6] ));
 sky130_fd_sc_hd__dfxtp_1 _0902_ (.CLK(clknet_3_6__leaf_clk),
    .D(_0079_),
    .Q(\aio_input_shift[7] ));
 sky130_fd_sc_hd__dfxtp_1 _0903_ (.CLK(clknet_3_5__leaf_clk),
    .D(_0080_),
    .Q(\bit_cnt[0] ));
 sky130_fd_sc_hd__dfxtp_1 _0904_ (.CLK(clknet_3_5__leaf_clk),
    .D(_0081_),
    .Q(\bit_cnt[1] ));
 sky130_fd_sc_hd__dfxtp_1 _0905_ (.CLK(clknet_3_5__leaf_clk),
    .D(_0082_),
    .Q(\bit_cnt[2] ));
 sky130_fd_sc_hd__dfxtp_1 _0906_ (.CLK(clknet_3_5__leaf_clk),
    .D(_0083_),
    .Q(\bit_cnt[3] ));
 sky130_fd_sc_hd__dfxtp_1 _0907_ (.CLK(clknet_3_5__leaf_clk),
    .D(_0084_),
    .Q(\proj_cnt[0] ));
 sky130_fd_sc_hd__dfxtp_1 _0908_ (.CLK(clknet_3_4__leaf_clk),
    .D(_0085_),
    .Q(\proj_cnt[1] ));
 sky130_fd_sc_hd__dfxtp_1 _0909_ (.CLK(clknet_3_5__leaf_clk),
    .D(_0086_),
    .Q(\proj_cnt[2] ));
 sky130_fd_sc_hd__dfxtp_1 _0910_ (.CLK(clknet_3_4__leaf_clk),
    .D(_0087_),
    .Q(\proj_cnt[3] ));
 sky130_fd_sc_hd__dfxtp_1 _0911_ (.CLK(clknet_3_4__leaf_clk),
    .D(_0088_),
    .Q(\proj_cnt[4] ));
 sky130_fd_sc_hd__dfxtp_1 _0912_ (.CLK(clknet_3_4__leaf_clk),
    .D(_0089_),
    .Q(\proj_cnt[5] ));
 sky130_fd_sc_hd__dfxtp_1 _0913_ (.CLK(clknet_3_5__leaf_clk),
    .D(_0090_),
    .Q(\proj_cnt[6] ));
 sky130_fd_sc_hd__dfxtp_1 _0914_ (.CLK(clknet_3_5__leaf_clk),
    .D(_0091_),
    .Q(\proj_cnt[7] ));
 sky130_fd_sc_hd__dfxtp_1 _0915_ (.CLK(clknet_3_5__leaf_clk),
    .D(_0092_),
    .Q(\proj_cnt[8] ));
 sky130_fd_sc_hd__dfxtp_1 _0916_ (.CLK(clknet_3_7__leaf_clk),
    .D(_0000_),
    .Q(int_scan_clk_out));
 sky130_fd_sc_hd__dfxtp_1 _0917_ (.CLK(clknet_3_3__leaf_clk),
    .D(\aio_input_shift[7] ),
    .Q(int_scan_data_out));
 sky130_fd_sc_hd__dfxtp_1 _0918_ (.CLK(clknet_3_7__leaf_clk),
    .D(_0001_),
    .Q(int_scan_select));
 sky130_fd_sc_hd__dfxtp_1 _0919_ (.CLK(clknet_3_6__leaf_clk),
    .D(\state[9] ),
    .Q(int_scan_latch_en));
 sky130_fd_sc_hd__dfxtp_1 _0920_ (.CLK(clknet_3_6__leaf_clk),
    .D(_0093_),
    .Q(\aio_input_reg[0] ));
 sky130_fd_sc_hd__dfxtp_1 _0921_ (.CLK(clknet_3_6__leaf_clk),
    .D(_0094_),
    .Q(\aio_input_reg[1] ));
 sky130_fd_sc_hd__dfxtp_1 _0922_ (.CLK(clknet_3_6__leaf_clk),
    .D(_0095_),
    .Q(\aio_input_reg[2] ));
 sky130_fd_sc_hd__dfxtp_1 _0923_ (.CLK(clknet_3_7__leaf_clk),
    .D(_0096_),
    .Q(\aio_input_reg[3] ));
 sky130_fd_sc_hd__dfxtp_1 _0924_ (.CLK(clknet_3_3__leaf_clk),
    .D(_0097_),
    .Q(\aio_input_reg[4] ));
 sky130_fd_sc_hd__dfxtp_1 _0925_ (.CLK(clknet_3_3__leaf_clk),
    .D(_0098_),
    .Q(\aio_input_reg[5] ));
 sky130_fd_sc_hd__dfxtp_1 _0926_ (.CLK(clknet_3_3__leaf_clk),
    .D(_0099_),
    .Q(\aio_input_reg[6] ));
 sky130_fd_sc_hd__dfxtp_1 _0927_ (.CLK(clknet_3_6__leaf_clk),
    .D(_0100_),
    .Q(\aio_input_reg[7] ));
 sky130_fd_sc_hd__dfxtp_1 _0928_ (.CLK(clknet_1_1__leaf_scan_clk_in),
    .D(net25),
    .Q(\aio_output_shift[0] ));
 sky130_fd_sc_hd__dfxtp_1 _0929_ (.CLK(clknet_1_1__leaf_scan_clk_in),
    .D(\aio_output_shift[0] ),
    .Q(\aio_output_shift[1] ));
 sky130_fd_sc_hd__dfxtp_1 _0930_ (.CLK(clknet_1_1__leaf_scan_clk_in),
    .D(\aio_output_shift[1] ),
    .Q(\aio_output_shift[2] ));
 sky130_fd_sc_hd__dfxtp_1 _0931_ (.CLK(clknet_1_0__leaf_scan_clk_in),
    .D(\aio_output_shift[2] ),
    .Q(\aio_output_shift[3] ));
 sky130_fd_sc_hd__dfxtp_1 _0932_ (.CLK(clknet_1_0__leaf_scan_clk_in),
    .D(\aio_output_shift[3] ),
    .Q(\aio_output_shift[4] ));
 sky130_fd_sc_hd__dfxtp_1 _0933_ (.CLK(clknet_1_0__leaf_scan_clk_in),
    .D(\aio_output_shift[4] ),
    .Q(\aio_output_shift[5] ));
 sky130_fd_sc_hd__dfxtp_1 _0934_ (.CLK(clknet_1_0__leaf_scan_clk_in),
    .D(\aio_output_shift[5] ),
    .Q(\aio_output_shift[6] ));
 sky130_fd_sc_hd__dfxtp_1 _0935_ (.CLK(clknet_1_1__leaf_scan_clk_in),
    .D(\aio_output_shift[6] ),
    .Q(\aio_output_shift[7] ));
 sky130_fd_sc_hd__dfxtp_1 _0936_ (.CLK(clknet_3_0__leaf_clk),
    .D(_0101_),
    .Q(\aio_output_reg[0] ));
 sky130_fd_sc_hd__dfxtp_1 _0937_ (.CLK(clknet_3_2__leaf_clk),
    .D(_0102_),
    .Q(\aio_output_reg[1] ));
 sky130_fd_sc_hd__dfxtp_1 _0938_ (.CLK(clknet_3_0__leaf_clk),
    .D(_0103_),
    .Q(\aio_output_reg[2] ));
 sky130_fd_sc_hd__dfxtp_1 _0939_ (.CLK(clknet_3_0__leaf_clk),
    .D(_0104_),
    .Q(\aio_output_reg[3] ));
 sky130_fd_sc_hd__dfxtp_1 _0940_ (.CLK(clknet_3_0__leaf_clk),
    .D(_0105_),
    .Q(\aio_output_reg[4] ));
 sky130_fd_sc_hd__dfxtp_1 _0941_ (.CLK(clknet_3_0__leaf_clk),
    .D(_0106_),
    .Q(\aio_output_reg[5] ));
 sky130_fd_sc_hd__dfxtp_1 _0942_ (.CLK(clknet_3_0__leaf_clk),
    .D(_0107_),
    .Q(\aio_output_reg[6] ));
 sky130_fd_sc_hd__dfxtp_1 _0943_ (.CLK(clknet_3_2__leaf_clk),
    .D(_0108_),
    .Q(\aio_output_reg[7] ));
 sky130_fd_sc_hd__dfrtp_1 _0944_ (.CLK(clknet_3_0__leaf_clk),
    .D(_0003_),
    .RESET_B(_0044_),
    .Q(\ws_set_sync[0] ));
 sky130_fd_sc_hd__dfrtp_1 _0945_ (.CLK(clknet_3_0__leaf_clk),
    .D(\ws_set_sync[0] ),
    .RESET_B(_0045_),
    .Q(\ws_set_sync[1] ));
 sky130_fd_sc_hd__dfrtp_1 _0946_ (.CLK(clknet_3_0__leaf_clk),
    .D(\ws_set_sync[1] ),
    .RESET_B(_0046_),
    .Q(\ws_set_sync[2] ));
 sky130_fd_sc_hd__dfxtp_2 _0947_ (.CLK(clknet_3_0__leaf_clk),
    .D(_0002_),
    .Q(ws_set_now));
 sky130_fd_sc_hd__dfxtp_1 _0948_ (.CLK(clknet_3_2__leaf_clk),
    .D(_0109_),
    .Q(\ws_cnt[0] ));
 sky130_fd_sc_hd__dfxtp_1 _0949_ (.CLK(clknet_3_2__leaf_clk),
    .D(_0110_),
    .Q(\ws_cnt[1] ));
 sky130_fd_sc_hd__dfxtp_1 _0950_ (.CLK(clknet_3_2__leaf_clk),
    .D(_0111_),
    .Q(\ws_cnt[2] ));
 sky130_fd_sc_hd__dfxtp_1 _0951_ (.CLK(clknet_3_2__leaf_clk),
    .D(_0112_),
    .Q(\ws_cnt[3] ));
 sky130_fd_sc_hd__dfxtp_1 _0952_ (.CLK(clknet_3_2__leaf_clk),
    .D(_0113_),
    .Q(\ws_cnt[4] ));
 sky130_fd_sc_hd__dfxtp_1 _0953_ (.CLK(clknet_3_2__leaf_clk),
    .D(_0114_),
    .Q(\ws_cnt[5] ));
 sky130_fd_sc_hd__dfxtp_1 _0954_ (.CLK(clknet_3_2__leaf_clk),
    .D(_0115_),
    .Q(\ws_cnt[6] ));
 sky130_fd_sc_hd__dfxtp_1 _0955_ (.CLK(clknet_3_2__leaf_clk),
    .D(_0116_),
    .Q(\ws_cnt[7] ));
 sky130_fd_sc_hd__dfxtp_2 _0956_ (.CLK(clknet_3_3__leaf_clk),
    .D(_0014_),
    .Q(\clk_divider_I.set_now ));
 sky130_fd_sc_hd__dfxtp_1 _0957_ (.CLK(clknet_3_3__leaf_clk),
    .D(net26),
    .Q(\clk_divider_I.set_sync[0] ));
 sky130_fd_sc_hd__dfxtp_1 _0958_ (.CLK(clknet_3_3__leaf_clk),
    .D(\clk_divider_I.set_sync[0] ),
    .Q(\clk_divider_I.set_sync[1] ));
 sky130_fd_sc_hd__dfxtp_1 _0959_ (.CLK(clknet_3_3__leaf_clk),
    .D(\clk_divider_I.set_sync[1] ),
    .Q(\clk_divider_I.active ));
 sky130_fd_sc_hd__dfrtp_1 _0960_ (.CLK(clknet_3_4__leaf_clk),
    .D(_0117_),
    .RESET_B(_0047_),
    .Q(\clk_divider_I.counter[0] ));
 sky130_fd_sc_hd__dfrtp_1 _0961_ (.CLK(clknet_3_4__leaf_clk),
    .D(_0118_),
    .RESET_B(_0048_),
    .Q(\clk_divider_I.counter[1] ));
 sky130_fd_sc_hd__dfrtp_1 _0962_ (.CLK(clknet_3_4__leaf_clk),
    .D(_0119_),
    .RESET_B(_0049_),
    .Q(\clk_divider_I.counter[2] ));
 sky130_fd_sc_hd__dfrtp_1 _0963_ (.CLK(clknet_3_4__leaf_clk),
    .D(_0120_),
    .RESET_B(_0050_),
    .Q(\clk_divider_I.counter[3] ));
 sky130_fd_sc_hd__dfrtp_1 _0964_ (.CLK(clknet_3_1__leaf_clk),
    .D(_0121_),
    .RESET_B(_0051_),
    .Q(\clk_divider_I.counter[4] ));
 sky130_fd_sc_hd__dfrtp_1 _0965_ (.CLK(clknet_3_1__leaf_clk),
    .D(_0122_),
    .RESET_B(_0052_),
    .Q(\clk_divider_I.counter[5] ));
 sky130_fd_sc_hd__dfrtp_1 _0966_ (.CLK(clknet_3_1__leaf_clk),
    .D(_0123_),
    .RESET_B(_0053_),
    .Q(\clk_divider_I.counter[6] ));
 sky130_fd_sc_hd__dfrtp_1 _0967_ (.CLK(clknet_3_1__leaf_clk),
    .D(_0124_),
    .RESET_B(_0054_),
    .Q(\clk_divider_I.counter[7] ));
 sky130_fd_sc_hd__dfrtp_4 _0968_ (.CLK(clknet_3_4__leaf_clk),
    .D(_0125_),
    .RESET_B(_0055_),
    .Q(net41));
 sky130_fd_sc_hd__dfxtp_1 _0969_ (.CLK(clknet_3_6__leaf_clk),
    .D(_0126_),
    .Q(\aio_input_shift[0] ));
 sky130_fd_sc_hd__clkbuf_1 _1009_ (.A(net25),
    .X(net27));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_scan_clk_in (.A(scan_clk_in),
    .X(clknet_0_scan_clk_in));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_scan_clk_in (.A(clknet_0_scan_clk_in),
    .X(clknet_1_0__leaf_scan_clk_in));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_scan_clk_in (.A(clknet_0_scan_clk_in),
    .X(clknet_1_1__leaf_scan_clk_in));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_0__f_clk (.A(clknet_0_clk),
    .X(clknet_3_0__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_1__f_clk (.A(clknet_0_clk),
    .X(clknet_3_1__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_2__f_clk (.A(clknet_0_clk),
    .X(clknet_3_2__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_3__f_clk (.A(clknet_0_clk),
    .X(clknet_3_3__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_4__f_clk (.A(clknet_0_clk),
    .X(clknet_3_4__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_5__f_clk (.A(clknet_0_clk),
    .X(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_6__f_clk (.A(clknet_0_clk),
    .X(clknet_3_6__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_7__f_clk (.A(clknet_0_clk),
    .X(clknet_3_7__leaf_clk));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1 (.A(\aio_output_shift[7] ),
    .X(net84));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2 (.A(\aio_output_shift[5] ),
    .X(net85));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3 (.A(\aio_output_shift[3] ),
    .X(net86));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4 (.A(\aio_output_shift[0] ),
    .X(net87));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5 (.A(\aio_output_shift[6] ),
    .X(net88));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6 (.A(\aio_output_shift[4] ),
    .X(net89));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7 (.A(\aio_output_shift[1] ),
    .X(net90));
 sky130_fd_sc_hd__dlygate4sd3_1 hold8 (.A(\aio_output_shift[2] ),
    .X(net91));
 sky130_fd_sc_hd__buf_2 input1 (.A(active_select[0]),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_4 input10 (.A(driver_sel[0]),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_2 input11 (.A(driver_sel[1]),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_2 input12 (.A(inputs[0]),
    .X(net12));
 sky130_fd_sc_hd__dlymetal6s2s_1 input13 (.A(inputs[1]),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_2 input14 (.A(inputs[2]),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_2 input15 (.A(inputs[3]),
    .X(net15));
 sky130_fd_sc_hd__dlymetal6s2s_1 input16 (.A(inputs[4]),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_1 input17 (.A(inputs[5]),
    .X(net17));
 sky130_fd_sc_hd__dlymetal6s2s_1 input18 (.A(inputs[6]),
    .X(net18));
 sky130_fd_sc_hd__clkbuf_2 input19 (.A(inputs[7]),
    .X(net19));
 sky130_fd_sc_hd__clkbuf_1 input2 (.A(active_select[1]),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_1 input20 (.A(la_scan_clk_in),
    .X(net20));
 sky130_fd_sc_hd__clkbuf_1 input21 (.A(la_scan_data_in),
    .X(net21));
 sky130_fd_sc_hd__clkbuf_1 input22 (.A(la_scan_latch_en),
    .X(net22));
 sky130_fd_sc_hd__clkbuf_1 input23 (.A(la_scan_select),
    .X(net23));
 sky130_fd_sc_hd__dlymetal6s2s_1 input24 (.A(reset),
    .X(net24));
 sky130_fd_sc_hd__clkbuf_2 input25 (.A(scan_data_in),
    .X(net25));
 sky130_fd_sc_hd__clkbuf_1 input26 (.A(set_clk_div),
    .X(net26));
 sky130_fd_sc_hd__clkbuf_1 input3 (.A(active_select[2]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_1 input4 (.A(active_select[3]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_1 input5 (.A(active_select[4]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_1 input6 (.A(active_select[5]),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_1 input7 (.A(active_select[6]),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_2 input8 (.A(active_select[7]),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_2 input9 (.A(active_select[8]),
    .X(net9));
 sky130_fd_sc_hd__buf_12 output27 (.A(net27),
    .X(la_scan_data_out));
 sky130_fd_sc_hd__clkbuf_1 output28 (.A(net28),
    .X(outputs[0]));
 sky130_fd_sc_hd__buf_12 output29 (.A(net29),
    .X(outputs[1]));
 sky130_fd_sc_hd__buf_12 output30 (.A(net30),
    .X(outputs[2]));
 sky130_fd_sc_hd__buf_12 output31 (.A(net31),
    .X(outputs[3]));
 sky130_fd_sc_hd__buf_12 output32 (.A(net32),
    .X(outputs[4]));
 sky130_fd_sc_hd__buf_12 output33 (.A(net33),
    .X(outputs[5]));
 sky130_fd_sc_hd__buf_12 output34 (.A(net34),
    .X(outputs[6]));
 sky130_fd_sc_hd__buf_12 output35 (.A(net35),
    .X(outputs[7]));
 sky130_fd_sc_hd__buf_12 output36 (.A(net36),
    .X(ready));
 sky130_fd_sc_hd__buf_12 output37 (.A(net37),
    .X(scan_clk_out));
 sky130_fd_sc_hd__buf_12 output38 (.A(net38),
    .X(scan_data_out));
 sky130_fd_sc_hd__buf_12 output39 (.A(net39),
    .X(scan_latch_en));
 sky130_fd_sc_hd__buf_12 output40 (.A(net40),
    .X(scan_select));
 sky130_fd_sc_hd__buf_12 output41 (.A(net41),
    .X(slow_clk));
 sky130_fd_sc_hd__conb_1 scan_controller_43 (.LO(net43));
 sky130_fd_sc_hd__conb_1 scan_controller_44 (.LO(net44));
 sky130_fd_sc_hd__conb_1 scan_controller_45 (.LO(net45));
 sky130_fd_sc_hd__conb_1 scan_controller_46 (.LO(net46));
 sky130_fd_sc_hd__conb_1 scan_controller_47 (.LO(net47));
 sky130_fd_sc_hd__conb_1 scan_controller_48 (.LO(net48));
 sky130_fd_sc_hd__conb_1 scan_controller_49 (.LO(net49));
 sky130_fd_sc_hd__conb_1 scan_controller_50 (.LO(net50));
 sky130_fd_sc_hd__conb_1 scan_controller_51 (.LO(net51));
 sky130_fd_sc_hd__conb_1 scan_controller_52 (.LO(net52));
 sky130_fd_sc_hd__conb_1 scan_controller_53 (.LO(net53));
 sky130_fd_sc_hd__conb_1 scan_controller_54 (.LO(net54));
 sky130_fd_sc_hd__conb_1 scan_controller_55 (.LO(net55));
 sky130_fd_sc_hd__conb_1 scan_controller_56 (.LO(net56));
 sky130_fd_sc_hd__conb_1 scan_controller_57 (.LO(net57));
 sky130_fd_sc_hd__conb_1 scan_controller_58 (.LO(net58));
 sky130_fd_sc_hd__conb_1 scan_controller_59 (.LO(net59));
 sky130_fd_sc_hd__conb_1 scan_controller_60 (.LO(net60));
 sky130_fd_sc_hd__conb_1 scan_controller_61 (.LO(net61));
 sky130_fd_sc_hd__conb_1 scan_controller_62 (.LO(net62));
 sky130_fd_sc_hd__conb_1 scan_controller_63 (.LO(net63));
 sky130_fd_sc_hd__conb_1 scan_controller_64 (.LO(net64));
 sky130_fd_sc_hd__conb_1 scan_controller_65 (.LO(net65));
 sky130_fd_sc_hd__conb_1 scan_controller_66 (.LO(net66));
 sky130_fd_sc_hd__conb_1 scan_controller_67 (.LO(net67));
 sky130_fd_sc_hd__conb_1 scan_controller_68 (.LO(net68));
 sky130_fd_sc_hd__conb_1 scan_controller_69 (.LO(net69));
 sky130_fd_sc_hd__conb_1 scan_controller_70 (.LO(net70));
 sky130_fd_sc_hd__conb_1 scan_controller_71 (.LO(net71));
 sky130_fd_sc_hd__conb_1 scan_controller_72 (.LO(net72));
 sky130_fd_sc_hd__conb_1 scan_controller_73 (.LO(net73));
 sky130_fd_sc_hd__conb_1 scan_controller_74 (.LO(net74));
 sky130_fd_sc_hd__conb_1 scan_controller_75 (.LO(net75));
 sky130_fd_sc_hd__conb_1 scan_controller_76 (.LO(net76));
 sky130_fd_sc_hd__conb_1 scan_controller_77 (.LO(net77));
 sky130_fd_sc_hd__conb_1 scan_controller_78 (.LO(net78));
 sky130_fd_sc_hd__conb_1 scan_controller_79 (.LO(net79));
 sky130_fd_sc_hd__conb_1 scan_controller_80 (.LO(net80));
 assign oeb[0] = net43;
 assign oeb[10] = net53;
 assign oeb[11] = net54;
 assign oeb[12] = net55;
 assign oeb[13] = net56;
 assign oeb[14] = net57;
 assign oeb[15] = net58;
 assign oeb[16] = net59;
 assign oeb[17] = net60;
 assign oeb[18] = net61;
 assign oeb[19] = net62;
 assign oeb[1] = net44;
 assign oeb[20] = net63;
 assign oeb[21] = net64;
 assign oeb[22] = net65;
 assign oeb[23] = net66;
 assign oeb[24] = net67;
 assign oeb[25] = net68;
 assign oeb[26] = net69;
 assign oeb[27] = net70;
 assign oeb[28] = net71;
 assign oeb[29] = net72;
 assign oeb[2] = net45;
 assign oeb[30] = net73;
 assign oeb[31] = net74;
 assign oeb[32] = net75;
 assign oeb[33] = net76;
 assign oeb[34] = net77;
 assign oeb[35] = net78;
 assign oeb[36] = net79;
 assign oeb[37] = net80;
 assign oeb[3] = net46;
 assign oeb[4] = net47;
 assign oeb[5] = net48;
 assign oeb[6] = net49;
 assign oeb[7] = net50;
 assign oeb[8] = net51;
 assign oeb[9] = net52;
endmodule

