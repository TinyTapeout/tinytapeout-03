magic
tech sky130A
magscale 1 2
timestamp 1682078255
<< viali >>
rect 17693 17289 17727 17323
rect 20913 17289 20947 17323
rect 40877 17289 40911 17323
rect 44281 17289 44315 17323
rect 1685 17221 1719 17255
rect 3249 17221 3283 17255
rect 4721 17221 4755 17255
rect 11805 17221 11839 17255
rect 16129 17221 16163 17255
rect 32413 17221 32447 17255
rect 38853 17221 38887 17255
rect 2421 17153 2455 17187
rect 6745 17153 6779 17187
rect 8033 17153 8067 17187
rect 9965 17153 9999 17187
rect 13185 17153 13219 17187
rect 14473 17153 14507 17187
rect 17509 17153 17543 17187
rect 19625 17153 19659 17187
rect 20729 17153 20763 17187
rect 22845 17153 22879 17187
rect 24777 17153 24811 17187
rect 26065 17153 26099 17187
rect 27997 17153 28031 17187
rect 29929 17153 29963 17187
rect 31217 17153 31251 17187
rect 35081 17153 35115 17187
rect 35725 17153 35759 17187
rect 37657 17153 37691 17187
rect 40693 17153 40727 17187
rect 42809 17153 42843 17187
rect 43637 17153 43671 17187
rect 44097 17153 44131 17187
rect 1869 17017 1903 17051
rect 3433 17017 3467 17051
rect 11989 17017 12023 17051
rect 16313 17017 16347 17051
rect 2513 16949 2547 16983
rect 4813 16949 4847 16983
rect 9781 16949 9815 16983
rect 24593 16949 24627 16983
rect 31033 16949 31067 16983
rect 32505 16949 32539 16983
rect 34897 16949 34931 16983
rect 38945 16949 38979 16983
rect 43729 16745 43763 16779
rect 44373 16745 44407 16779
rect 1869 16609 1903 16643
rect 1685 16541 1719 16575
rect 14565 16541 14599 16575
rect 28549 16541 28583 16575
rect 14381 16405 14415 16439
rect 28365 16405 28399 16439
rect 42993 16201 43027 16235
rect 1777 16065 1811 16099
rect 42809 16065 42843 16099
rect 43269 16065 43303 16099
rect 44373 15861 44407 15895
rect 32321 15657 32355 15691
rect 1593 15453 1627 15487
rect 32137 15385 32171 15419
rect 1777 15317 1811 15351
rect 32337 15317 32371 15351
rect 32505 15317 32539 15351
rect 23305 15113 23339 15147
rect 26341 15113 26375 15147
rect 26249 15045 26283 15079
rect 32597 15045 32631 15079
rect 23213 14977 23247 15011
rect 31493 14977 31527 15011
rect 33609 14977 33643 15011
rect 33885 14977 33919 15011
rect 34345 14977 34379 15011
rect 34529 14977 34563 15011
rect 36369 14977 36403 15011
rect 36553 14977 36587 15011
rect 37657 14977 37691 15011
rect 18153 14909 18187 14943
rect 18429 14909 18463 14943
rect 23397 14909 23431 14943
rect 26525 14909 26559 14943
rect 31769 14909 31803 14943
rect 32321 14909 32355 14943
rect 32689 14909 32723 14943
rect 32806 14909 32840 14943
rect 33793 14909 33827 14943
rect 31585 14841 31619 14875
rect 19901 14773 19935 14807
rect 22845 14773 22879 14807
rect 25881 14773 25915 14807
rect 31493 14773 31527 14807
rect 32965 14773 32999 14807
rect 33425 14773 33459 14807
rect 34713 14773 34747 14807
rect 36461 14773 36495 14807
rect 37473 14773 37507 14807
rect 33241 14569 33275 14603
rect 34897 14569 34931 14603
rect 41337 14569 41371 14603
rect 18797 14501 18831 14535
rect 42809 14501 42843 14535
rect 22753 14433 22787 14467
rect 9873 14365 9907 14399
rect 10129 14365 10163 14399
rect 18245 14365 18279 14399
rect 18705 14365 18739 14399
rect 19441 14365 19475 14399
rect 20361 14365 20395 14399
rect 26157 14365 26191 14399
rect 31309 14365 31343 14399
rect 31565 14365 31599 14399
rect 33425 14365 33459 14399
rect 33609 14365 33643 14399
rect 34897 14365 34931 14399
rect 35081 14365 35115 14399
rect 36829 14365 36863 14399
rect 37096 14365 37130 14399
rect 40969 14365 41003 14399
rect 42165 14365 42199 14399
rect 42993 14365 43027 14399
rect 44097 14365 44131 14399
rect 20606 14297 20640 14331
rect 22661 14297 22695 14331
rect 26424 14297 26458 14331
rect 33149 14297 33183 14331
rect 36001 14297 36035 14331
rect 36185 14297 36219 14331
rect 11253 14229 11287 14263
rect 18061 14229 18095 14263
rect 19533 14229 19567 14263
rect 21741 14229 21775 14263
rect 22201 14229 22235 14263
rect 22569 14229 22603 14263
rect 27537 14229 27571 14263
rect 32689 14229 32723 14263
rect 33793 14229 33827 14263
rect 36369 14229 36403 14263
rect 38209 14229 38243 14263
rect 41337 14229 41371 14263
rect 41521 14229 41555 14263
rect 41981 14229 42015 14263
rect 44281 14229 44315 14263
rect 6643 14025 6677 14059
rect 17325 14025 17359 14059
rect 20085 14025 20119 14059
rect 21373 14025 21407 14059
rect 22293 14025 22327 14059
rect 24317 14025 24351 14059
rect 25145 14025 25179 14059
rect 27629 14025 27663 14059
rect 31591 14025 31625 14059
rect 34253 14025 34287 14059
rect 36553 14025 36587 14059
rect 36645 14025 36679 14059
rect 36921 14025 36955 14059
rect 7113 13957 7147 13991
rect 20453 13957 20487 13991
rect 23182 13957 23216 13991
rect 25237 13957 25271 13991
rect 26065 13957 26099 13991
rect 30205 13957 30239 13991
rect 31493 13957 31527 13991
rect 36762 13957 36796 13991
rect 37657 13957 37691 13991
rect 40960 13957 40994 13991
rect 5365 13889 5399 13923
rect 6929 13889 6963 13923
rect 12633 13889 12667 13923
rect 13360 13889 13394 13923
rect 17233 13889 17267 13923
rect 17877 13889 17911 13923
rect 20269 13889 20303 13923
rect 20545 13889 20579 13923
rect 21189 13889 21223 13923
rect 22477 13889 22511 13923
rect 22937 13889 22971 13923
rect 26249 13889 26283 13923
rect 27537 13889 27571 13923
rect 28365 13889 28399 13923
rect 28632 13889 28666 13923
rect 30481 13889 30515 13923
rect 30573 13889 30607 13923
rect 30665 13889 30699 13923
rect 30849 13889 30883 13923
rect 31677 13889 31711 13923
rect 31769 13889 31803 13923
rect 32873 13889 32907 13923
rect 33140 13889 33174 13923
rect 34805 13889 34839 13923
rect 34989 13889 35023 13923
rect 35449 13889 35483 13923
rect 35541 13889 35575 13923
rect 37473 13889 37507 13923
rect 37749 13889 37783 13923
rect 38209 13889 38243 13923
rect 38393 13889 38427 13923
rect 1777 13821 1811 13855
rect 5181 13821 5215 13855
rect 7205 13821 7239 13855
rect 13093 13821 13127 13855
rect 18153 13821 18187 13855
rect 21005 13821 21039 13855
rect 25329 13821 25363 13855
rect 27721 13821 27755 13855
rect 34897 13821 34931 13855
rect 36277 13821 36311 13855
rect 38301 13821 38335 13855
rect 40693 13821 40727 13855
rect 27169 13753 27203 13787
rect 5549 13685 5583 13719
rect 12449 13685 12483 13719
rect 14473 13685 14507 13719
rect 19625 13685 19659 13719
rect 24777 13685 24811 13719
rect 26433 13685 26467 13719
rect 29745 13685 29779 13719
rect 37473 13685 37507 13719
rect 42073 13685 42107 13719
rect 14657 13481 14691 13515
rect 19625 13481 19659 13515
rect 20545 13481 20579 13515
rect 21557 13481 21591 13515
rect 26341 13481 26375 13515
rect 26801 13481 26835 13515
rect 29745 13481 29779 13515
rect 32137 13481 32171 13515
rect 35541 13481 35575 13515
rect 42809 13481 42843 13515
rect 6929 13413 6963 13447
rect 18889 13413 18923 13447
rect 28825 13413 28859 13447
rect 31861 13413 31895 13447
rect 40233 13413 40267 13447
rect 7573 13345 7607 13379
rect 10885 13345 10919 13379
rect 11437 13345 11471 13379
rect 17141 13345 17175 13379
rect 20729 13345 20763 13379
rect 22201 13345 22235 13379
rect 30941 13345 30975 13379
rect 36093 13345 36127 13379
rect 36921 13345 36955 13379
rect 4629 13277 4663 13311
rect 5089 13277 5123 13311
rect 11693 13277 11727 13311
rect 14381 13277 14415 13311
rect 14473 13277 14507 13311
rect 19809 13277 19843 13311
rect 19993 13277 20027 13311
rect 20085 13277 20119 13311
rect 20821 13277 20855 13311
rect 21465 13277 21499 13311
rect 22385 13277 22419 13311
rect 22569 13277 22603 13311
rect 23765 13277 23799 13311
rect 24593 13277 24627 13311
rect 26985 13277 27019 13311
rect 28733 13277 28767 13311
rect 28917 13277 28951 13311
rect 29929 13277 29963 13311
rect 30021 13277 30055 13311
rect 31033 13277 31067 13311
rect 32316 13277 32350 13311
rect 32688 13277 32722 13311
rect 32781 13277 32815 13311
rect 33241 13277 33275 13311
rect 33425 13277 33459 13311
rect 35449 13277 35483 13311
rect 36277 13277 36311 13311
rect 37188 13277 37222 13311
rect 40509 13277 40543 13311
rect 40969 13277 41003 13311
rect 41225 13277 41259 13311
rect 42993 13277 43027 13311
rect 43269 13277 43303 13311
rect 5334 13209 5368 13243
rect 7297 13209 7331 13243
rect 10609 13209 10643 13243
rect 17417 13209 17451 13243
rect 20545 13209 20579 13243
rect 24869 13209 24903 13243
rect 29745 13209 29779 13243
rect 32413 13209 32447 13243
rect 32505 13209 32539 13243
rect 40233 13209 40267 13243
rect 43177 13209 43211 13243
rect 4445 13141 4479 13175
rect 6469 13141 6503 13175
rect 7389 13141 7423 13175
rect 10241 13141 10275 13175
rect 10701 13141 10735 13175
rect 12817 13141 12851 13175
rect 21005 13141 21039 13175
rect 23581 13141 23615 13175
rect 31401 13141 31435 13175
rect 33333 13141 33367 13175
rect 36461 13141 36495 13175
rect 38301 13141 38335 13175
rect 40417 13141 40451 13175
rect 42349 13141 42383 13175
rect 5457 12937 5491 12971
rect 11713 12937 11747 12971
rect 12173 12937 12207 12971
rect 14565 12937 14599 12971
rect 15025 12937 15059 12971
rect 20269 12937 20303 12971
rect 22385 12937 22419 12971
rect 27353 12937 27387 12971
rect 31401 12937 31435 12971
rect 33625 12937 33659 12971
rect 33793 12937 33827 12971
rect 37473 12937 37507 12971
rect 38393 12937 38427 12971
rect 40233 12937 40267 12971
rect 40417 12937 40451 12971
rect 41245 12937 41279 12971
rect 41613 12937 41647 12971
rect 13452 12869 13486 12903
rect 17969 12869 18003 12903
rect 31493 12869 31527 12903
rect 32321 12869 32355 12903
rect 33425 12869 33459 12903
rect 34437 12869 34471 12903
rect 40141 12869 40175 12903
rect 3157 12801 3191 12835
rect 4077 12801 4111 12835
rect 4344 12801 4378 12835
rect 6828 12801 6862 12835
rect 8585 12801 8619 12835
rect 9781 12801 9815 12835
rect 10048 12801 10082 12835
rect 12081 12801 12115 12835
rect 15209 12801 15243 12835
rect 17877 12801 17911 12835
rect 18521 12801 18555 12835
rect 20913 12801 20947 12835
rect 21005 12801 21039 12835
rect 21097 12801 21131 12835
rect 21235 12801 21269 12835
rect 22017 12801 22051 12835
rect 24869 12801 24903 12835
rect 25881 12801 25915 12835
rect 26065 12801 26099 12835
rect 26249 12801 26283 12835
rect 27261 12801 27295 12835
rect 29193 12801 29227 12835
rect 29460 12801 29494 12835
rect 31585 12801 31619 12835
rect 31769 12801 31803 12835
rect 32689 12801 32723 12835
rect 32781 12801 32815 12835
rect 35449 12801 35483 12835
rect 35633 12801 35667 12835
rect 36093 12801 36127 12835
rect 36277 12801 36311 12835
rect 36461 12801 36495 12835
rect 36645 12801 36679 12835
rect 37657 12801 37691 12835
rect 37841 12801 37875 12835
rect 37933 12801 37967 12835
rect 38577 12801 38611 12835
rect 38761 12801 38795 12835
rect 38853 12801 38887 12835
rect 39313 12801 39347 12835
rect 39497 12801 39531 12835
rect 40049 12801 40083 12835
rect 41521 12801 41555 12835
rect 6561 12733 6595 12767
rect 12357 12733 12391 12767
rect 13185 12733 13219 12767
rect 18797 12733 18831 12767
rect 20729 12733 20763 12767
rect 21373 12733 21407 12767
rect 22109 12733 22143 12767
rect 24961 12733 24995 12767
rect 35541 12733 35575 12767
rect 36369 12733 36403 12767
rect 39405 12733 39439 12767
rect 40417 12733 40451 12767
rect 41429 12733 41463 12767
rect 41797 12733 41831 12767
rect 41889 12733 41923 12767
rect 8401 12665 8435 12699
rect 31217 12665 31251 12699
rect 34621 12665 34655 12699
rect 2973 12597 3007 12631
rect 7941 12597 7975 12631
rect 11161 12597 11195 12631
rect 22201 12597 22235 12631
rect 30573 12597 30607 12631
rect 32965 12597 32999 12631
rect 33609 12597 33643 12631
rect 36829 12597 36863 12631
rect 44373 12597 44407 12631
rect 2973 12393 3007 12427
rect 7389 12393 7423 12427
rect 10149 12393 10183 12427
rect 12173 12393 12207 12427
rect 13001 12393 13035 12427
rect 21189 12393 21223 12427
rect 26893 12393 26927 12427
rect 32965 12393 32999 12427
rect 35449 12393 35483 12427
rect 36461 12393 36495 12427
rect 36921 12393 36955 12427
rect 31033 12325 31067 12359
rect 4905 12257 4939 12291
rect 8033 12257 8067 12291
rect 13645 12257 13679 12291
rect 15209 12257 15243 12291
rect 19441 12257 19475 12291
rect 19717 12257 19751 12291
rect 21649 12257 21683 12291
rect 22293 12257 22327 12291
rect 24593 12257 24627 12291
rect 30021 12257 30055 12291
rect 36093 12257 36127 12291
rect 40509 12257 40543 12291
rect 40718 12257 40752 12291
rect 3157 12189 3191 12223
rect 5457 12189 5491 12223
rect 7757 12189 7791 12223
rect 10333 12189 10367 12223
rect 10793 12189 10827 12223
rect 15025 12189 15059 12223
rect 18705 12189 18739 12223
rect 21833 12189 21867 12223
rect 22017 12189 22051 12223
rect 22753 12189 22787 12223
rect 23029 12189 23063 12223
rect 23121 12189 23155 12223
rect 26801 12189 26835 12223
rect 29745 12189 29779 12223
rect 31309 12189 31343 12223
rect 31769 12189 31803 12223
rect 31953 12189 31987 12223
rect 32045 12189 32079 12223
rect 32321 12189 32355 12223
rect 34069 12189 34103 12223
rect 36277 12189 36311 12223
rect 37197 12189 37231 12223
rect 37289 12189 37323 12223
rect 37381 12189 37415 12223
rect 37565 12189 37599 12223
rect 38025 12189 38059 12223
rect 38209 12189 38243 12223
rect 38853 12189 38887 12223
rect 38945 12189 38979 12223
rect 39129 12189 39163 12223
rect 39221 12189 39255 12223
rect 39313 12189 39347 12223
rect 40233 12189 40267 12223
rect 41797 12189 41831 12223
rect 42073 12189 42107 12223
rect 42257 12189 42291 12223
rect 5724 12121 5758 12155
rect 11060 12121 11094 12155
rect 21925 12121 21959 12155
rect 22135 12121 22169 12155
rect 22937 12121 22971 12155
rect 24869 12121 24903 12155
rect 31033 12121 31067 12155
rect 32137 12121 32171 12155
rect 32781 12121 32815 12155
rect 32997 12121 33031 12155
rect 35265 12121 35299 12155
rect 35481 12121 35515 12155
rect 40601 12121 40635 12155
rect 4261 12053 4295 12087
rect 4629 12053 4663 12087
rect 4721 12053 4755 12087
rect 6837 12053 6871 12087
rect 7849 12053 7883 12087
rect 13369 12053 13403 12087
rect 13461 12053 13495 12087
rect 14657 12053 14691 12087
rect 15117 12053 15151 12087
rect 18797 12053 18831 12087
rect 23305 12053 23339 12087
rect 26341 12053 26375 12087
rect 31217 12053 31251 12087
rect 33149 12053 33183 12087
rect 34253 12053 34287 12087
rect 35633 12053 35667 12087
rect 38393 12053 38427 12087
rect 38853 12053 38887 12087
rect 40877 12053 40911 12087
rect 41613 12053 41647 12087
rect 3985 11849 4019 11883
rect 6009 11849 6043 11883
rect 7389 11849 7423 11883
rect 7481 11849 7515 11883
rect 8217 11849 8251 11883
rect 14565 11849 14599 11883
rect 15025 11849 15059 11883
rect 19717 11849 19751 11883
rect 20085 11849 20119 11883
rect 22937 11849 22971 11883
rect 26617 11849 26651 11883
rect 29377 11849 29411 11883
rect 32689 11849 32723 11883
rect 33517 11849 33551 11883
rect 37841 11849 37875 11883
rect 38117 11849 38151 11883
rect 38577 11849 38611 11883
rect 38945 11849 38979 11883
rect 41429 11849 41463 11883
rect 8677 11781 8711 11815
rect 13452 11781 13486 11815
rect 20177 11781 20211 11815
rect 25145 11781 25179 11815
rect 28825 11781 28859 11815
rect 33149 11781 33183 11815
rect 33365 11781 33399 11815
rect 36461 11781 36495 11815
rect 37749 11781 37783 11815
rect 37958 11781 37992 11815
rect 41797 11781 41831 11815
rect 3433 11713 3467 11747
rect 4169 11713 4203 11747
rect 4896 11713 4930 11747
rect 8585 11713 8619 11747
rect 10333 11713 10367 11747
rect 13185 11713 13219 11747
rect 15209 11713 15243 11747
rect 17233 11713 17267 11747
rect 19257 11713 19291 11747
rect 21373 11713 21407 11747
rect 21465 11713 21499 11747
rect 22109 11713 22143 11747
rect 22201 11713 22235 11747
rect 22845 11713 22879 11747
rect 23029 11713 23063 11747
rect 28641 11713 28675 11747
rect 28917 11713 28951 11747
rect 29561 11713 29595 11747
rect 30564 11713 30598 11747
rect 32505 11713 32539 11747
rect 34244 11713 34278 11747
rect 35817 11713 35851 11747
rect 36645 11713 36679 11747
rect 38853 11713 38887 11747
rect 39037 11713 39071 11747
rect 40785 11713 40819 11747
rect 41613 11713 41647 11747
rect 41889 11713 41923 11747
rect 4629 11645 4663 11679
rect 7665 11645 7699 11679
rect 8861 11645 8895 11679
rect 17325 11645 17359 11679
rect 17509 11645 17543 11679
rect 20269 11645 20303 11679
rect 21189 11645 21223 11679
rect 24869 11645 24903 11679
rect 29745 11645 29779 11679
rect 29837 11645 29871 11679
rect 30297 11645 30331 11679
rect 32321 11645 32355 11679
rect 33977 11645 34011 11679
rect 36829 11645 36863 11679
rect 37473 11645 37507 11679
rect 39221 11645 39255 11679
rect 39313 11645 39347 11679
rect 35357 11577 35391 11611
rect 40877 11577 40911 11611
rect 3249 11509 3283 11543
rect 7021 11509 7055 11543
rect 10149 11509 10183 11543
rect 16865 11509 16899 11543
rect 19073 11509 19107 11543
rect 21005 11509 21039 11543
rect 22385 11509 22419 11543
rect 28641 11509 28675 11543
rect 31677 11509 31711 11543
rect 33333 11509 33367 11543
rect 35909 11509 35943 11543
rect 36737 11509 36771 11543
rect 36921 11509 36955 11543
rect 3433 11305 3467 11339
rect 5549 11305 5583 11339
rect 6009 11305 6043 11339
rect 14657 11305 14691 11339
rect 17141 11305 17175 11339
rect 21189 11305 21223 11339
rect 25513 11305 25547 11339
rect 26157 11305 26191 11339
rect 32597 11305 32631 11339
rect 35173 11305 35207 11339
rect 35265 11305 35299 11339
rect 39221 11305 39255 11339
rect 6745 11237 6779 11271
rect 13737 11237 13771 11271
rect 32689 11237 32723 11271
rect 37381 11237 37415 11271
rect 7205 11169 7239 11203
rect 7389 11169 7423 11203
rect 9965 11169 9999 11203
rect 12357 11169 12391 11203
rect 19717 11169 19751 11203
rect 24777 11169 24811 11203
rect 41429 11169 41463 11203
rect 3157 11101 3191 11135
rect 3249 11101 3283 11135
rect 4169 11101 4203 11135
rect 4425 11101 4459 11135
rect 6193 11101 6227 11135
rect 7941 11101 7975 11135
rect 10232 11101 10266 11135
rect 12624 11101 12658 11135
rect 14381 11101 14415 11135
rect 14473 11101 14507 11135
rect 15761 11101 15795 11135
rect 19441 11101 19475 11135
rect 22661 11101 22695 11135
rect 24593 11101 24627 11135
rect 24685 11101 24719 11135
rect 24961 11101 24995 11135
rect 25421 11101 25455 11135
rect 26065 11101 26099 11135
rect 30297 11101 30331 11135
rect 30665 11101 30699 11135
rect 32091 11101 32125 11135
rect 32597 11101 32631 11135
rect 32873 11101 32907 11135
rect 35081 11101 35115 11135
rect 35265 11101 35299 11135
rect 36553 11101 36587 11135
rect 36829 11101 36863 11135
rect 37289 11101 37323 11135
rect 37565 11101 37599 11135
rect 38025 11101 38059 11135
rect 38209 11101 38243 11135
rect 38301 11101 38335 11135
rect 38393 11101 38427 11135
rect 38577 11101 38611 11135
rect 39221 11101 39255 11135
rect 39405 11101 39439 11135
rect 39497 11101 39531 11135
rect 41696 11101 41730 11135
rect 44373 11101 44407 11135
rect 7113 11033 7147 11067
rect 16006 11033 16040 11067
rect 34897 11033 34931 11067
rect 36737 11033 36771 11067
rect 37473 11033 37507 11067
rect 38761 11033 38795 11067
rect 8585 10965 8619 10999
rect 11345 10965 11379 10999
rect 22477 10965 22511 10999
rect 24869 10965 24903 10999
rect 36369 10965 36403 10999
rect 42809 10965 42843 10999
rect 2329 10761 2363 10795
rect 5365 10761 5399 10795
rect 8309 10761 8343 10795
rect 9597 10761 9631 10795
rect 10333 10761 10367 10795
rect 10793 10761 10827 10795
rect 13093 10761 13127 10795
rect 14013 10761 14047 10795
rect 15485 10761 15519 10795
rect 16129 10761 16163 10795
rect 16957 10761 16991 10795
rect 17325 10761 17359 10795
rect 20821 10761 20855 10795
rect 26157 10761 26191 10795
rect 27353 10761 27387 10795
rect 30849 10761 30883 10795
rect 31217 10761 31251 10795
rect 32413 10761 32447 10795
rect 36369 10761 36403 10795
rect 38853 10761 38887 10795
rect 39773 10761 39807 10795
rect 43177 10761 43211 10795
rect 10701 10693 10735 10727
rect 11958 10693 11992 10727
rect 20269 10693 20303 10727
rect 23121 10693 23155 10727
rect 25513 10693 25547 10727
rect 33793 10693 33827 10727
rect 39313 10693 39347 10727
rect 2145 10625 2179 10659
rect 3985 10625 4019 10659
rect 4252 10625 4286 10659
rect 6929 10625 6963 10659
rect 7196 10625 7230 10659
rect 9505 10625 9539 10659
rect 11713 10625 11747 10659
rect 13921 10625 13955 10659
rect 15025 10625 15059 10659
rect 15669 10625 15703 10659
rect 16313 10625 16347 10659
rect 18889 10625 18923 10659
rect 20085 10625 20119 10659
rect 20729 10625 20763 10659
rect 22109 10625 22143 10659
rect 25421 10625 25455 10659
rect 26065 10625 26099 10659
rect 26249 10625 26283 10659
rect 27261 10625 27295 10659
rect 28641 10625 28675 10659
rect 31033 10625 31067 10659
rect 31309 10625 31343 10659
rect 32321 10625 32355 10659
rect 36001 10625 36035 10659
rect 37473 10625 37507 10659
rect 37729 10625 37763 10659
rect 42809 10625 42843 10659
rect 2973 10557 3007 10591
rect 9781 10557 9815 10591
rect 10885 10557 10919 10591
rect 14105 10557 14139 10591
rect 17417 10557 17451 10591
rect 17509 10557 17543 10591
rect 22845 10557 22879 10591
rect 24869 10557 24903 10591
rect 42901 10557 42935 10591
rect 9137 10489 9171 10523
rect 13553 10489 13587 10523
rect 39589 10489 39623 10523
rect 3525 10421 3559 10455
rect 14841 10421 14875 10455
rect 18705 10421 18739 10455
rect 22201 10421 22235 10455
rect 29929 10421 29963 10455
rect 35081 10421 35115 10455
rect 36369 10421 36403 10455
rect 36553 10421 36587 10455
rect 1777 10217 1811 10251
rect 7941 10217 7975 10251
rect 8401 10217 8435 10251
rect 11713 10217 11747 10251
rect 24685 10217 24719 10251
rect 32045 10217 32079 10251
rect 38209 10217 38243 10251
rect 38761 10217 38795 10251
rect 42901 10217 42935 10251
rect 13737 10149 13771 10183
rect 14933 10149 14967 10183
rect 17141 10149 17175 10183
rect 22937 10149 22971 10183
rect 3157 10081 3191 10115
rect 3249 10081 3283 10115
rect 9597 10081 9631 10115
rect 9781 10081 9815 10115
rect 18521 10081 18555 10115
rect 18705 10081 18739 10115
rect 21465 10081 21499 10115
rect 25697 10081 25731 10115
rect 31861 10081 31895 10115
rect 36829 10081 36863 10115
rect 1593 10013 1627 10047
rect 4537 10013 4571 10047
rect 4793 10013 4827 10047
rect 6561 10013 6595 10047
rect 8585 10013 8619 10047
rect 13369 10013 13403 10047
rect 13553 10013 13587 10047
rect 14657 10013 14691 10047
rect 14749 10013 14783 10047
rect 19441 10013 19475 10047
rect 21189 10013 21223 10047
rect 23581 10013 23615 10047
rect 24593 10013 24627 10047
rect 29745 10013 29779 10047
rect 30001 10013 30035 10047
rect 31769 10013 31803 10047
rect 32689 10013 32723 10047
rect 32781 10013 32815 10047
rect 38669 10013 38703 10047
rect 42809 10013 42843 10047
rect 6806 9945 6840 9979
rect 10425 9945 10459 9979
rect 15669 9945 15703 9979
rect 25964 9945 25998 9979
rect 37074 9945 37108 9979
rect 2697 9877 2731 9911
rect 3065 9877 3099 9911
rect 5917 9877 5951 9911
rect 9137 9877 9171 9911
rect 9505 9877 9539 9911
rect 18061 9877 18095 9911
rect 18429 9877 18463 9911
rect 19533 9877 19567 9911
rect 23673 9877 23707 9911
rect 27077 9877 27111 9911
rect 31125 9877 31159 9911
rect 32965 9877 32999 9911
rect 4721 9673 4755 9707
rect 14289 9673 14323 9707
rect 26433 9673 26467 9707
rect 31677 9673 31711 9707
rect 36737 9673 36771 9707
rect 5549 9605 5583 9639
rect 15200 9605 15234 9639
rect 22845 9605 22879 9639
rect 24593 9605 24627 9639
rect 26157 9605 26191 9639
rect 30665 9605 30699 9639
rect 2237 9537 2271 9571
rect 2881 9537 2915 9571
rect 3341 9537 3375 9571
rect 3608 9537 3642 9571
rect 5641 9537 5675 9571
rect 7205 9537 7239 9571
rect 7472 9537 7506 9571
rect 9689 9537 9723 9571
rect 9956 9537 9990 9571
rect 11897 9537 11931 9571
rect 12909 9537 12943 9571
rect 13176 9537 13210 9571
rect 14933 9537 14967 9571
rect 17141 9537 17175 9571
rect 17601 9537 17635 9571
rect 18613 9537 18647 9571
rect 22569 9537 22603 9571
rect 25421 9537 25455 9571
rect 25881 9537 25915 9571
rect 26065 9537 26099 9571
rect 26249 9537 26283 9571
rect 28457 9537 28491 9571
rect 31585 9537 31619 9571
rect 32505 9537 32539 9571
rect 32965 9537 32999 9571
rect 35817 9537 35851 9571
rect 36921 9537 36955 9571
rect 37749 9537 37783 9571
rect 5825 9469 5859 9503
rect 18245 9469 18279 9503
rect 28733 9469 28767 9503
rect 30205 9469 30239 9503
rect 33241 9469 33275 9503
rect 34989 9469 35023 9503
rect 35909 9469 35943 9503
rect 36001 9469 36035 9503
rect 5181 9401 5215 9435
rect 11069 9401 11103 9435
rect 16313 9401 16347 9435
rect 30941 9401 30975 9435
rect 32321 9401 32355 9435
rect 2053 9333 2087 9367
rect 2697 9333 2731 9367
rect 8585 9333 8619 9367
rect 11713 9333 11747 9367
rect 16957 9333 16991 9367
rect 17693 9333 17727 9367
rect 20039 9333 20073 9367
rect 25237 9333 25271 9367
rect 31125 9333 31159 9367
rect 35449 9333 35483 9367
rect 37565 9333 37599 9367
rect 7849 9129 7883 9163
rect 11621 9129 11655 9163
rect 14289 9129 14323 9163
rect 18843 9129 18877 9163
rect 19441 9129 19475 9163
rect 33057 9129 33091 9163
rect 34161 9129 34195 9163
rect 36369 9129 36403 9163
rect 2697 9061 2731 9095
rect 22017 9061 22051 9095
rect 27261 9061 27295 9095
rect 29101 9061 29135 9095
rect 29837 9061 29871 9095
rect 32413 9061 32447 9095
rect 3341 8993 3375 9027
rect 8493 8993 8527 9027
rect 9781 8993 9815 9027
rect 14933 8993 14967 9027
rect 17417 8993 17451 9027
rect 19993 8993 20027 9027
rect 25053 8993 25087 9027
rect 27813 8993 27847 9027
rect 30481 8993 30515 9027
rect 2237 8925 2271 8959
rect 4077 8925 4111 8959
rect 5641 8925 5675 8959
rect 8309 8925 8343 8959
rect 9321 8925 9355 8959
rect 10048 8925 10082 8959
rect 11805 8925 11839 8959
rect 14657 8925 14691 8959
rect 16405 8925 16439 8959
rect 17049 8925 17083 8959
rect 22661 8925 22695 8959
rect 24777 8925 24811 8959
rect 29009 8925 29043 8959
rect 31033 8925 31067 8959
rect 32965 8925 32999 8959
rect 34345 8925 34379 8959
rect 34989 8925 35023 8959
rect 37473 8925 37507 8959
rect 37729 8925 37763 8959
rect 44373 8925 44407 8959
rect 3065 8857 3099 8891
rect 19809 8857 19843 8891
rect 21741 8857 21775 8891
rect 22906 8857 22940 8891
rect 27721 8857 27755 8891
rect 31300 8857 31334 8891
rect 35234 8857 35268 8891
rect 2053 8789 2087 8823
rect 3157 8789 3191 8823
rect 4629 8789 4663 8823
rect 6929 8789 6963 8823
rect 8217 8789 8251 8823
rect 9137 8789 9171 8823
rect 11161 8789 11195 8823
rect 14749 8789 14783 8823
rect 16221 8789 16255 8823
rect 19901 8789 19935 8823
rect 22201 8789 22235 8823
rect 24041 8789 24075 8823
rect 26525 8789 26559 8823
rect 27629 8789 27663 8823
rect 30205 8789 30239 8823
rect 30297 8789 30331 8823
rect 38853 8789 38887 8823
rect 44189 8789 44223 8823
rect 5365 8585 5399 8619
rect 8217 8585 8251 8619
rect 10057 8585 10091 8619
rect 25605 8585 25639 8619
rect 25973 8585 26007 8619
rect 31033 8585 31067 8619
rect 31493 8585 31527 8619
rect 33977 8585 34011 8619
rect 37473 8585 37507 8619
rect 37933 8585 37967 8619
rect 4230 8517 4264 8551
rect 8944 8517 8978 8551
rect 19993 8517 20027 8551
rect 20821 8517 20855 8551
rect 22201 8517 22235 8551
rect 24777 8517 24811 8551
rect 34866 8517 34900 8551
rect 2145 8449 2179 8483
rect 2401 8449 2435 8483
rect 3985 8449 4019 8483
rect 7113 8449 7147 8483
rect 14197 8449 14231 8483
rect 14381 8449 14415 8483
rect 16129 8449 16163 8483
rect 16865 8449 16899 8483
rect 19073 8449 19107 8483
rect 19165 8449 19199 8483
rect 19717 8449 19751 8483
rect 19901 8449 19935 8483
rect 20085 8449 20119 8483
rect 20729 8449 20763 8483
rect 22017 8449 22051 8483
rect 23121 8449 23155 8483
rect 26065 8449 26099 8483
rect 28080 8449 28114 8483
rect 29909 8449 29943 8483
rect 31677 8449 31711 8483
rect 34161 8449 34195 8483
rect 34621 8449 34655 8483
rect 37841 8449 37875 8483
rect 40509 8449 40543 8483
rect 7665 8381 7699 8415
rect 8677 8381 8711 8415
rect 17141 8381 17175 8415
rect 26157 8381 26191 8415
rect 27813 8381 27847 8415
rect 29653 8381 29687 8415
rect 38025 8381 38059 8415
rect 3525 8313 3559 8347
rect 6929 8313 6963 8347
rect 18613 8313 18647 8347
rect 36001 8313 36035 8347
rect 40601 8313 40635 8347
rect 14289 8245 14323 8279
rect 16221 8245 16255 8279
rect 20269 8245 20303 8279
rect 22385 8245 22419 8279
rect 29193 8245 29227 8279
rect 5365 8041 5399 8075
rect 6469 8041 6503 8075
rect 8401 8041 8435 8075
rect 12449 8041 12483 8075
rect 25053 8041 25087 8075
rect 25697 8041 25731 8075
rect 29745 8041 29779 8075
rect 34897 8041 34931 8075
rect 3985 7905 4019 7939
rect 5917 7905 5951 7939
rect 9137 7905 9171 7939
rect 19993 7905 20027 7939
rect 20085 7905 20119 7939
rect 21557 7905 21591 7939
rect 24685 7905 24719 7939
rect 28733 7905 28767 7939
rect 31401 7905 31435 7939
rect 35357 7905 35391 7939
rect 35541 7905 35575 7939
rect 38209 7905 38243 7939
rect 39497 7905 39531 7939
rect 42257 7905 42291 7939
rect 2053 7837 2087 7871
rect 4252 7837 4286 7871
rect 6929 7837 6963 7871
rect 8033 7837 8067 7871
rect 8217 7837 8251 7871
rect 10977 7837 11011 7871
rect 12081 7837 12115 7871
rect 12265 7837 12299 7871
rect 13277 7837 13311 7871
rect 13369 7837 13403 7871
rect 14565 7837 14599 7871
rect 15393 7837 15427 7871
rect 16037 7837 16071 7871
rect 16497 7837 16531 7871
rect 17141 7837 17175 7871
rect 19717 7837 19751 7871
rect 19901 7837 19935 7871
rect 20269 7837 20303 7871
rect 20913 7837 20947 7871
rect 21097 7837 21131 7871
rect 23581 7837 23615 7871
rect 24777 7837 24811 7871
rect 25605 7837 25639 7871
rect 28917 7837 28951 7871
rect 29929 7837 29963 7871
rect 31125 7837 31159 7871
rect 32597 7837 32631 7871
rect 35265 7837 35299 7871
rect 38301 7837 38335 7871
rect 39221 7837 39255 7871
rect 39313 7837 39347 7871
rect 40049 7837 40083 7871
rect 2320 7769 2354 7803
rect 9382 7769 9416 7803
rect 17417 7769 17451 7803
rect 21824 7769 21858 7803
rect 29101 7769 29135 7803
rect 40325 7769 40359 7803
rect 42533 7769 42567 7803
rect 3433 7701 3467 7735
rect 7573 7701 7607 7735
rect 10517 7701 10551 7735
rect 11621 7701 11655 7735
rect 13553 7701 13587 7735
rect 14657 7701 14691 7735
rect 15209 7701 15243 7735
rect 15853 7701 15887 7735
rect 16589 7701 16623 7735
rect 18889 7701 18923 7735
rect 20453 7701 20487 7735
rect 21005 7701 21039 7735
rect 22937 7701 22971 7735
rect 23397 7701 23431 7735
rect 32413 7701 32447 7735
rect 38669 7701 38703 7735
rect 39497 7701 39531 7735
rect 41797 7701 41831 7735
rect 44005 7701 44039 7735
rect 3893 7497 3927 7531
rect 5641 7497 5675 7531
rect 6929 7497 6963 7531
rect 9137 7497 9171 7531
rect 10057 7497 10091 7531
rect 10517 7497 10551 7531
rect 14473 7497 14507 7531
rect 16865 7497 16899 7531
rect 17325 7497 17359 7531
rect 18153 7497 18187 7531
rect 18521 7497 18555 7531
rect 20269 7497 20303 7531
rect 22217 7497 22251 7531
rect 22385 7497 22419 7531
rect 22845 7497 22879 7531
rect 29929 7497 29963 7531
rect 30757 7497 30791 7531
rect 39497 7497 39531 7531
rect 40617 7497 40651 7531
rect 41245 7497 41279 7531
rect 42717 7497 42751 7531
rect 44189 7497 44223 7531
rect 2605 7429 2639 7463
rect 7849 7429 7883 7463
rect 13360 7429 13394 7463
rect 17233 7429 17267 7463
rect 22017 7429 22051 7463
rect 30849 7429 30883 7463
rect 32566 7429 32600 7463
rect 37565 7429 37599 7463
rect 38761 7429 38795 7463
rect 38945 7429 38979 7463
rect 40417 7429 40451 7463
rect 1777 7361 1811 7395
rect 5549 7361 5583 7395
rect 6745 7361 6779 7395
rect 10425 7361 10459 7395
rect 12633 7361 12667 7395
rect 14933 7361 14967 7395
rect 15117 7361 15151 7395
rect 19625 7361 19659 7395
rect 20085 7361 20119 7395
rect 20729 7361 20763 7395
rect 23029 7361 23063 7395
rect 23765 7361 23799 7395
rect 24685 7361 24719 7395
rect 24961 7361 24995 7395
rect 25605 7361 25639 7395
rect 28816 7361 28850 7395
rect 34345 7361 34379 7395
rect 35541 7361 35575 7395
rect 35725 7361 35759 7395
rect 36093 7361 36127 7395
rect 37473 7361 37507 7395
rect 39037 7361 39071 7395
rect 39681 7361 39715 7395
rect 39865 7361 39899 7395
rect 39957 7361 39991 7395
rect 41429 7361 41463 7395
rect 42625 7361 42659 7395
rect 44373 7361 44407 7395
rect 5825 7293 5859 7327
rect 6561 7293 6595 7327
rect 10609 7293 10643 7327
rect 13093 7293 13127 7327
rect 17509 7293 17543 7327
rect 18613 7293 18647 7327
rect 18797 7293 18831 7327
rect 19993 7293 20027 7327
rect 21005 7293 21039 7327
rect 23949 7293 23983 7327
rect 28549 7293 28583 7327
rect 30941 7293 30975 7327
rect 32321 7293 32355 7327
rect 34253 7293 34287 7327
rect 35817 7293 35851 7327
rect 35909 7293 35943 7327
rect 1593 7225 1627 7259
rect 21281 7225 21315 7259
rect 38761 7225 38795 7259
rect 40785 7225 40819 7259
rect 5181 7157 5215 7191
rect 12449 7157 12483 7191
rect 14933 7157 14967 7191
rect 20085 7157 20119 7191
rect 20821 7157 20855 7191
rect 22201 7157 22235 7191
rect 25697 7157 25731 7191
rect 30389 7157 30423 7191
rect 33701 7157 33735 7191
rect 34713 7157 34747 7191
rect 36277 7157 36311 7191
rect 40601 7157 40635 7191
rect 8585 6953 8619 6987
rect 13737 6953 13771 6987
rect 14657 6953 14691 6987
rect 17601 6953 17635 6987
rect 20913 6953 20947 6987
rect 28641 6953 28675 6987
rect 32413 6953 32447 6987
rect 39129 6953 39163 6987
rect 40233 6953 40267 6987
rect 11713 6885 11747 6919
rect 17049 6885 17083 6919
rect 2697 6817 2731 6851
rect 3985 6817 4019 6851
rect 15393 6817 15427 6851
rect 17693 6817 17727 6851
rect 18889 6817 18923 6851
rect 19993 6817 20027 6851
rect 32965 6817 32999 6851
rect 40969 6817 41003 6851
rect 41153 6817 41187 6851
rect 41705 6817 41739 6851
rect 7205 6749 7239 6783
rect 9505 6749 9539 6783
rect 9781 6749 9815 6783
rect 11713 6749 11747 6783
rect 11897 6749 11931 6783
rect 12357 6749 12391 6783
rect 12613 6749 12647 6783
rect 14289 6749 14323 6783
rect 15301 6749 15335 6783
rect 17230 6749 17264 6783
rect 18153 6749 18187 6783
rect 18337 6749 18371 6783
rect 18429 6749 18463 6783
rect 18521 6749 18555 6783
rect 18705 6749 18739 6783
rect 19625 6749 19659 6783
rect 19717 6749 19751 6783
rect 20085 6749 20119 6783
rect 20821 6749 20855 6783
rect 21005 6749 21039 6783
rect 21741 6749 21775 6783
rect 21833 6749 21867 6783
rect 21925 6749 21959 6783
rect 22109 6749 22143 6783
rect 22661 6749 22695 6783
rect 24041 6749 24075 6783
rect 24593 6749 24627 6783
rect 28181 6749 28215 6783
rect 28825 6749 28859 6783
rect 31217 6749 31251 6783
rect 32781 6749 32815 6783
rect 33609 6749 33643 6783
rect 33977 6749 34011 6783
rect 35265 6749 35299 6783
rect 35413 6749 35447 6783
rect 35541 6749 35575 6783
rect 35771 6749 35805 6783
rect 38301 6749 38335 6783
rect 38485 6749 38519 6783
rect 40877 6749 40911 6783
rect 41613 6749 41647 6783
rect 42257 6749 42291 6783
rect 2513 6681 2547 6715
rect 4230 6681 4264 6715
rect 7472 6681 7506 6715
rect 24869 6681 24903 6715
rect 32873 6681 32907 6715
rect 33793 6681 33827 6715
rect 33885 6681 33919 6715
rect 35633 6681 35667 6715
rect 38945 6681 38979 6715
rect 40049 6681 40083 6715
rect 40265 6681 40299 6715
rect 2145 6613 2179 6647
rect 2605 6613 2639 6647
rect 5365 6613 5399 6647
rect 9219 6613 9253 6647
rect 9689 6613 9723 6647
rect 14657 6613 14691 6647
rect 14841 6613 14875 6647
rect 17233 6613 17267 6647
rect 19441 6613 19475 6647
rect 21465 6613 21499 6647
rect 22753 6613 22787 6647
rect 23857 6613 23891 6647
rect 26341 6613 26375 6647
rect 27997 6613 28031 6647
rect 31309 6613 31343 6647
rect 34161 6613 34195 6647
rect 35909 6613 35943 6647
rect 38393 6613 38427 6647
rect 39145 6613 39179 6647
rect 39313 6613 39347 6647
rect 40417 6613 40451 6647
rect 41153 6613 41187 6647
rect 42349 6613 42383 6647
rect 2881 6409 2915 6443
rect 4721 6409 4755 6443
rect 9321 6409 9355 6443
rect 11161 6409 11195 6443
rect 13553 6409 13587 6443
rect 15041 6409 15075 6443
rect 20269 6409 20303 6443
rect 23397 6409 23431 6443
rect 24869 6409 24903 6443
rect 25237 6409 25271 6443
rect 38577 6409 38611 6443
rect 8186 6341 8220 6375
rect 12173 6341 12207 6375
rect 12389 6341 12423 6375
rect 13369 6341 13403 6375
rect 14013 6341 14047 6375
rect 14841 6341 14875 6375
rect 17693 6341 17727 6375
rect 18889 6341 18923 6375
rect 22262 6341 22296 6375
rect 27721 6341 27755 6375
rect 28794 6341 28828 6375
rect 32781 6341 32815 6375
rect 42717 6341 42751 6375
rect 1777 6273 1811 6307
rect 2329 6273 2363 6307
rect 3341 6273 3375 6307
rect 3608 6273 3642 6307
rect 7941 6273 7975 6307
rect 9781 6273 9815 6307
rect 10048 6273 10082 6307
rect 14197 6273 14231 6307
rect 19717 6273 19751 6307
rect 19901 6273 19935 6307
rect 19993 6273 20027 6307
rect 20085 6273 20119 6307
rect 20913 6273 20947 6307
rect 22017 6273 22051 6307
rect 24225 6273 24259 6307
rect 27629 6273 27663 6307
rect 31493 6273 31527 6307
rect 31677 6273 31711 6307
rect 31769 6273 31803 6307
rect 33057 6273 33091 6307
rect 33149 6273 33183 6307
rect 33241 6273 33275 6307
rect 33425 6273 33459 6307
rect 34069 6273 34103 6307
rect 34161 6273 34195 6307
rect 34437 6273 34471 6307
rect 34989 6273 35023 6307
rect 35081 6273 35115 6307
rect 35173 6273 35207 6307
rect 35909 6273 35943 6307
rect 36093 6273 36127 6307
rect 38485 6273 38519 6307
rect 39497 6273 39531 6307
rect 39589 6273 39623 6307
rect 40325 6273 40359 6307
rect 42625 6273 42659 6307
rect 17785 6205 17819 6239
rect 17969 6205 18003 6239
rect 18981 6205 19015 6239
rect 19165 6205 19199 6239
rect 21005 6205 21039 6239
rect 25329 6205 25363 6239
rect 25513 6205 25547 6239
rect 27813 6205 27847 6239
rect 28549 6205 28583 6239
rect 33885 6205 33919 6239
rect 34345 6205 34379 6239
rect 39313 6205 39347 6239
rect 39405 6205 39439 6239
rect 40601 6205 40635 6239
rect 12541 6137 12575 6171
rect 13001 6137 13035 6171
rect 14381 6137 14415 6171
rect 21281 6137 21315 6171
rect 24317 6137 24351 6171
rect 12357 6069 12391 6103
rect 13369 6069 13403 6103
rect 15025 6069 15059 6103
rect 15209 6069 15243 6103
rect 17325 6069 17359 6103
rect 18521 6069 18555 6103
rect 27261 6069 27295 6103
rect 29929 6069 29963 6103
rect 35357 6069 35391 6103
rect 36001 6069 36035 6103
rect 39129 6069 39163 6103
rect 42073 6069 42107 6103
rect 3249 5865 3283 5899
rect 5365 5865 5399 5899
rect 11713 5865 11747 5899
rect 14381 5865 14415 5899
rect 14473 5865 14507 5899
rect 18245 5865 18279 5899
rect 29745 5865 29779 5899
rect 32689 5865 32723 5899
rect 34069 5865 34103 5899
rect 34989 5865 35023 5899
rect 40141 5865 40175 5899
rect 42625 5865 42659 5899
rect 28181 5797 28215 5831
rect 35633 5797 35667 5831
rect 39497 5797 39531 5831
rect 3985 5729 4019 5763
rect 5825 5729 5859 5763
rect 14565 5729 14599 5763
rect 16497 5729 16531 5763
rect 21281 5729 21315 5763
rect 26801 5729 26835 5763
rect 30297 5729 30331 5763
rect 33333 5729 33367 5763
rect 34161 5729 34195 5763
rect 37749 5729 37783 5763
rect 40325 5729 40359 5763
rect 40877 5729 40911 5763
rect 2789 5661 2823 5695
rect 3433 5661 3467 5695
rect 6009 5661 6043 5695
rect 9597 5661 9631 5695
rect 9781 5661 9815 5695
rect 10425 5661 10459 5695
rect 14289 5661 14323 5695
rect 16037 5661 16071 5695
rect 18705 5661 18739 5695
rect 20453 5661 20487 5695
rect 20545 5661 20579 5695
rect 20637 5661 20671 5695
rect 20821 5661 20855 5695
rect 26341 5661 26375 5695
rect 28825 5661 28859 5695
rect 30113 5661 30147 5695
rect 31401 5661 31435 5695
rect 32045 5661 32079 5695
rect 32229 5661 32263 5695
rect 32870 5661 32904 5695
rect 33241 5661 33275 5695
rect 34897 5661 34931 5695
rect 35541 5661 35575 5695
rect 40049 5661 40083 5695
rect 44097 5661 44131 5695
rect 4230 5593 4264 5627
rect 16773 5593 16807 5627
rect 18797 5593 18831 5627
rect 20177 5593 20211 5627
rect 21526 5593 21560 5627
rect 27046 5593 27080 5627
rect 30205 5593 30239 5627
rect 31493 5593 31527 5627
rect 33793 5593 33827 5627
rect 34253 5593 34287 5627
rect 36553 5593 36587 5627
rect 36737 5593 36771 5627
rect 38025 5593 38059 5627
rect 41153 5593 41187 5627
rect 2605 5525 2639 5559
rect 6193 5525 6227 5559
rect 9965 5525 9999 5559
rect 15853 5525 15887 5559
rect 22661 5525 22695 5559
rect 26157 5525 26191 5559
rect 28641 5525 28675 5559
rect 32137 5525 32171 5559
rect 32873 5525 32907 5559
rect 33885 5525 33919 5559
rect 36921 5525 36955 5559
rect 40325 5525 40359 5559
rect 44281 5525 44315 5559
rect 5365 5321 5399 5355
rect 13645 5321 13679 5355
rect 18613 5321 18647 5355
rect 21097 5321 21131 5355
rect 24409 5321 24443 5355
rect 29929 5321 29963 5355
rect 35081 5321 35115 5355
rect 36211 5321 36245 5355
rect 38695 5321 38729 5355
rect 40509 5321 40543 5355
rect 41153 5321 41187 5355
rect 28641 5253 28675 5287
rect 33793 5253 33827 5287
rect 36001 5253 36035 5287
rect 38485 5253 38519 5287
rect 40325 5253 40359 5287
rect 3985 5185 4019 5219
rect 4252 5185 4286 5219
rect 9229 5185 9263 5219
rect 9413 5185 9447 5219
rect 12265 5185 12299 5219
rect 12532 5185 12566 5219
rect 14105 5185 14139 5219
rect 15301 5185 15335 5219
rect 15485 5185 15519 5219
rect 16865 5185 16899 5219
rect 19257 5185 19291 5219
rect 21005 5185 21039 5219
rect 21189 5185 21223 5219
rect 23029 5185 23063 5219
rect 23296 5185 23330 5219
rect 32413 5185 32447 5219
rect 32505 5185 32539 5219
rect 32689 5185 32723 5219
rect 32781 5185 32815 5219
rect 32873 5185 32907 5219
rect 37841 5185 37875 5219
rect 37933 5185 37967 5219
rect 39497 5185 39531 5219
rect 40601 5185 40635 5219
rect 41061 5185 41095 5219
rect 41245 5185 41279 5219
rect 42993 5185 43027 5219
rect 1593 5117 1627 5151
rect 1869 5117 1903 5151
rect 14197 5117 14231 5151
rect 14381 5117 14415 5151
rect 17141 5117 17175 5151
rect 19073 5049 19107 5083
rect 36369 5049 36403 5083
rect 39313 5049 39347 5083
rect 40325 5049 40359 5083
rect 9597 4981 9631 5015
rect 14289 4981 14323 5015
rect 15669 4981 15703 5015
rect 32413 4981 32447 5015
rect 36185 4981 36219 5015
rect 38669 4981 38703 5015
rect 38853 4981 38887 5015
rect 42809 4981 42843 5015
rect 13185 4777 13219 4811
rect 18429 4777 18463 4811
rect 28549 4777 28583 4811
rect 32965 4777 32999 4811
rect 37197 4777 37231 4811
rect 38393 4777 38427 4811
rect 23029 4709 23063 4743
rect 4905 4641 4939 4675
rect 20545 4641 20579 4675
rect 20821 4641 20855 4675
rect 22293 4641 22327 4675
rect 22753 4641 22787 4675
rect 27169 4641 27203 4675
rect 31217 4641 31251 4675
rect 31493 4641 31527 4675
rect 33425 4641 33459 4675
rect 35449 4641 35483 4675
rect 5089 4573 5123 4607
rect 11805 4573 11839 4607
rect 15209 4573 15243 4607
rect 15669 4573 15703 4607
rect 18337 4573 18371 4607
rect 19441 4573 19475 4607
rect 27436 4573 27470 4607
rect 33793 4573 33827 4607
rect 33885 4573 33919 4607
rect 37657 4573 37691 4607
rect 38577 4573 38611 4607
rect 44097 4573 44131 4607
rect 12050 4505 12084 4539
rect 17417 4505 17451 4539
rect 35725 4505 35759 4539
rect 37749 4505 37783 4539
rect 5273 4437 5307 4471
rect 15025 4437 15059 4471
rect 19533 4437 19567 4471
rect 23213 4437 23247 4471
rect 33701 4437 33735 4471
rect 44281 4437 44315 4471
rect 13093 4233 13127 4267
rect 14841 4165 14875 4199
rect 27813 4165 27847 4199
rect 13001 4097 13035 4131
rect 13185 4097 13219 4131
rect 16865 4097 16899 4131
rect 17509 4097 17543 4131
rect 22017 4097 22051 4131
rect 22109 4097 22143 4131
rect 22937 4097 22971 4131
rect 27905 4097 27939 4131
rect 31585 4097 31619 4131
rect 32505 4097 32539 4131
rect 33425 4097 33459 4131
rect 33517 4097 33551 4131
rect 35265 4097 35299 4131
rect 36369 4097 36403 4131
rect 37473 4097 37507 4131
rect 14565 4029 14599 4063
rect 18153 4029 18187 4063
rect 18429 4029 18463 4063
rect 19901 4029 19935 4063
rect 27997 4029 28031 4063
rect 32689 4029 32723 4063
rect 32781 4029 32815 4063
rect 36277 4029 36311 4063
rect 37749 4029 37783 4063
rect 16313 3961 16347 3995
rect 22753 3961 22787 3995
rect 27445 3961 27479 3995
rect 35081 3961 35115 3995
rect 36737 3961 36771 3995
rect 16957 3893 16991 3927
rect 17601 3893 17635 3927
rect 31677 3893 31711 3927
rect 32321 3893 32355 3927
rect 39221 3893 39255 3927
rect 31388 3689 31422 3723
rect 32873 3689 32907 3723
rect 37565 3689 37599 3723
rect 22385 3621 22419 3655
rect 1777 3485 1811 3519
rect 5917 3485 5951 3519
rect 14565 3485 14599 3519
rect 15669 3485 15703 3519
rect 16681 3485 16715 3519
rect 17049 3485 17083 3519
rect 19441 3485 19475 3519
rect 31125 3485 31159 3519
rect 37473 3485 37507 3519
rect 44373 3485 44407 3519
rect 18475 3417 18509 3451
rect 22109 3417 22143 3451
rect 5733 3349 5767 3383
rect 14657 3349 14691 3383
rect 19533 3349 19567 3383
rect 9689 3145 9723 3179
rect 16267 3145 16301 3179
rect 16957 3145 16991 3179
rect 17601 3145 17635 3179
rect 20315 3145 20349 3179
rect 33885 3145 33919 3179
rect 44189 3145 44223 3179
rect 7757 3009 7791 3043
rect 9505 3009 9539 3043
rect 14013 3009 14047 3043
rect 14473 3009 14507 3043
rect 14841 3009 14875 3043
rect 16865 3009 16899 3043
rect 17509 3009 17543 3043
rect 18521 3009 18555 3043
rect 18889 3009 18923 3043
rect 22477 3009 22511 3043
rect 34253 3009 34287 3043
rect 44373 3009 44407 3043
rect 1777 2805 1811 2839
rect 7573 2805 7607 2839
rect 13829 2805 13863 2839
rect 22293 2805 22327 2839
rect 34437 2805 34471 2839
rect 16957 2601 16991 2635
rect 27353 2601 27387 2635
rect 37473 2601 37507 2635
rect 43453 2601 43487 2635
rect 42901 2533 42935 2567
rect 2421 2465 2455 2499
rect 13185 2465 13219 2499
rect 17785 2465 17819 2499
rect 32597 2465 32631 2499
rect 1777 2397 1811 2431
rect 4169 2397 4203 2431
rect 4813 2397 4847 2431
rect 6561 2397 6595 2431
rect 8033 2397 8067 2431
rect 9781 2397 9815 2431
rect 11897 2397 11931 2431
rect 12909 2397 12943 2431
rect 15669 2397 15703 2431
rect 16865 2397 16899 2431
rect 17509 2397 17543 2431
rect 19625 2397 19659 2431
rect 20913 2397 20947 2431
rect 22661 2397 22695 2431
rect 24777 2397 24811 2431
rect 26065 2397 26099 2431
rect 27169 2397 27203 2431
rect 29929 2397 29963 2431
rect 30573 2397 30607 2431
rect 32321 2397 32355 2431
rect 35541 2397 35575 2431
rect 37657 2397 37691 2431
rect 38945 2397 38979 2431
rect 40233 2397 40267 2431
rect 43637 2397 43671 2431
rect 44097 2397 44131 2431
rect 42717 2329 42751 2363
rect 6745 2261 6779 2295
rect 9965 2261 9999 2295
rect 22845 2261 22879 2295
rect 25881 2261 25915 2295
rect 35725 2261 35759 2295
rect 44281 2261 44315 2295
<< metal1 >>
rect 34146 19048 34152 19100
rect 34204 19088 34210 19100
rect 35066 19088 35072 19100
rect 34204 19060 35072 19088
rect 34204 19048 34210 19060
rect 35066 19048 35072 19060
rect 35124 19048 35130 19100
rect 41874 19048 41880 19100
rect 41932 19088 41938 19100
rect 42794 19088 42800 19100
rect 41932 19060 42800 19088
rect 41932 19048 41938 19060
rect 42794 19048 42800 19060
rect 42852 19048 42858 19100
rect 43714 17960 43720 18012
rect 43772 18000 43778 18012
rect 45002 18000 45008 18012
rect 43772 17972 45008 18000
rect 43772 17960 43778 17972
rect 45002 17960 45008 17972
rect 45060 17960 45066 18012
rect 1104 17434 45051 17456
rect 1104 17382 11896 17434
rect 11948 17382 11960 17434
rect 12012 17382 12024 17434
rect 12076 17382 12088 17434
rect 12140 17382 12152 17434
rect 12204 17382 22843 17434
rect 22895 17382 22907 17434
rect 22959 17382 22971 17434
rect 23023 17382 23035 17434
rect 23087 17382 23099 17434
rect 23151 17382 33790 17434
rect 33842 17382 33854 17434
rect 33906 17382 33918 17434
rect 33970 17382 33982 17434
rect 34034 17382 34046 17434
rect 34098 17382 44737 17434
rect 44789 17382 44801 17434
rect 44853 17382 44865 17434
rect 44917 17382 44929 17434
rect 44981 17382 44993 17434
rect 45045 17382 45051 17434
rect 1104 17360 45051 17382
rect 17402 17280 17408 17332
rect 17460 17320 17466 17332
rect 17681 17323 17739 17329
rect 17681 17320 17693 17323
rect 17460 17292 17693 17320
rect 17460 17280 17466 17292
rect 17681 17289 17693 17292
rect 17727 17289 17739 17323
rect 17681 17283 17739 17289
rect 20714 17280 20720 17332
rect 20772 17320 20778 17332
rect 20901 17323 20959 17329
rect 20901 17320 20913 17323
rect 20772 17292 20913 17320
rect 20772 17280 20778 17292
rect 20901 17289 20913 17292
rect 20947 17289 20959 17323
rect 20901 17283 20959 17289
rect 40586 17280 40592 17332
rect 40644 17320 40650 17332
rect 40865 17323 40923 17329
rect 40865 17320 40877 17323
rect 40644 17292 40877 17320
rect 40644 17280 40650 17292
rect 40865 17289 40877 17292
rect 40911 17289 40923 17323
rect 40865 17283 40923 17289
rect 44266 17280 44272 17332
rect 44324 17280 44330 17332
rect 1302 17212 1308 17264
rect 1360 17252 1366 17264
rect 1673 17255 1731 17261
rect 1673 17252 1685 17255
rect 1360 17224 1685 17252
rect 1360 17212 1366 17224
rect 1673 17221 1685 17224
rect 1719 17221 1731 17255
rect 1673 17215 1731 17221
rect 3234 17212 3240 17264
rect 3292 17212 3298 17264
rect 4522 17212 4528 17264
rect 4580 17252 4586 17264
rect 4709 17255 4767 17261
rect 4709 17252 4721 17255
rect 4580 17224 4721 17252
rect 4580 17212 4586 17224
rect 4709 17221 4721 17224
rect 4755 17221 4767 17255
rect 4709 17215 4767 17221
rect 11054 17212 11060 17264
rect 11112 17252 11118 17264
rect 11793 17255 11851 17261
rect 11793 17252 11805 17255
rect 11112 17224 11805 17252
rect 11112 17212 11118 17224
rect 11793 17221 11805 17224
rect 11839 17221 11851 17255
rect 11793 17215 11851 17221
rect 16114 17212 16120 17264
rect 16172 17212 16178 17264
rect 32214 17212 32220 17264
rect 32272 17252 32278 17264
rect 32401 17255 32459 17261
rect 32401 17252 32413 17255
rect 32272 17224 32413 17252
rect 32272 17212 32278 17224
rect 32401 17221 32413 17224
rect 32447 17221 32459 17255
rect 32401 17215 32459 17221
rect 38654 17212 38660 17264
rect 38712 17252 38718 17264
rect 38841 17255 38899 17261
rect 38841 17252 38853 17255
rect 38712 17224 38853 17252
rect 38712 17212 38718 17224
rect 38841 17221 38853 17224
rect 38887 17221 38899 17255
rect 38841 17215 38899 17221
rect 934 17144 940 17196
rect 992 17184 998 17196
rect 2409 17187 2467 17193
rect 2409 17184 2421 17187
rect 992 17156 2421 17184
rect 992 17144 998 17156
rect 2409 17153 2421 17156
rect 2455 17153 2467 17187
rect 2409 17147 2467 17153
rect 6454 17144 6460 17196
rect 6512 17184 6518 17196
rect 6733 17187 6791 17193
rect 6733 17184 6745 17187
rect 6512 17156 6745 17184
rect 6512 17144 6518 17156
rect 6733 17153 6745 17156
rect 6779 17153 6791 17187
rect 6733 17147 6791 17153
rect 7742 17144 7748 17196
rect 7800 17184 7806 17196
rect 8021 17187 8079 17193
rect 8021 17184 8033 17187
rect 7800 17156 8033 17184
rect 7800 17144 7806 17156
rect 8021 17153 8033 17156
rect 8067 17153 8079 17187
rect 8021 17147 8079 17153
rect 9674 17144 9680 17196
rect 9732 17184 9738 17196
rect 9953 17187 10011 17193
rect 9953 17184 9965 17187
rect 9732 17156 9965 17184
rect 9732 17144 9738 17156
rect 9953 17153 9965 17156
rect 9999 17153 10011 17187
rect 9953 17147 10011 17153
rect 12894 17144 12900 17196
rect 12952 17184 12958 17196
rect 13173 17187 13231 17193
rect 13173 17184 13185 17187
rect 12952 17156 13185 17184
rect 12952 17144 12958 17156
rect 13173 17153 13185 17156
rect 13219 17153 13231 17187
rect 13173 17147 13231 17153
rect 14182 17144 14188 17196
rect 14240 17184 14246 17196
rect 14461 17187 14519 17193
rect 14461 17184 14473 17187
rect 14240 17156 14473 17184
rect 14240 17144 14246 17156
rect 14461 17153 14473 17156
rect 14507 17153 14519 17187
rect 14461 17147 14519 17153
rect 16574 17144 16580 17196
rect 16632 17184 16638 17196
rect 17497 17187 17555 17193
rect 17497 17184 17509 17187
rect 16632 17156 17509 17184
rect 16632 17144 16638 17156
rect 17497 17153 17509 17156
rect 17543 17153 17555 17187
rect 17497 17147 17555 17153
rect 19334 17144 19340 17196
rect 19392 17184 19398 17196
rect 19613 17187 19671 17193
rect 19613 17184 19625 17187
rect 19392 17156 19625 17184
rect 19392 17144 19398 17156
rect 19613 17153 19625 17156
rect 19659 17153 19671 17187
rect 19613 17147 19671 17153
rect 20714 17144 20720 17196
rect 20772 17144 20778 17196
rect 22554 17144 22560 17196
rect 22612 17184 22618 17196
rect 22833 17187 22891 17193
rect 22833 17184 22845 17187
rect 22612 17156 22845 17184
rect 22612 17144 22618 17156
rect 22833 17153 22845 17156
rect 22879 17153 22891 17187
rect 22833 17147 22891 17153
rect 23842 17144 23848 17196
rect 23900 17184 23906 17196
rect 24765 17187 24823 17193
rect 24765 17184 24777 17187
rect 23900 17156 24777 17184
rect 23900 17144 23906 17156
rect 24765 17153 24777 17156
rect 24811 17153 24823 17187
rect 24765 17147 24823 17153
rect 25774 17144 25780 17196
rect 25832 17184 25838 17196
rect 26053 17187 26111 17193
rect 26053 17184 26065 17187
rect 25832 17156 26065 17184
rect 25832 17144 25838 17156
rect 26053 17153 26065 17156
rect 26099 17153 26111 17187
rect 26053 17147 26111 17153
rect 27706 17144 27712 17196
rect 27764 17184 27770 17196
rect 27985 17187 28043 17193
rect 27985 17184 27997 17187
rect 27764 17156 27997 17184
rect 27764 17144 27770 17156
rect 27985 17153 27997 17156
rect 28031 17153 28043 17187
rect 27985 17147 28043 17153
rect 28994 17144 29000 17196
rect 29052 17184 29058 17196
rect 29917 17187 29975 17193
rect 29917 17184 29929 17187
rect 29052 17156 29929 17184
rect 29052 17144 29058 17156
rect 29917 17153 29929 17156
rect 29963 17153 29975 17187
rect 29917 17147 29975 17153
rect 30926 17144 30932 17196
rect 30984 17184 30990 17196
rect 31205 17187 31263 17193
rect 31205 17184 31217 17187
rect 30984 17156 31217 17184
rect 30984 17144 30990 17156
rect 31205 17153 31217 17156
rect 31251 17153 31263 17187
rect 31205 17147 31263 17153
rect 35066 17144 35072 17196
rect 35124 17144 35130 17196
rect 35434 17144 35440 17196
rect 35492 17184 35498 17196
rect 35713 17187 35771 17193
rect 35713 17184 35725 17187
rect 35492 17156 35725 17184
rect 35492 17144 35498 17156
rect 35713 17153 35725 17156
rect 35759 17153 35771 17187
rect 35713 17147 35771 17153
rect 37366 17144 37372 17196
rect 37424 17184 37430 17196
rect 37645 17187 37703 17193
rect 37645 17184 37657 17187
rect 37424 17156 37657 17184
rect 37424 17144 37430 17156
rect 37645 17153 37657 17156
rect 37691 17153 37703 17187
rect 37645 17147 37703 17153
rect 40678 17144 40684 17196
rect 40736 17144 40742 17196
rect 42794 17144 42800 17196
rect 42852 17144 42858 17196
rect 43625 17187 43683 17193
rect 43625 17153 43637 17187
rect 43671 17184 43683 17187
rect 43806 17184 43812 17196
rect 43671 17156 43812 17184
rect 43671 17153 43683 17156
rect 43625 17147 43683 17153
rect 43806 17144 43812 17156
rect 43864 17144 43870 17196
rect 44082 17144 44088 17196
rect 44140 17144 44146 17196
rect 1854 17008 1860 17060
rect 1912 17008 1918 17060
rect 3421 17051 3479 17057
rect 3421 17017 3433 17051
rect 3467 17048 3479 17051
rect 4062 17048 4068 17060
rect 3467 17020 4068 17048
rect 3467 17017 3479 17020
rect 3421 17011 3479 17017
rect 4062 17008 4068 17020
rect 4120 17008 4126 17060
rect 11977 17051 12035 17057
rect 11977 17017 11989 17051
rect 12023 17048 12035 17051
rect 13078 17048 13084 17060
rect 12023 17020 13084 17048
rect 12023 17017 12035 17020
rect 11977 17011 12035 17017
rect 13078 17008 13084 17020
rect 13136 17008 13142 17060
rect 16298 17008 16304 17060
rect 16356 17008 16362 17060
rect 2498 16940 2504 16992
rect 2556 16940 2562 16992
rect 4798 16940 4804 16992
rect 4856 16940 4862 16992
rect 9769 16983 9827 16989
rect 9769 16949 9781 16983
rect 9815 16980 9827 16983
rect 9950 16980 9956 16992
rect 9815 16952 9956 16980
rect 9815 16949 9827 16952
rect 9769 16943 9827 16949
rect 9950 16940 9956 16952
rect 10008 16940 10014 16992
rect 23290 16940 23296 16992
rect 23348 16980 23354 16992
rect 24581 16983 24639 16989
rect 24581 16980 24593 16983
rect 23348 16952 24593 16980
rect 23348 16940 23354 16952
rect 24581 16949 24593 16952
rect 24627 16949 24639 16983
rect 24581 16943 24639 16949
rect 30926 16940 30932 16992
rect 30984 16980 30990 16992
rect 31021 16983 31079 16989
rect 31021 16980 31033 16983
rect 30984 16952 31033 16980
rect 30984 16940 30990 16952
rect 31021 16949 31033 16952
rect 31067 16949 31079 16983
rect 31021 16943 31079 16949
rect 32214 16940 32220 16992
rect 32272 16980 32278 16992
rect 32493 16983 32551 16989
rect 32493 16980 32505 16983
rect 32272 16952 32505 16980
rect 32272 16940 32278 16952
rect 32493 16949 32505 16952
rect 32539 16949 32551 16983
rect 32493 16943 32551 16949
rect 34882 16940 34888 16992
rect 34940 16940 34946 16992
rect 38930 16940 38936 16992
rect 38988 16940 38994 16992
rect 1104 16890 44896 16912
rect 1104 16838 6423 16890
rect 6475 16838 6487 16890
rect 6539 16838 6551 16890
rect 6603 16838 6615 16890
rect 6667 16838 6679 16890
rect 6731 16838 17370 16890
rect 17422 16838 17434 16890
rect 17486 16838 17498 16890
rect 17550 16838 17562 16890
rect 17614 16838 17626 16890
rect 17678 16838 28317 16890
rect 28369 16838 28381 16890
rect 28433 16838 28445 16890
rect 28497 16838 28509 16890
rect 28561 16838 28573 16890
rect 28625 16838 39264 16890
rect 39316 16838 39328 16890
rect 39380 16838 39392 16890
rect 39444 16838 39456 16890
rect 39508 16838 39520 16890
rect 39572 16838 44896 16890
rect 1104 16816 44896 16838
rect 2498 16736 2504 16788
rect 2556 16776 2562 16788
rect 34790 16776 34796 16788
rect 2556 16748 34796 16776
rect 2556 16736 2562 16748
rect 34790 16736 34796 16748
rect 34848 16736 34854 16788
rect 43714 16736 43720 16788
rect 43772 16736 43778 16788
rect 44361 16779 44419 16785
rect 44361 16745 44373 16779
rect 44407 16776 44419 16779
rect 45094 16776 45100 16788
rect 44407 16748 45100 16776
rect 44407 16745 44419 16748
rect 44361 16739 44419 16745
rect 45094 16736 45100 16748
rect 45152 16736 45158 16788
rect 1857 16643 1915 16649
rect 1857 16609 1869 16643
rect 1903 16640 1915 16643
rect 1946 16640 1952 16652
rect 1903 16612 1952 16640
rect 1903 16609 1915 16612
rect 1857 16603 1915 16609
rect 1946 16600 1952 16612
rect 2004 16600 2010 16652
rect 14 16532 20 16584
rect 72 16572 78 16584
rect 1673 16575 1731 16581
rect 1673 16572 1685 16575
rect 72 16544 1685 16572
rect 72 16532 78 16544
rect 1673 16541 1685 16544
rect 1719 16541 1731 16575
rect 1673 16535 1731 16541
rect 14182 16532 14188 16584
rect 14240 16572 14246 16584
rect 14553 16575 14611 16581
rect 14553 16572 14565 16575
rect 14240 16544 14565 16572
rect 14240 16532 14246 16544
rect 14553 16541 14565 16544
rect 14599 16541 14611 16575
rect 14553 16535 14611 16541
rect 27614 16532 27620 16584
rect 27672 16572 27678 16584
rect 28537 16575 28595 16581
rect 28537 16572 28549 16575
rect 27672 16544 28549 16572
rect 27672 16532 27678 16544
rect 28537 16541 28549 16544
rect 28583 16541 28595 16575
rect 28537 16535 28595 16541
rect 14369 16439 14427 16445
rect 14369 16405 14381 16439
rect 14415 16436 14427 16439
rect 20714 16436 20720 16448
rect 14415 16408 20720 16436
rect 14415 16405 14427 16408
rect 14369 16399 14427 16405
rect 20714 16396 20720 16408
rect 20772 16396 20778 16448
rect 28353 16439 28411 16445
rect 28353 16405 28365 16439
rect 28399 16436 28411 16439
rect 40678 16436 40684 16448
rect 28399 16408 40684 16436
rect 28399 16405 28411 16408
rect 28353 16399 28411 16405
rect 40678 16396 40684 16408
rect 40736 16396 40742 16448
rect 1104 16346 45051 16368
rect 1104 16294 11896 16346
rect 11948 16294 11960 16346
rect 12012 16294 12024 16346
rect 12076 16294 12088 16346
rect 12140 16294 12152 16346
rect 12204 16294 22843 16346
rect 22895 16294 22907 16346
rect 22959 16294 22971 16346
rect 23023 16294 23035 16346
rect 23087 16294 23099 16346
rect 23151 16294 33790 16346
rect 33842 16294 33854 16346
rect 33906 16294 33918 16346
rect 33970 16294 33982 16346
rect 34034 16294 34046 16346
rect 34098 16294 44737 16346
rect 44789 16294 44801 16346
rect 44853 16294 44865 16346
rect 44917 16294 44929 16346
rect 44981 16294 44993 16346
rect 45045 16294 45051 16346
rect 1104 16272 45051 16294
rect 42981 16235 43039 16241
rect 42981 16201 42993 16235
rect 43027 16232 43039 16235
rect 44082 16232 44088 16244
rect 43027 16204 44088 16232
rect 43027 16201 43039 16204
rect 42981 16195 43039 16201
rect 44082 16192 44088 16204
rect 44140 16192 44146 16244
rect 1026 16056 1032 16108
rect 1084 16096 1090 16108
rect 1765 16099 1823 16105
rect 1765 16096 1777 16099
rect 1084 16068 1777 16096
rect 1084 16056 1090 16068
rect 1765 16065 1777 16068
rect 1811 16065 1823 16099
rect 42797 16099 42855 16105
rect 42797 16096 42809 16099
rect 1765 16059 1823 16065
rect 26206 16068 42809 16096
rect 6822 15852 6828 15904
rect 6880 15892 6886 15904
rect 26206 15892 26234 16068
rect 42797 16065 42809 16068
rect 42843 16096 42855 16099
rect 43257 16099 43315 16105
rect 43257 16096 43269 16099
rect 42843 16068 43269 16096
rect 42843 16065 42855 16068
rect 42797 16059 42855 16065
rect 43257 16065 43269 16068
rect 43303 16065 43315 16099
rect 43257 16059 43315 16065
rect 6880 15864 26234 15892
rect 6880 15852 6886 15864
rect 44358 15852 44364 15904
rect 44416 15852 44422 15904
rect 1104 15802 44896 15824
rect 1104 15750 6423 15802
rect 6475 15750 6487 15802
rect 6539 15750 6551 15802
rect 6603 15750 6615 15802
rect 6667 15750 6679 15802
rect 6731 15750 17370 15802
rect 17422 15750 17434 15802
rect 17486 15750 17498 15802
rect 17550 15750 17562 15802
rect 17614 15750 17626 15802
rect 17678 15750 28317 15802
rect 28369 15750 28381 15802
rect 28433 15750 28445 15802
rect 28497 15750 28509 15802
rect 28561 15750 28573 15802
rect 28625 15750 39264 15802
rect 39316 15750 39328 15802
rect 39380 15750 39392 15802
rect 39444 15750 39456 15802
rect 39508 15750 39520 15802
rect 39572 15750 44896 15802
rect 1104 15728 44896 15750
rect 32309 15691 32367 15697
rect 32309 15657 32321 15691
rect 32355 15688 32367 15691
rect 32950 15688 32956 15700
rect 32355 15660 32956 15688
rect 32355 15657 32367 15660
rect 32309 15651 32367 15657
rect 32950 15648 32956 15660
rect 33008 15648 33014 15700
rect 1581 15487 1639 15493
rect 1581 15453 1593 15487
rect 1627 15484 1639 15487
rect 2958 15484 2964 15496
rect 1627 15456 2964 15484
rect 1627 15453 1639 15456
rect 1581 15447 1639 15453
rect 2958 15444 2964 15456
rect 3016 15444 3022 15496
rect 32125 15419 32183 15425
rect 32125 15385 32137 15419
rect 32171 15416 32183 15419
rect 32674 15416 32680 15428
rect 32171 15388 32680 15416
rect 32171 15385 32183 15388
rect 32125 15379 32183 15385
rect 32674 15376 32680 15388
rect 32732 15376 32738 15428
rect 934 15308 940 15360
rect 992 15348 998 15360
rect 1765 15351 1823 15357
rect 1765 15348 1777 15351
rect 992 15320 1777 15348
rect 992 15308 998 15320
rect 1765 15317 1777 15320
rect 1811 15317 1823 15351
rect 1765 15311 1823 15317
rect 31754 15308 31760 15360
rect 31812 15348 31818 15360
rect 32325 15351 32383 15357
rect 32325 15348 32337 15351
rect 31812 15320 32337 15348
rect 31812 15308 31818 15320
rect 32325 15317 32337 15320
rect 32371 15317 32383 15351
rect 32325 15311 32383 15317
rect 32490 15308 32496 15360
rect 32548 15308 32554 15360
rect 1104 15258 45051 15280
rect 1104 15206 11896 15258
rect 11948 15206 11960 15258
rect 12012 15206 12024 15258
rect 12076 15206 12088 15258
rect 12140 15206 12152 15258
rect 12204 15206 22843 15258
rect 22895 15206 22907 15258
rect 22959 15206 22971 15258
rect 23023 15206 23035 15258
rect 23087 15206 23099 15258
rect 23151 15206 33790 15258
rect 33842 15206 33854 15258
rect 33906 15206 33918 15258
rect 33970 15206 33982 15258
rect 34034 15206 34046 15258
rect 34098 15206 44737 15258
rect 44789 15206 44801 15258
rect 44853 15206 44865 15258
rect 44917 15206 44929 15258
rect 44981 15206 44993 15258
rect 45045 15206 45051 15258
rect 1104 15184 45051 15206
rect 23290 15104 23296 15156
rect 23348 15104 23354 15156
rect 26329 15147 26387 15153
rect 26329 15113 26341 15147
rect 26375 15144 26387 15147
rect 34882 15144 34888 15156
rect 26375 15116 34888 15144
rect 26375 15113 26387 15116
rect 26329 15107 26387 15113
rect 34882 15104 34888 15116
rect 34940 15104 34946 15156
rect 18874 15036 18880 15088
rect 18932 15036 18938 15088
rect 26234 15036 26240 15088
rect 26292 15076 26298 15088
rect 32214 15076 32220 15088
rect 26292 15048 32220 15076
rect 26292 15036 26298 15048
rect 32214 15036 32220 15048
rect 32272 15036 32278 15088
rect 32585 15079 32643 15085
rect 32585 15045 32597 15079
rect 32631 15076 32643 15079
rect 33502 15076 33508 15088
rect 32631 15048 33508 15076
rect 32631 15045 32643 15048
rect 32585 15039 32643 15045
rect 33502 15036 33508 15048
rect 33560 15076 33566 15088
rect 33560 15048 33916 15076
rect 33560 15036 33566 15048
rect 23201 15011 23259 15017
rect 23201 14977 23213 15011
rect 23247 14977 23259 15011
rect 23201 14971 23259 14977
rect 31481 15011 31539 15017
rect 31481 14977 31493 15011
rect 31527 15008 31539 15011
rect 32490 15008 32496 15020
rect 31527 14980 32496 15008
rect 31527 14977 31539 14980
rect 31481 14971 31539 14977
rect 18138 14900 18144 14952
rect 18196 14900 18202 14952
rect 18417 14943 18475 14949
rect 18417 14909 18429 14943
rect 18463 14940 18475 14943
rect 20070 14940 20076 14952
rect 18463 14912 20076 14940
rect 18463 14909 18475 14912
rect 18417 14903 18475 14909
rect 20070 14900 20076 14912
rect 20128 14900 20134 14952
rect 23216 14872 23244 14971
rect 32490 14968 32496 14980
rect 32548 15008 32554 15020
rect 32548 14980 33180 15008
rect 32548 14968 32554 14980
rect 23385 14943 23443 14949
rect 23385 14909 23397 14943
rect 23431 14940 23443 14943
rect 26513 14943 26571 14949
rect 26513 14940 26525 14943
rect 23431 14912 26525 14940
rect 23431 14909 23443 14912
rect 23385 14903 23443 14909
rect 26513 14909 26525 14912
rect 26559 14940 26571 14943
rect 26602 14940 26608 14952
rect 26559 14912 26608 14940
rect 26559 14909 26571 14912
rect 26513 14903 26571 14909
rect 26602 14900 26608 14912
rect 26660 14900 26666 14952
rect 31757 14943 31815 14949
rect 30760 14912 31708 14940
rect 30760 14872 30788 14912
rect 19444 14844 30788 14872
rect 18414 14764 18420 14816
rect 18472 14804 18478 14816
rect 19444 14804 19472 14844
rect 31570 14832 31576 14884
rect 31628 14832 31634 14884
rect 31680 14872 31708 14912
rect 31757 14909 31769 14943
rect 31803 14940 31815 14943
rect 31846 14940 31852 14952
rect 31803 14912 31852 14940
rect 31803 14909 31815 14912
rect 31757 14903 31815 14909
rect 31846 14900 31852 14912
rect 31904 14900 31910 14952
rect 32306 14900 32312 14952
rect 32364 14900 32370 14952
rect 32674 14900 32680 14952
rect 32732 14900 32738 14952
rect 32794 14943 32852 14949
rect 32794 14909 32806 14943
rect 32840 14940 32852 14943
rect 32950 14940 32956 14952
rect 32840 14912 32956 14940
rect 32840 14909 32852 14912
rect 32794 14903 32852 14909
rect 32950 14900 32956 14912
rect 33008 14900 33014 14952
rect 33152 14940 33180 14980
rect 33594 14968 33600 15020
rect 33652 14968 33658 15020
rect 33888 15017 33916 15048
rect 33962 15036 33968 15088
rect 34020 15076 34026 15088
rect 37826 15076 37832 15088
rect 34020 15048 37832 15076
rect 34020 15036 34026 15048
rect 37826 15036 37832 15048
rect 37884 15036 37890 15088
rect 33873 15011 33931 15017
rect 33873 14977 33885 15011
rect 33919 15008 33931 15011
rect 34333 15011 34391 15017
rect 34333 15008 34345 15011
rect 33919 14980 34345 15008
rect 33919 14977 33931 14980
rect 33873 14971 33931 14977
rect 34333 14977 34345 14980
rect 34379 14977 34391 15011
rect 34333 14971 34391 14977
rect 34517 15011 34575 15017
rect 34517 14977 34529 15011
rect 34563 14977 34575 15011
rect 36357 15011 36415 15017
rect 36357 15008 36369 15011
rect 34517 14971 34575 14977
rect 34900 14980 36369 15008
rect 33781 14943 33839 14949
rect 33781 14940 33793 14943
rect 33152 14912 33793 14940
rect 33781 14909 33793 14912
rect 33827 14940 33839 14943
rect 34532 14940 34560 14971
rect 33827 14912 34560 14940
rect 33827 14909 33839 14912
rect 33781 14903 33839 14909
rect 32582 14872 32588 14884
rect 31680 14844 32588 14872
rect 32582 14832 32588 14844
rect 32640 14832 32646 14884
rect 34514 14872 34520 14884
rect 32692 14844 34520 14872
rect 18472 14776 19472 14804
rect 19889 14807 19947 14813
rect 18472 14764 18478 14776
rect 19889 14773 19901 14807
rect 19935 14804 19947 14807
rect 20438 14804 20444 14816
rect 19935 14776 20444 14804
rect 19935 14773 19947 14776
rect 19889 14767 19947 14773
rect 20438 14764 20444 14776
rect 20496 14764 20502 14816
rect 22830 14764 22836 14816
rect 22888 14764 22894 14816
rect 25130 14764 25136 14816
rect 25188 14804 25194 14816
rect 25869 14807 25927 14813
rect 25869 14804 25881 14807
rect 25188 14776 25881 14804
rect 25188 14764 25194 14776
rect 25869 14773 25881 14776
rect 25915 14773 25927 14807
rect 25869 14767 25927 14773
rect 31386 14764 31392 14816
rect 31444 14804 31450 14816
rect 31481 14807 31539 14813
rect 31481 14804 31493 14807
rect 31444 14776 31493 14804
rect 31444 14764 31450 14776
rect 31481 14773 31493 14776
rect 31527 14773 31539 14807
rect 31481 14767 31539 14773
rect 32214 14764 32220 14816
rect 32272 14804 32278 14816
rect 32692 14804 32720 14844
rect 34514 14832 34520 14844
rect 34572 14832 34578 14884
rect 34900 14816 34928 14980
rect 36357 14977 36369 14980
rect 36403 14977 36415 15011
rect 36357 14971 36415 14977
rect 36538 14968 36544 15020
rect 36596 14968 36602 15020
rect 36906 14968 36912 15020
rect 36964 15008 36970 15020
rect 37645 15011 37703 15017
rect 37645 15008 37657 15011
rect 36964 14980 37657 15008
rect 36964 14968 36970 14980
rect 37645 14977 37657 14980
rect 37691 14977 37703 15011
rect 37645 14971 37703 14977
rect 32272 14776 32720 14804
rect 32272 14764 32278 14776
rect 32766 14764 32772 14816
rect 32824 14804 32830 14816
rect 32953 14807 33011 14813
rect 32953 14804 32965 14807
rect 32824 14776 32965 14804
rect 32824 14764 32830 14776
rect 32953 14773 32965 14776
rect 32999 14773 33011 14807
rect 32953 14767 33011 14773
rect 33410 14764 33416 14816
rect 33468 14764 33474 14816
rect 34701 14807 34759 14813
rect 34701 14773 34713 14807
rect 34747 14804 34759 14807
rect 34882 14804 34888 14816
rect 34747 14776 34888 14804
rect 34747 14773 34759 14776
rect 34701 14767 34759 14773
rect 34882 14764 34888 14776
rect 34940 14764 34946 14816
rect 36449 14807 36507 14813
rect 36449 14773 36461 14807
rect 36495 14804 36507 14807
rect 36630 14804 36636 14816
rect 36495 14776 36636 14804
rect 36495 14773 36507 14776
rect 36449 14767 36507 14773
rect 36630 14764 36636 14776
rect 36688 14764 36694 14816
rect 37458 14764 37464 14816
rect 37516 14764 37522 14816
rect 37826 14764 37832 14816
rect 37884 14804 37890 14816
rect 38930 14804 38936 14816
rect 37884 14776 38936 14804
rect 37884 14764 37890 14776
rect 38930 14764 38936 14776
rect 38988 14764 38994 14816
rect 1104 14714 44896 14736
rect 1104 14662 6423 14714
rect 6475 14662 6487 14714
rect 6539 14662 6551 14714
rect 6603 14662 6615 14714
rect 6667 14662 6679 14714
rect 6731 14662 17370 14714
rect 17422 14662 17434 14714
rect 17486 14662 17498 14714
rect 17550 14662 17562 14714
rect 17614 14662 17626 14714
rect 17678 14662 28317 14714
rect 28369 14662 28381 14714
rect 28433 14662 28445 14714
rect 28497 14662 28509 14714
rect 28561 14662 28573 14714
rect 28625 14662 39264 14714
rect 39316 14662 39328 14714
rect 39380 14662 39392 14714
rect 39444 14662 39456 14714
rect 39508 14662 39520 14714
rect 39572 14662 44896 14714
rect 1104 14640 44896 14662
rect 1946 14560 1952 14612
rect 2004 14600 2010 14612
rect 27246 14600 27252 14612
rect 2004 14572 22094 14600
rect 2004 14560 2010 14572
rect 18785 14535 18843 14541
rect 18785 14501 18797 14535
rect 18831 14532 18843 14535
rect 18874 14532 18880 14544
rect 18831 14504 18880 14532
rect 18831 14501 18843 14504
rect 18785 14495 18843 14501
rect 18874 14492 18880 14504
rect 18932 14492 18938 14544
rect 18138 14424 18144 14476
rect 18196 14464 18202 14476
rect 22066 14464 22094 14572
rect 22756 14572 27252 14600
rect 22756 14473 22784 14572
rect 27246 14560 27252 14572
rect 27304 14560 27310 14612
rect 30282 14560 30288 14612
rect 30340 14600 30346 14612
rect 30340 14572 32628 14600
rect 30340 14560 30346 14572
rect 32600 14532 32628 14572
rect 32674 14560 32680 14612
rect 32732 14600 32738 14612
rect 33229 14603 33287 14609
rect 33229 14600 33241 14603
rect 32732 14572 33241 14600
rect 32732 14560 32738 14572
rect 33229 14569 33241 14572
rect 33275 14569 33287 14603
rect 33229 14563 33287 14569
rect 33594 14560 33600 14612
rect 33652 14600 33658 14612
rect 34885 14603 34943 14609
rect 34885 14600 34897 14603
rect 33652 14572 34897 14600
rect 33652 14560 33658 14572
rect 34885 14569 34897 14572
rect 34931 14569 34943 14603
rect 34885 14563 34943 14569
rect 41325 14603 41383 14609
rect 41325 14569 41337 14603
rect 41371 14600 41383 14603
rect 42702 14600 42708 14612
rect 41371 14572 42708 14600
rect 41371 14569 41383 14572
rect 41325 14563 41383 14569
rect 42702 14560 42708 14572
rect 42760 14560 42766 14612
rect 36446 14532 36452 14544
rect 32600 14504 36452 14532
rect 36446 14492 36452 14504
rect 36504 14492 36510 14544
rect 42797 14535 42855 14541
rect 42797 14501 42809 14535
rect 42843 14501 42855 14535
rect 42797 14495 42855 14501
rect 22741 14467 22799 14473
rect 22741 14464 22753 14467
rect 18196 14436 20392 14464
rect 22066 14436 22753 14464
rect 18196 14424 18202 14436
rect 9858 14356 9864 14408
rect 9916 14356 9922 14408
rect 9950 14356 9956 14408
rect 10008 14396 10014 14408
rect 10117 14399 10175 14405
rect 10117 14396 10129 14399
rect 10008 14368 10129 14396
rect 10008 14356 10014 14368
rect 10117 14365 10129 14368
rect 10163 14365 10175 14399
rect 10117 14359 10175 14365
rect 18233 14399 18291 14405
rect 18233 14365 18245 14399
rect 18279 14365 18291 14399
rect 18233 14359 18291 14365
rect 13354 14288 13360 14340
rect 13412 14328 13418 14340
rect 18248 14328 18276 14359
rect 18690 14356 18696 14408
rect 18748 14396 18754 14408
rect 20364 14405 20392 14436
rect 22741 14433 22753 14436
rect 22787 14433 22799 14467
rect 22741 14427 22799 14433
rect 32950 14424 32956 14476
rect 33008 14464 33014 14476
rect 42812 14464 42840 14495
rect 33008 14436 33364 14464
rect 42812 14436 44128 14464
rect 33008 14424 33014 14436
rect 19429 14399 19487 14405
rect 19429 14396 19441 14399
rect 18748 14368 19441 14396
rect 18748 14356 18754 14368
rect 19429 14365 19441 14368
rect 19475 14365 19487 14399
rect 19429 14359 19487 14365
rect 20349 14399 20407 14405
rect 20349 14365 20361 14399
rect 20395 14396 20407 14399
rect 22554 14396 22560 14408
rect 20395 14368 22560 14396
rect 20395 14365 20407 14368
rect 20349 14359 20407 14365
rect 22554 14356 22560 14368
rect 22612 14356 22618 14408
rect 26145 14399 26203 14405
rect 26145 14365 26157 14399
rect 26191 14396 26203 14399
rect 26191 14368 26556 14396
rect 26191 14365 26203 14368
rect 26145 14359 26203 14365
rect 26528 14340 26556 14368
rect 29178 14356 29184 14408
rect 29236 14396 29242 14408
rect 31297 14399 31355 14405
rect 31297 14396 31309 14399
rect 29236 14368 31309 14396
rect 29236 14356 29242 14368
rect 31297 14365 31309 14368
rect 31343 14365 31355 14399
rect 31297 14359 31355 14365
rect 31386 14356 31392 14408
rect 31444 14396 31450 14408
rect 31553 14399 31611 14405
rect 31553 14396 31565 14399
rect 31444 14368 31565 14396
rect 31444 14356 31450 14368
rect 31553 14365 31565 14368
rect 31599 14365 31611 14399
rect 33336 14396 33364 14436
rect 33413 14399 33471 14405
rect 33413 14396 33425 14399
rect 33336 14368 33425 14396
rect 31553 14359 31611 14365
rect 33413 14365 33425 14368
rect 33459 14365 33471 14399
rect 33413 14359 33471 14365
rect 33502 14356 33508 14408
rect 33560 14396 33566 14408
rect 33597 14399 33655 14405
rect 33597 14396 33609 14399
rect 33560 14368 33609 14396
rect 33560 14356 33566 14368
rect 33597 14365 33609 14368
rect 33643 14365 33655 14399
rect 33597 14359 33655 14365
rect 34882 14356 34888 14408
rect 34940 14356 34946 14408
rect 35069 14399 35127 14405
rect 35069 14365 35081 14399
rect 35115 14396 35127 14399
rect 35158 14396 35164 14408
rect 35115 14368 35164 14396
rect 35115 14365 35127 14368
rect 35069 14359 35127 14365
rect 35158 14356 35164 14368
rect 35216 14356 35222 14408
rect 36814 14356 36820 14408
rect 36872 14356 36878 14408
rect 37084 14399 37142 14405
rect 37084 14365 37096 14399
rect 37130 14396 37142 14399
rect 37458 14396 37464 14408
rect 37130 14368 37464 14396
rect 37130 14365 37142 14368
rect 37084 14359 37142 14365
rect 37458 14356 37464 14368
rect 37516 14356 37522 14408
rect 40954 14356 40960 14408
rect 41012 14356 41018 14408
rect 42153 14399 42211 14405
rect 42153 14396 42165 14399
rect 41524 14368 42165 14396
rect 20162 14328 20168 14340
rect 13412 14300 18184 14328
rect 18248 14300 20168 14328
rect 13412 14288 13418 14300
rect 11238 14220 11244 14272
rect 11296 14220 11302 14272
rect 11330 14220 11336 14272
rect 11388 14260 11394 14272
rect 14366 14260 14372 14272
rect 11388 14232 14372 14260
rect 11388 14220 11394 14232
rect 14366 14220 14372 14232
rect 14424 14220 14430 14272
rect 18046 14220 18052 14272
rect 18104 14220 18110 14272
rect 18156 14260 18184 14300
rect 20162 14288 20168 14300
rect 20220 14288 20226 14340
rect 20254 14288 20260 14340
rect 20312 14328 20318 14340
rect 26418 14337 26424 14340
rect 20594 14331 20652 14337
rect 20594 14328 20606 14331
rect 20312 14300 20606 14328
rect 20312 14288 20318 14300
rect 20594 14297 20606 14300
rect 20640 14297 20652 14331
rect 22649 14331 22707 14337
rect 22649 14328 22661 14331
rect 20594 14291 20652 14297
rect 22066 14300 22661 14328
rect 18414 14260 18420 14272
rect 18156 14232 18420 14260
rect 18414 14220 18420 14232
rect 18472 14220 18478 14272
rect 19518 14220 19524 14272
rect 19576 14220 19582 14272
rect 21729 14263 21787 14269
rect 21729 14229 21741 14263
rect 21775 14260 21787 14263
rect 22066 14260 22094 14300
rect 22649 14297 22661 14300
rect 22695 14297 22707 14331
rect 22649 14291 22707 14297
rect 26412 14291 26424 14337
rect 26418 14288 26424 14291
rect 26476 14288 26482 14340
rect 26510 14288 26516 14340
rect 26568 14288 26574 14340
rect 32306 14288 32312 14340
rect 32364 14328 32370 14340
rect 33137 14331 33195 14337
rect 33137 14328 33149 14331
rect 32364 14300 33149 14328
rect 32364 14288 32370 14300
rect 33137 14297 33149 14300
rect 33183 14328 33195 14331
rect 34900 14328 34928 14356
rect 35989 14331 36047 14337
rect 35989 14328 36001 14331
rect 33183 14300 34836 14328
rect 34900 14300 36001 14328
rect 33183 14297 33195 14300
rect 33137 14291 33195 14297
rect 21775 14232 22094 14260
rect 22189 14263 22247 14269
rect 21775 14229 21787 14232
rect 21729 14223 21787 14229
rect 22189 14229 22201 14263
rect 22235 14260 22247 14263
rect 22370 14260 22376 14272
rect 22235 14232 22376 14260
rect 22235 14229 22247 14232
rect 22189 14223 22247 14229
rect 22370 14220 22376 14232
rect 22428 14220 22434 14272
rect 22557 14263 22615 14269
rect 22557 14229 22569 14263
rect 22603 14260 22615 14263
rect 22830 14260 22836 14272
rect 22603 14232 22836 14260
rect 22603 14229 22615 14232
rect 22557 14223 22615 14229
rect 22830 14220 22836 14232
rect 22888 14220 22894 14272
rect 27522 14220 27528 14272
rect 27580 14220 27586 14272
rect 32674 14220 32680 14272
rect 32732 14220 32738 14272
rect 33226 14220 33232 14272
rect 33284 14260 33290 14272
rect 33781 14263 33839 14269
rect 33781 14260 33793 14263
rect 33284 14232 33793 14260
rect 33284 14220 33290 14232
rect 33781 14229 33793 14232
rect 33827 14229 33839 14263
rect 34808 14260 34836 14300
rect 35989 14297 36001 14300
rect 36035 14297 36047 14331
rect 35989 14291 36047 14297
rect 36173 14331 36231 14337
rect 36173 14297 36185 14331
rect 36219 14328 36231 14331
rect 36538 14328 36544 14340
rect 36219 14300 36544 14328
rect 36219 14297 36231 14300
rect 36173 14291 36231 14297
rect 36188 14260 36216 14291
rect 36538 14288 36544 14300
rect 36596 14288 36602 14340
rect 34808 14232 36216 14260
rect 33781 14223 33839 14229
rect 36354 14220 36360 14272
rect 36412 14220 36418 14272
rect 36556 14260 36584 14288
rect 38197 14263 38255 14269
rect 38197 14260 38209 14263
rect 36556 14232 38209 14260
rect 38197 14229 38209 14232
rect 38243 14229 38255 14263
rect 38197 14223 38255 14229
rect 40494 14220 40500 14272
rect 40552 14260 40558 14272
rect 41524 14269 41552 14368
rect 42153 14365 42165 14368
rect 42199 14365 42211 14399
rect 42153 14359 42211 14365
rect 42978 14356 42984 14408
rect 43036 14356 43042 14408
rect 44100 14405 44128 14436
rect 44085 14399 44143 14405
rect 44085 14365 44097 14399
rect 44131 14365 44143 14399
rect 44085 14359 44143 14365
rect 41325 14263 41383 14269
rect 41325 14260 41337 14263
rect 40552 14232 41337 14260
rect 40552 14220 40558 14232
rect 41325 14229 41337 14232
rect 41371 14229 41383 14263
rect 41325 14223 41383 14229
rect 41509 14263 41567 14269
rect 41509 14229 41521 14263
rect 41555 14229 41567 14263
rect 41509 14223 41567 14229
rect 41966 14220 41972 14272
rect 42024 14220 42030 14272
rect 44266 14220 44272 14272
rect 44324 14220 44330 14272
rect 1104 14170 45051 14192
rect 1104 14118 11896 14170
rect 11948 14118 11960 14170
rect 12012 14118 12024 14170
rect 12076 14118 12088 14170
rect 12140 14118 12152 14170
rect 12204 14118 22843 14170
rect 22895 14118 22907 14170
rect 22959 14118 22971 14170
rect 23023 14118 23035 14170
rect 23087 14118 23099 14170
rect 23151 14118 33790 14170
rect 33842 14118 33854 14170
rect 33906 14118 33918 14170
rect 33970 14118 33982 14170
rect 34034 14118 34046 14170
rect 34098 14118 44737 14170
rect 44789 14118 44801 14170
rect 44853 14118 44865 14170
rect 44917 14118 44929 14170
rect 44981 14118 44993 14170
rect 45045 14118 45051 14170
rect 1104 14096 45051 14118
rect 6631 14059 6689 14065
rect 6631 14025 6643 14059
rect 6677 14056 6689 14059
rect 6822 14056 6828 14068
rect 6677 14028 6828 14056
rect 6677 14025 6689 14028
rect 6631 14019 6689 14025
rect 6822 14016 6828 14028
rect 6880 14016 6886 14068
rect 16298 14056 16304 14068
rect 12360 14028 16304 14056
rect 5534 13948 5540 14000
rect 5592 13988 5598 14000
rect 7101 13991 7159 13997
rect 7101 13988 7113 13991
rect 5592 13960 7113 13988
rect 5592 13948 5598 13960
rect 7101 13957 7113 13960
rect 7147 13957 7159 13991
rect 7101 13951 7159 13957
rect 5350 13880 5356 13932
rect 5408 13880 5414 13932
rect 6914 13880 6920 13932
rect 6972 13920 6978 13932
rect 12360 13920 12388 14028
rect 16298 14016 16304 14028
rect 16356 14016 16362 14068
rect 17313 14059 17371 14065
rect 17313 14025 17325 14059
rect 17359 14056 17371 14059
rect 17954 14056 17960 14068
rect 17359 14028 17960 14056
rect 17359 14025 17371 14028
rect 17313 14019 17371 14025
rect 17954 14016 17960 14028
rect 18012 14016 18018 14068
rect 20070 14016 20076 14068
rect 20128 14016 20134 14068
rect 20162 14016 20168 14068
rect 20220 14056 20226 14068
rect 21361 14059 21419 14065
rect 21361 14056 21373 14059
rect 20220 14028 21373 14056
rect 20220 14016 20226 14028
rect 21361 14025 21373 14028
rect 21407 14025 21419 14059
rect 21361 14019 21419 14025
rect 22281 14059 22339 14065
rect 22281 14025 22293 14059
rect 22327 14025 22339 14059
rect 22281 14019 22339 14025
rect 24305 14059 24363 14065
rect 24305 14025 24317 14059
rect 24351 14025 24363 14059
rect 24305 14019 24363 14025
rect 14642 13988 14648 14000
rect 12636 13960 14648 13988
rect 12636 13929 12664 13960
rect 14642 13948 14648 13960
rect 14700 13948 14706 14000
rect 18138 13988 18144 14000
rect 17880 13960 18144 13988
rect 13354 13929 13360 13932
rect 6972 13892 12388 13920
rect 12621 13923 12679 13929
rect 6972 13880 6978 13892
rect 12621 13889 12633 13923
rect 12667 13889 12679 13923
rect 13348 13920 13360 13929
rect 13315 13892 13360 13920
rect 12621 13883 12679 13889
rect 13348 13883 13360 13892
rect 13354 13880 13360 13883
rect 13412 13880 13418 13932
rect 17218 13880 17224 13932
rect 17276 13880 17282 13932
rect 17880 13929 17908 13960
rect 18138 13948 18144 13960
rect 18196 13948 18202 14000
rect 19518 13988 19524 14000
rect 19366 13960 19524 13988
rect 19518 13948 19524 13960
rect 19576 13948 19582 14000
rect 20438 13948 20444 14000
rect 20496 13948 20502 14000
rect 22296 13988 22324 14019
rect 23170 13991 23228 13997
rect 23170 13988 23182 13991
rect 22296 13960 23182 13988
rect 23170 13957 23182 13960
rect 23216 13957 23228 13991
rect 24320 13988 24348 14019
rect 25130 14016 25136 14068
rect 25188 14016 25194 14068
rect 27430 14056 27436 14068
rect 25332 14028 27436 14056
rect 25225 13991 25283 13997
rect 25225 13988 25237 13991
rect 24320 13960 25237 13988
rect 23170 13951 23228 13957
rect 25225 13957 25237 13960
rect 25271 13957 25283 13991
rect 25225 13951 25283 13957
rect 17865 13923 17923 13929
rect 17865 13889 17877 13923
rect 17911 13889 17923 13923
rect 17865 13883 17923 13889
rect 20254 13880 20260 13932
rect 20312 13880 20318 13932
rect 20533 13923 20591 13929
rect 20533 13889 20545 13923
rect 20579 13920 20591 13923
rect 20622 13920 20628 13932
rect 20579 13892 20628 13920
rect 20579 13889 20591 13892
rect 20533 13883 20591 13889
rect 20622 13880 20628 13892
rect 20680 13880 20686 13932
rect 21174 13880 21180 13932
rect 21232 13880 21238 13932
rect 22462 13880 22468 13932
rect 22520 13880 22526 13932
rect 22554 13880 22560 13932
rect 22612 13920 22618 13932
rect 22925 13923 22983 13929
rect 22925 13920 22937 13923
rect 22612 13892 22937 13920
rect 22612 13880 22618 13892
rect 22925 13889 22937 13892
rect 22971 13889 22983 13923
rect 25332 13920 25360 14028
rect 27430 14016 27436 14028
rect 27488 14016 27494 14068
rect 27522 14016 27528 14068
rect 27580 14056 27586 14068
rect 27617 14059 27675 14065
rect 27617 14056 27629 14059
rect 27580 14028 27629 14056
rect 27580 14016 27586 14028
rect 27617 14025 27629 14028
rect 27663 14025 27675 14059
rect 27617 14019 27675 14025
rect 31570 14016 31576 14068
rect 31628 14065 31634 14068
rect 31628 14056 31637 14065
rect 31628 14028 31673 14056
rect 31628 14019 31637 14028
rect 31628 14016 31634 14019
rect 33502 14016 33508 14068
rect 33560 14056 33566 14068
rect 34241 14059 34299 14065
rect 34241 14056 34253 14059
rect 33560 14028 34253 14056
rect 33560 14016 33566 14028
rect 34241 14025 34253 14028
rect 34287 14025 34299 14059
rect 34241 14019 34299 14025
rect 34790 14016 34796 14068
rect 34848 14056 34854 14068
rect 36262 14056 36268 14068
rect 34848 14028 36268 14056
rect 34848 14016 34854 14028
rect 36262 14016 36268 14028
rect 36320 14016 36326 14068
rect 36446 14016 36452 14068
rect 36504 14056 36510 14068
rect 36541 14059 36599 14065
rect 36541 14056 36553 14059
rect 36504 14028 36553 14056
rect 36504 14016 36510 14028
rect 36541 14025 36553 14028
rect 36587 14025 36599 14059
rect 36541 14019 36599 14025
rect 36630 14016 36636 14068
rect 36688 14016 36694 14068
rect 36906 14016 36912 14068
rect 36964 14016 36970 14068
rect 37274 14016 37280 14068
rect 37332 14056 37338 14068
rect 37332 14028 38240 14056
rect 37332 14016 37338 14028
rect 26053 13991 26111 13997
rect 26053 13957 26065 13991
rect 26099 13988 26111 13991
rect 26099 13960 26464 13988
rect 26099 13957 26111 13960
rect 26053 13951 26111 13957
rect 22925 13883 22983 13889
rect 23032 13892 25360 13920
rect 934 13812 940 13864
rect 992 13852 998 13864
rect 1765 13855 1823 13861
rect 1765 13852 1777 13855
rect 992 13824 1777 13852
rect 992 13812 998 13824
rect 1765 13821 1777 13824
rect 1811 13821 1823 13855
rect 1765 13815 1823 13821
rect 5169 13855 5227 13861
rect 5169 13821 5181 13855
rect 5215 13852 5227 13855
rect 7193 13855 7251 13861
rect 7193 13852 7205 13855
rect 5215 13824 7205 13852
rect 5215 13821 5227 13824
rect 5169 13815 5227 13821
rect 7193 13821 7205 13824
rect 7239 13852 7251 13855
rect 11330 13852 11336 13864
rect 7239 13824 11336 13852
rect 7239 13821 7251 13824
rect 7193 13815 7251 13821
rect 11330 13812 11336 13824
rect 11388 13812 11394 13864
rect 11422 13812 11428 13864
rect 11480 13852 11486 13864
rect 13081 13855 13139 13861
rect 13081 13852 13093 13855
rect 11480 13824 13093 13852
rect 11480 13812 11486 13824
rect 13081 13821 13093 13824
rect 13127 13821 13139 13855
rect 13081 13815 13139 13821
rect 18141 13855 18199 13861
rect 18141 13821 18153 13855
rect 18187 13852 18199 13855
rect 18506 13852 18512 13864
rect 18187 13824 18512 13852
rect 18187 13821 18199 13824
rect 18141 13815 18199 13821
rect 18506 13812 18512 13824
rect 18564 13812 18570 13864
rect 20806 13812 20812 13864
rect 20864 13852 20870 13864
rect 20993 13855 21051 13861
rect 20993 13852 21005 13855
rect 20864 13824 21005 13852
rect 20864 13812 20870 13824
rect 20993 13821 21005 13824
rect 21039 13821 21051 13855
rect 20993 13815 21051 13821
rect 21266 13812 21272 13864
rect 21324 13852 21330 13864
rect 23032 13852 23060 13892
rect 25332 13861 25360 13892
rect 26237 13923 26295 13929
rect 26237 13889 26249 13923
rect 26283 13920 26295 13923
rect 26326 13920 26332 13932
rect 26283 13892 26332 13920
rect 26283 13889 26295 13892
rect 26237 13883 26295 13889
rect 26326 13880 26332 13892
rect 26384 13880 26390 13932
rect 26436 13920 26464 13960
rect 26510 13948 26516 14000
rect 26568 13988 26574 14000
rect 29178 13988 29184 14000
rect 26568 13960 29184 13988
rect 26568 13948 26574 13960
rect 27154 13920 27160 13932
rect 26436 13892 27160 13920
rect 27154 13880 27160 13892
rect 27212 13880 27218 13932
rect 27522 13880 27528 13932
rect 27580 13880 27586 13932
rect 28368 13929 28396 13960
rect 29178 13948 29184 13960
rect 29236 13948 29242 14000
rect 30193 13991 30251 13997
rect 30193 13957 30205 13991
rect 30239 13957 30251 13991
rect 30193 13951 30251 13957
rect 28353 13923 28411 13929
rect 28353 13889 28365 13923
rect 28399 13889 28411 13923
rect 28353 13883 28411 13889
rect 28620 13923 28678 13929
rect 28620 13889 28632 13923
rect 28666 13920 28678 13923
rect 30208 13920 30236 13951
rect 30282 13948 30288 14000
rect 30340 13988 30346 14000
rect 31481 13991 31539 13997
rect 30340 13960 30696 13988
rect 30340 13948 30346 13960
rect 28666 13892 30236 13920
rect 30469 13923 30527 13929
rect 28666 13889 28678 13892
rect 28620 13883 28678 13889
rect 30469 13889 30481 13923
rect 30515 13889 30527 13923
rect 30469 13883 30527 13889
rect 21324 13824 23060 13852
rect 25317 13855 25375 13861
rect 21324 13812 21330 13824
rect 25317 13821 25329 13855
rect 25363 13821 25375 13855
rect 27614 13852 27620 13864
rect 25317 13815 25375 13821
rect 27172 13824 27620 13852
rect 1854 13744 1860 13796
rect 1912 13784 1918 13796
rect 27172 13793 27200 13824
rect 27614 13812 27620 13824
rect 27672 13812 27678 13864
rect 27709 13855 27767 13861
rect 27709 13821 27721 13855
rect 27755 13821 27767 13855
rect 27709 13815 27767 13821
rect 27157 13787 27215 13793
rect 1912 13756 13124 13784
rect 1912 13744 1918 13756
rect 5537 13719 5595 13725
rect 5537 13685 5549 13719
rect 5583 13716 5595 13719
rect 5626 13716 5632 13728
rect 5583 13688 5632 13716
rect 5583 13685 5595 13688
rect 5537 13679 5595 13685
rect 5626 13676 5632 13688
rect 5684 13676 5690 13728
rect 12434 13676 12440 13728
rect 12492 13676 12498 13728
rect 13096 13716 13124 13756
rect 14016 13756 17448 13784
rect 14016 13716 14044 13756
rect 13096 13688 14044 13716
rect 14458 13676 14464 13728
rect 14516 13676 14522 13728
rect 17420 13716 17448 13756
rect 19168 13756 22416 13784
rect 19168 13716 19196 13756
rect 17420 13688 19196 13716
rect 19613 13719 19671 13725
rect 19613 13685 19625 13719
rect 19659 13716 19671 13719
rect 19978 13716 19984 13728
rect 19659 13688 19984 13716
rect 19659 13685 19671 13688
rect 19613 13679 19671 13685
rect 19978 13676 19984 13688
rect 20036 13676 20042 13728
rect 22388 13716 22416 13756
rect 23860 13756 27108 13784
rect 23860 13716 23888 13756
rect 22388 13688 23888 13716
rect 24762 13676 24768 13728
rect 24820 13676 24826 13728
rect 26421 13719 26479 13725
rect 26421 13685 26433 13719
rect 26467 13716 26479 13719
rect 26970 13716 26976 13728
rect 26467 13688 26976 13716
rect 26467 13685 26479 13688
rect 26421 13679 26479 13685
rect 26970 13676 26976 13688
rect 27028 13676 27034 13728
rect 27080 13716 27108 13756
rect 27157 13753 27169 13787
rect 27203 13753 27215 13787
rect 27157 13747 27215 13753
rect 27430 13744 27436 13796
rect 27488 13784 27494 13796
rect 27724 13784 27752 13815
rect 29914 13812 29920 13864
rect 29972 13852 29978 13864
rect 30484 13852 30512 13883
rect 30558 13880 30564 13932
rect 30616 13880 30622 13932
rect 30668 13929 30696 13960
rect 31481 13957 31493 13991
rect 31527 13988 31539 13991
rect 32674 13988 32680 14000
rect 31527 13960 32680 13988
rect 31527 13957 31539 13960
rect 31481 13951 31539 13957
rect 32674 13948 32680 13960
rect 32732 13948 32738 14000
rect 33686 13988 33692 14000
rect 32876 13960 33692 13988
rect 30653 13923 30711 13929
rect 30653 13889 30665 13923
rect 30699 13889 30711 13923
rect 30653 13883 30711 13889
rect 30834 13880 30840 13932
rect 30892 13880 30898 13932
rect 31665 13923 31723 13929
rect 31665 13889 31677 13923
rect 31711 13889 31723 13923
rect 31665 13883 31723 13889
rect 31680 13852 31708 13883
rect 31754 13880 31760 13932
rect 31812 13880 31818 13932
rect 32876 13929 32904 13960
rect 33686 13948 33692 13960
rect 33744 13948 33750 14000
rect 34440 13960 35480 13988
rect 32861 13923 32919 13929
rect 32861 13889 32873 13923
rect 32907 13889 32919 13923
rect 32861 13883 32919 13889
rect 32950 13880 32956 13932
rect 33008 13880 33014 13932
rect 33128 13923 33186 13929
rect 33128 13889 33140 13923
rect 33174 13920 33186 13923
rect 33410 13920 33416 13932
rect 33174 13892 33416 13920
rect 33174 13889 33186 13892
rect 33128 13883 33186 13889
rect 33410 13880 33416 13892
rect 33468 13880 33474 13932
rect 32968 13852 32996 13880
rect 29972 13824 32996 13852
rect 29972 13812 29978 13824
rect 31754 13784 31760 13796
rect 27488 13756 27752 13784
rect 29656 13756 31760 13784
rect 27488 13744 27494 13756
rect 29656 13716 29684 13756
rect 31754 13744 31760 13756
rect 31812 13744 31818 13796
rect 27080 13688 29684 13716
rect 29733 13719 29791 13725
rect 29733 13685 29745 13719
rect 29779 13716 29791 13719
rect 29914 13716 29920 13728
rect 29779 13688 29920 13716
rect 29779 13685 29791 13688
rect 29733 13679 29791 13685
rect 29914 13676 29920 13688
rect 29972 13676 29978 13728
rect 32674 13676 32680 13728
rect 32732 13716 32738 13728
rect 34440 13716 34468 13960
rect 35452 13932 35480 13960
rect 36354 13948 36360 14000
rect 36412 13988 36418 14000
rect 36750 13991 36808 13997
rect 36750 13988 36762 13991
rect 36412 13960 36762 13988
rect 36412 13948 36418 13960
rect 36750 13957 36762 13960
rect 36796 13957 36808 13991
rect 37642 13988 37648 14000
rect 36750 13951 36808 13957
rect 37108 13960 37648 13988
rect 34790 13880 34796 13932
rect 34848 13880 34854 13932
rect 34977 13923 35035 13929
rect 34977 13889 34989 13923
rect 35023 13920 35035 13923
rect 35023 13892 35388 13920
rect 35023 13889 35035 13892
rect 34977 13883 35035 13889
rect 34885 13855 34943 13861
rect 34885 13821 34897 13855
rect 34931 13852 34943 13855
rect 34931 13824 35296 13852
rect 34931 13821 34943 13824
rect 34885 13815 34943 13821
rect 32732 13688 34468 13716
rect 35268 13716 35296 13824
rect 35360 13784 35388 13892
rect 35434 13880 35440 13932
rect 35492 13880 35498 13932
rect 35529 13923 35587 13929
rect 35529 13889 35541 13923
rect 35575 13920 35587 13923
rect 37108 13920 37136 13960
rect 37642 13948 37648 13960
rect 37700 13948 37706 14000
rect 35575 13892 37136 13920
rect 37461 13923 37519 13929
rect 35575 13889 35587 13892
rect 35529 13883 35587 13889
rect 37461 13889 37473 13923
rect 37507 13920 37519 13923
rect 37550 13920 37556 13932
rect 37507 13892 37556 13920
rect 37507 13889 37519 13892
rect 37461 13883 37519 13889
rect 37550 13880 37556 13892
rect 37608 13880 37614 13932
rect 38212 13929 38240 14028
rect 40948 13991 41006 13997
rect 40948 13957 40960 13991
rect 40994 13988 41006 13991
rect 41966 13988 41972 14000
rect 40994 13960 41972 13988
rect 40994 13957 41006 13960
rect 40948 13951 41006 13957
rect 41966 13948 41972 13960
rect 42024 13948 42030 14000
rect 37737 13923 37795 13929
rect 37737 13889 37749 13923
rect 37783 13889 37795 13923
rect 37737 13883 37795 13889
rect 38197 13923 38255 13929
rect 38197 13889 38209 13923
rect 38243 13889 38255 13923
rect 38197 13883 38255 13889
rect 36265 13855 36323 13861
rect 36265 13821 36277 13855
rect 36311 13852 36323 13855
rect 36354 13852 36360 13864
rect 36311 13824 36360 13852
rect 36311 13821 36323 13824
rect 36265 13815 36323 13821
rect 36354 13812 36360 13824
rect 36412 13812 36418 13864
rect 36446 13812 36452 13864
rect 36504 13852 36510 13864
rect 37752 13852 37780 13883
rect 38378 13880 38384 13932
rect 38436 13880 38442 13932
rect 36504 13824 37780 13852
rect 38289 13855 38347 13861
rect 36504 13812 36510 13824
rect 38289 13821 38301 13855
rect 38335 13852 38347 13855
rect 38930 13852 38936 13864
rect 38335 13824 38936 13852
rect 38335 13821 38347 13824
rect 38289 13815 38347 13821
rect 38930 13812 38936 13824
rect 38988 13812 38994 13864
rect 40681 13855 40739 13861
rect 40681 13852 40693 13855
rect 40604 13824 40693 13852
rect 40604 13796 40632 13824
rect 40681 13821 40693 13824
rect 40727 13821 40739 13855
rect 40681 13815 40739 13821
rect 36078 13784 36084 13796
rect 35360 13756 36084 13784
rect 36078 13744 36084 13756
rect 36136 13744 36142 13796
rect 36814 13744 36820 13796
rect 36872 13784 36878 13796
rect 40586 13784 40592 13796
rect 36872 13756 40592 13784
rect 36872 13744 36878 13756
rect 40586 13744 40592 13756
rect 40644 13744 40650 13796
rect 36630 13716 36636 13728
rect 35268 13688 36636 13716
rect 32732 13676 32738 13688
rect 36630 13676 36636 13688
rect 36688 13676 36694 13728
rect 37458 13676 37464 13728
rect 37516 13676 37522 13728
rect 42058 13676 42064 13728
rect 42116 13676 42122 13728
rect 1104 13626 44896 13648
rect 1104 13574 6423 13626
rect 6475 13574 6487 13626
rect 6539 13574 6551 13626
rect 6603 13574 6615 13626
rect 6667 13574 6679 13626
rect 6731 13574 17370 13626
rect 17422 13574 17434 13626
rect 17486 13574 17498 13626
rect 17550 13574 17562 13626
rect 17614 13574 17626 13626
rect 17678 13574 28317 13626
rect 28369 13574 28381 13626
rect 28433 13574 28445 13626
rect 28497 13574 28509 13626
rect 28561 13574 28573 13626
rect 28625 13574 39264 13626
rect 39316 13574 39328 13626
rect 39380 13574 39392 13626
rect 39444 13574 39456 13626
rect 39508 13574 39520 13626
rect 39572 13574 44896 13626
rect 1104 13552 44896 13574
rect 14642 13472 14648 13524
rect 14700 13472 14706 13524
rect 18506 13472 18512 13524
rect 18564 13512 18570 13524
rect 19613 13515 19671 13521
rect 19613 13512 19625 13515
rect 18564 13484 19625 13512
rect 18564 13472 18570 13484
rect 19613 13481 19625 13484
rect 19659 13481 19671 13515
rect 19613 13475 19671 13481
rect 20438 13472 20444 13524
rect 20496 13512 20502 13524
rect 20533 13515 20591 13521
rect 20533 13512 20545 13515
rect 20496 13484 20545 13512
rect 20496 13472 20502 13484
rect 20533 13481 20545 13484
rect 20579 13512 20591 13515
rect 20579 13484 21128 13512
rect 20579 13481 20591 13484
rect 20533 13475 20591 13481
rect 6917 13447 6975 13453
rect 6917 13413 6929 13447
rect 6963 13444 6975 13447
rect 8570 13444 8576 13456
rect 6963 13416 8576 13444
rect 6963 13413 6975 13416
rect 6917 13407 6975 13413
rect 8570 13404 8576 13416
rect 8628 13404 8634 13456
rect 18877 13447 18935 13453
rect 18877 13413 18889 13447
rect 18923 13444 18935 13447
rect 20254 13444 20260 13456
rect 18923 13416 20260 13444
rect 18923 13413 18935 13416
rect 18877 13407 18935 13413
rect 20254 13404 20260 13416
rect 20312 13404 20318 13456
rect 21100 13444 21128 13484
rect 21174 13472 21180 13524
rect 21232 13512 21238 13524
rect 21545 13515 21603 13521
rect 21545 13512 21557 13515
rect 21232 13484 21557 13512
rect 21232 13472 21238 13484
rect 21545 13481 21557 13484
rect 21591 13512 21603 13515
rect 21591 13484 22094 13512
rect 21591 13481 21603 13484
rect 21545 13475 21603 13481
rect 22066 13444 22094 13484
rect 26326 13472 26332 13524
rect 26384 13472 26390 13524
rect 26418 13472 26424 13524
rect 26476 13512 26482 13524
rect 26789 13515 26847 13521
rect 26789 13512 26801 13515
rect 26476 13484 26801 13512
rect 26476 13472 26482 13484
rect 26789 13481 26801 13484
rect 26835 13481 26847 13515
rect 26789 13475 26847 13481
rect 29733 13515 29791 13521
rect 29733 13481 29745 13515
rect 29779 13512 29791 13515
rect 30834 13512 30840 13524
rect 29779 13484 30840 13512
rect 29779 13481 29791 13484
rect 29733 13475 29791 13481
rect 30834 13472 30840 13484
rect 30892 13472 30898 13524
rect 32122 13472 32128 13524
rect 32180 13512 32186 13524
rect 33410 13512 33416 13524
rect 32180 13484 33416 13512
rect 32180 13472 32186 13484
rect 33410 13472 33416 13484
rect 33468 13472 33474 13524
rect 35529 13515 35587 13521
rect 35529 13481 35541 13515
rect 35575 13512 35587 13515
rect 37274 13512 37280 13524
rect 35575 13484 37280 13512
rect 35575 13481 35587 13484
rect 35529 13475 35587 13481
rect 37274 13472 37280 13484
rect 37332 13472 37338 13524
rect 42702 13472 42708 13524
rect 42760 13512 42766 13524
rect 42797 13515 42855 13521
rect 42797 13512 42809 13515
rect 42760 13484 42809 13512
rect 42760 13472 42766 13484
rect 42797 13481 42809 13484
rect 42843 13481 42855 13515
rect 42797 13475 42855 13481
rect 28813 13447 28871 13453
rect 20640 13416 21036 13444
rect 21100 13416 21680 13444
rect 22066 13416 22416 13444
rect 4632 13348 5212 13376
rect 4632 13317 4660 13348
rect 4617 13311 4675 13317
rect 4617 13277 4629 13311
rect 4663 13277 4675 13311
rect 4617 13271 4675 13277
rect 5074 13268 5080 13320
rect 5132 13268 5138 13320
rect 5184 13308 5212 13348
rect 7558 13336 7564 13388
rect 7616 13376 7622 13388
rect 10873 13379 10931 13385
rect 10873 13376 10885 13379
rect 7616 13348 10885 13376
rect 7616 13336 7622 13348
rect 10873 13345 10885 13348
rect 10919 13376 10931 13379
rect 11054 13376 11060 13388
rect 10919 13348 11060 13376
rect 10919 13345 10931 13348
rect 10873 13339 10931 13345
rect 11054 13336 11060 13348
rect 11112 13336 11118 13388
rect 11422 13336 11428 13388
rect 11480 13336 11486 13388
rect 17129 13379 17187 13385
rect 17129 13345 17141 13379
rect 17175 13376 17187 13379
rect 18138 13376 18144 13388
rect 17175 13348 18144 13376
rect 17175 13345 17187 13348
rect 17129 13339 17187 13345
rect 18138 13336 18144 13348
rect 18196 13336 18202 13388
rect 20640 13376 20668 13416
rect 19996 13348 20668 13376
rect 19996 13320 20024 13348
rect 20714 13336 20720 13388
rect 20772 13336 20778 13388
rect 21008 13376 21036 13416
rect 21542 13376 21548 13388
rect 21008 13348 21548 13376
rect 5626 13308 5632 13320
rect 5184 13280 5632 13308
rect 5626 13268 5632 13280
rect 5684 13268 5690 13320
rect 11238 13268 11244 13320
rect 11296 13308 11302 13320
rect 11681 13311 11739 13317
rect 11681 13308 11693 13311
rect 11296 13280 11693 13308
rect 11296 13268 11302 13280
rect 11681 13277 11693 13280
rect 11727 13277 11739 13311
rect 11681 13271 11739 13277
rect 14366 13268 14372 13320
rect 14424 13268 14430 13320
rect 14458 13268 14464 13320
rect 14516 13268 14522 13320
rect 19797 13311 19855 13317
rect 19797 13277 19809 13311
rect 19843 13277 19855 13311
rect 19797 13271 19855 13277
rect 5322 13243 5380 13249
rect 5322 13240 5334 13243
rect 4448 13212 5334 13240
rect 4448 13181 4476 13212
rect 5322 13209 5334 13212
rect 5368 13209 5380 13243
rect 7285 13243 7343 13249
rect 7285 13240 7297 13243
rect 5322 13203 5380 13209
rect 6886 13212 7297 13240
rect 4433 13175 4491 13181
rect 4433 13141 4445 13175
rect 4479 13141 4491 13175
rect 4433 13135 4491 13141
rect 6457 13175 6515 13181
rect 6457 13141 6469 13175
rect 6503 13172 6515 13175
rect 6886 13172 6914 13212
rect 7285 13209 7297 13212
rect 7331 13209 7343 13243
rect 7285 13203 7343 13209
rect 10597 13243 10655 13249
rect 10597 13209 10609 13243
rect 10643 13240 10655 13243
rect 11790 13240 11796 13252
rect 10643 13212 11796 13240
rect 10643 13209 10655 13212
rect 10597 13203 10655 13209
rect 11790 13200 11796 13212
rect 11848 13200 11854 13252
rect 17405 13243 17463 13249
rect 17405 13209 17417 13243
rect 17451 13209 17463 13243
rect 17405 13203 17463 13209
rect 6503 13144 6914 13172
rect 6503 13141 6515 13144
rect 6457 13135 6515 13141
rect 7374 13132 7380 13184
rect 7432 13132 7438 13184
rect 10229 13175 10287 13181
rect 10229 13141 10241 13175
rect 10275 13172 10287 13175
rect 10318 13172 10324 13184
rect 10275 13144 10324 13172
rect 10275 13141 10287 13144
rect 10229 13135 10287 13141
rect 10318 13132 10324 13144
rect 10376 13132 10382 13184
rect 10689 13175 10747 13181
rect 10689 13141 10701 13175
rect 10735 13172 10747 13175
rect 11698 13172 11704 13184
rect 10735 13144 11704 13172
rect 10735 13141 10747 13144
rect 10689 13135 10747 13141
rect 11698 13132 11704 13144
rect 11756 13132 11762 13184
rect 12802 13132 12808 13184
rect 12860 13132 12866 13184
rect 17420 13172 17448 13203
rect 17954 13200 17960 13252
rect 18012 13200 18018 13252
rect 19812 13240 19840 13271
rect 19978 13268 19984 13320
rect 20036 13268 20042 13320
rect 20073 13311 20131 13317
rect 20073 13277 20085 13311
rect 20119 13308 20131 13311
rect 20622 13308 20628 13320
rect 20119 13280 20628 13308
rect 20119 13277 20131 13280
rect 20073 13271 20131 13277
rect 20622 13268 20628 13280
rect 20680 13268 20686 13320
rect 20809 13311 20867 13317
rect 20809 13277 20821 13311
rect 20855 13308 20867 13311
rect 21008 13308 21036 13348
rect 21542 13336 21548 13348
rect 21600 13336 21606 13388
rect 21652 13376 21680 13416
rect 22002 13376 22008 13388
rect 21652 13348 22008 13376
rect 22002 13336 22008 13348
rect 22060 13376 22066 13388
rect 22189 13379 22247 13385
rect 22189 13376 22201 13379
rect 22060 13348 22201 13376
rect 22060 13336 22066 13348
rect 22189 13345 22201 13348
rect 22235 13345 22247 13379
rect 22189 13339 22247 13345
rect 20855 13280 21036 13308
rect 20855 13277 20867 13280
rect 20809 13271 20867 13277
rect 21450 13268 21456 13320
rect 21508 13268 21514 13320
rect 22278 13268 22284 13320
rect 22336 13308 22342 13320
rect 22388 13317 22416 13416
rect 28813 13413 28825 13447
rect 28859 13444 28871 13447
rect 30282 13444 30288 13456
rect 28859 13416 30288 13444
rect 28859 13413 28871 13416
rect 28813 13407 28871 13413
rect 30282 13404 30288 13416
rect 30340 13404 30346 13456
rect 30558 13444 30564 13456
rect 30484 13416 30564 13444
rect 22646 13336 22652 13388
rect 22704 13376 22710 13388
rect 26326 13376 26332 13388
rect 22704 13348 26332 13376
rect 22704 13336 22710 13348
rect 26326 13336 26332 13348
rect 26384 13336 26390 13388
rect 30484 13376 30512 13416
rect 30558 13404 30564 13416
rect 30616 13444 30622 13456
rect 31478 13444 31484 13456
rect 30616 13416 31484 13444
rect 30616 13404 30622 13416
rect 31478 13404 31484 13416
rect 31536 13404 31542 13456
rect 31754 13404 31760 13456
rect 31812 13444 31818 13456
rect 31849 13447 31907 13453
rect 31849 13444 31861 13447
rect 31812 13416 31861 13444
rect 31812 13404 31818 13416
rect 31849 13413 31861 13416
rect 31895 13444 31907 13447
rect 32398 13444 32404 13456
rect 31895 13416 32404 13444
rect 31895 13413 31907 13416
rect 31849 13407 31907 13413
rect 32398 13404 32404 13416
rect 32456 13444 32462 13456
rect 40221 13447 40279 13453
rect 32456 13416 33456 13444
rect 32456 13404 32462 13416
rect 28736 13348 30512 13376
rect 22373 13311 22431 13317
rect 22373 13308 22385 13311
rect 22336 13280 22385 13308
rect 22336 13268 22342 13280
rect 22373 13277 22385 13280
rect 22419 13277 22431 13311
rect 22373 13271 22431 13277
rect 22557 13311 22615 13317
rect 22557 13277 22569 13311
rect 22603 13308 22615 13311
rect 23753 13311 23811 13317
rect 23753 13308 23765 13311
rect 22603 13280 23765 13308
rect 22603 13277 22615 13280
rect 22557 13271 22615 13277
rect 23753 13277 23765 13280
rect 23799 13277 23811 13311
rect 23753 13271 23811 13277
rect 24578 13268 24584 13320
rect 24636 13268 24642 13320
rect 26970 13268 26976 13320
rect 27028 13268 27034 13320
rect 27154 13268 27160 13320
rect 27212 13308 27218 13320
rect 28736 13317 28764 13348
rect 28721 13311 28779 13317
rect 28721 13308 28733 13311
rect 27212 13280 28733 13308
rect 27212 13268 27218 13280
rect 28721 13277 28733 13280
rect 28767 13277 28779 13311
rect 28721 13271 28779 13277
rect 28902 13268 28908 13320
rect 28960 13268 28966 13320
rect 29914 13268 29920 13320
rect 29972 13268 29978 13320
rect 30024 13317 30052 13348
rect 30926 13336 30932 13388
rect 30984 13336 30990 13388
rect 32508 13348 33180 13376
rect 30009 13311 30067 13317
rect 30009 13277 30021 13311
rect 30055 13277 30067 13311
rect 30009 13271 30067 13277
rect 30558 13268 30564 13320
rect 30616 13308 30622 13320
rect 31021 13311 31079 13317
rect 31021 13308 31033 13311
rect 30616 13280 31033 13308
rect 30616 13268 30622 13280
rect 31021 13277 31033 13280
rect 31067 13277 31079 13311
rect 31021 13271 31079 13277
rect 32304 13311 32362 13317
rect 32304 13277 32316 13311
rect 32350 13308 32362 13311
rect 32508 13308 32536 13348
rect 33152 13320 33180 13348
rect 32350 13280 32536 13308
rect 32350 13277 32362 13280
rect 32304 13271 32362 13277
rect 32674 13268 32680 13320
rect 32732 13268 32738 13320
rect 32766 13268 32772 13320
rect 32824 13268 32830 13320
rect 33134 13268 33140 13320
rect 33192 13308 33198 13320
rect 33428 13317 33456 13416
rect 40221 13413 40233 13447
rect 40267 13413 40279 13447
rect 40221 13407 40279 13413
rect 36078 13336 36084 13388
rect 36136 13336 36142 13388
rect 36814 13336 36820 13388
rect 36872 13376 36878 13388
rect 36909 13379 36967 13385
rect 36909 13376 36921 13379
rect 36872 13348 36921 13376
rect 36872 13336 36878 13348
rect 36909 13345 36921 13348
rect 36955 13345 36967 13379
rect 40236 13376 40264 13407
rect 40236 13348 41092 13376
rect 36909 13339 36967 13345
rect 33229 13311 33287 13317
rect 33229 13308 33241 13311
rect 33192 13280 33241 13308
rect 33192 13268 33198 13280
rect 33229 13277 33241 13280
rect 33275 13277 33287 13311
rect 33229 13271 33287 13277
rect 33413 13311 33471 13317
rect 33413 13277 33425 13311
rect 33459 13308 33471 13311
rect 35437 13311 35495 13317
rect 35437 13308 35449 13311
rect 33459 13280 35449 13308
rect 33459 13277 33471 13280
rect 33413 13271 33471 13277
rect 35437 13277 35449 13280
rect 35483 13277 35495 13311
rect 35437 13271 35495 13277
rect 20533 13243 20591 13249
rect 19812 13212 20116 13240
rect 18046 13172 18052 13184
rect 17420 13144 18052 13172
rect 18046 13132 18052 13144
rect 18104 13132 18110 13184
rect 20088 13172 20116 13212
rect 20533 13209 20545 13243
rect 20579 13240 20591 13243
rect 20714 13240 20720 13252
rect 20579 13212 20720 13240
rect 20579 13209 20591 13212
rect 20533 13203 20591 13209
rect 20714 13200 20720 13212
rect 20772 13200 20778 13252
rect 22646 13240 22652 13252
rect 20824 13212 22652 13240
rect 20824 13172 20852 13212
rect 22646 13200 22652 13212
rect 22704 13200 22710 13252
rect 24857 13243 24915 13249
rect 24857 13209 24869 13243
rect 24903 13209 24915 13243
rect 26878 13240 26884 13252
rect 26082 13212 26884 13240
rect 24857 13203 24915 13209
rect 20088 13144 20852 13172
rect 20990 13132 20996 13184
rect 21048 13132 21054 13184
rect 23569 13175 23627 13181
rect 23569 13141 23581 13175
rect 23615 13172 23627 13175
rect 24872 13172 24900 13203
rect 26878 13200 26884 13212
rect 26936 13200 26942 13252
rect 29733 13243 29791 13249
rect 29733 13209 29745 13243
rect 29779 13240 29791 13243
rect 30926 13240 30932 13252
rect 29779 13212 30932 13240
rect 29779 13209 29791 13212
rect 29733 13203 29791 13209
rect 30926 13200 30932 13212
rect 30984 13240 30990 13252
rect 31846 13240 31852 13252
rect 30984 13212 31852 13240
rect 30984 13200 30990 13212
rect 31846 13200 31852 13212
rect 31904 13200 31910 13252
rect 32048 13212 32260 13240
rect 23615 13144 24900 13172
rect 31389 13175 31447 13181
rect 23615 13141 23627 13144
rect 23569 13135 23627 13141
rect 31389 13141 31401 13175
rect 31435 13172 31447 13175
rect 32048 13172 32076 13212
rect 31435 13144 32076 13172
rect 32232 13172 32260 13212
rect 32398 13200 32404 13252
rect 32456 13200 32462 13252
rect 32490 13200 32496 13252
rect 32548 13200 32554 13252
rect 35710 13240 35716 13252
rect 32600 13212 35716 13240
rect 32600 13172 32628 13212
rect 35710 13200 35716 13212
rect 35768 13200 35774 13252
rect 36096 13240 36124 13336
rect 36262 13268 36268 13320
rect 36320 13268 36326 13320
rect 37176 13311 37234 13317
rect 37176 13277 37188 13311
rect 37222 13308 37234 13311
rect 37458 13308 37464 13320
rect 37222 13280 37464 13308
rect 37222 13277 37234 13280
rect 37176 13271 37234 13277
rect 37458 13268 37464 13280
rect 37516 13268 37522 13320
rect 40494 13268 40500 13320
rect 40552 13268 40558 13320
rect 40586 13268 40592 13320
rect 40644 13308 40650 13320
rect 40957 13311 41015 13317
rect 40957 13308 40969 13311
rect 40644 13280 40969 13308
rect 40644 13268 40650 13280
rect 40957 13277 40969 13280
rect 41003 13277 41015 13311
rect 41064 13308 41092 13348
rect 41966 13336 41972 13388
rect 42024 13376 42030 13388
rect 42024 13348 43300 13376
rect 42024 13336 42030 13348
rect 41213 13311 41271 13317
rect 41213 13308 41225 13311
rect 41064 13280 41225 13308
rect 40957 13271 41015 13277
rect 41213 13277 41225 13280
rect 41259 13277 41271 13311
rect 41213 13271 41271 13277
rect 42058 13268 42064 13320
rect 42116 13308 42122 13320
rect 43272 13317 43300 13348
rect 42981 13311 43039 13317
rect 42981 13308 42993 13311
rect 42116 13280 42993 13308
rect 42116 13268 42122 13280
rect 42981 13277 42993 13280
rect 43027 13277 43039 13311
rect 42981 13271 43039 13277
rect 43257 13311 43315 13317
rect 43257 13277 43269 13311
rect 43303 13277 43315 13311
rect 43257 13271 43315 13277
rect 40126 13240 40132 13252
rect 36096 13212 40132 13240
rect 40126 13200 40132 13212
rect 40184 13200 40190 13252
rect 40221 13243 40279 13249
rect 40221 13209 40233 13243
rect 40267 13240 40279 13243
rect 41046 13240 41052 13252
rect 40267 13212 41052 13240
rect 40267 13209 40279 13212
rect 40221 13203 40279 13209
rect 41046 13200 41052 13212
rect 41104 13200 41110 13252
rect 41690 13200 41696 13252
rect 41748 13240 41754 13252
rect 43165 13243 43223 13249
rect 43165 13240 43177 13243
rect 41748 13212 43177 13240
rect 41748 13200 41754 13212
rect 43165 13209 43177 13212
rect 43211 13209 43223 13243
rect 43165 13203 43223 13209
rect 32232 13144 32628 13172
rect 31435 13141 31447 13144
rect 31389 13135 31447 13141
rect 32674 13132 32680 13184
rect 32732 13172 32738 13184
rect 33321 13175 33379 13181
rect 33321 13172 33333 13175
rect 32732 13144 33333 13172
rect 32732 13132 32738 13144
rect 33321 13141 33333 13144
rect 33367 13141 33379 13175
rect 33321 13135 33379 13141
rect 36446 13132 36452 13184
rect 36504 13132 36510 13184
rect 38289 13175 38347 13181
rect 38289 13141 38301 13175
rect 38335 13172 38347 13175
rect 38378 13172 38384 13184
rect 38335 13144 38384 13172
rect 38335 13141 38347 13144
rect 38289 13135 38347 13141
rect 38378 13132 38384 13144
rect 38436 13172 38442 13184
rect 38654 13172 38660 13184
rect 38436 13144 38660 13172
rect 38436 13132 38442 13144
rect 38654 13132 38660 13144
rect 38712 13132 38718 13184
rect 40402 13132 40408 13184
rect 40460 13132 40466 13184
rect 42334 13132 42340 13184
rect 42392 13132 42398 13184
rect 1104 13082 45051 13104
rect 1104 13030 11896 13082
rect 11948 13030 11960 13082
rect 12012 13030 12024 13082
rect 12076 13030 12088 13082
rect 12140 13030 12152 13082
rect 12204 13030 22843 13082
rect 22895 13030 22907 13082
rect 22959 13030 22971 13082
rect 23023 13030 23035 13082
rect 23087 13030 23099 13082
rect 23151 13030 33790 13082
rect 33842 13030 33854 13082
rect 33906 13030 33918 13082
rect 33970 13030 33982 13082
rect 34034 13030 34046 13082
rect 34098 13030 44737 13082
rect 44789 13030 44801 13082
rect 44853 13030 44865 13082
rect 44917 13030 44929 13082
rect 44981 13030 44993 13082
rect 45045 13030 45051 13082
rect 1104 13008 45051 13030
rect 5350 12928 5356 12980
rect 5408 12968 5414 12980
rect 5445 12971 5503 12977
rect 5445 12968 5457 12971
rect 5408 12940 5457 12968
rect 5408 12928 5414 12940
rect 5445 12937 5457 12940
rect 5491 12937 5503 12971
rect 5445 12931 5503 12937
rect 11698 12928 11704 12980
rect 11756 12928 11762 12980
rect 12161 12971 12219 12977
rect 12161 12937 12173 12971
rect 12207 12968 12219 12971
rect 14550 12968 14556 12980
rect 12207 12940 14556 12968
rect 12207 12937 12219 12940
rect 12161 12931 12219 12937
rect 14550 12928 14556 12940
rect 14608 12928 14614 12980
rect 15013 12971 15071 12977
rect 15013 12937 15025 12971
rect 15059 12937 15071 12971
rect 15013 12931 15071 12937
rect 20257 12971 20315 12977
rect 20257 12937 20269 12971
rect 20303 12968 20315 12971
rect 20806 12968 20812 12980
rect 20303 12940 20812 12968
rect 20303 12937 20315 12940
rect 20257 12931 20315 12937
rect 9858 12900 9864 12912
rect 6564 12872 9864 12900
rect 3142 12792 3148 12844
rect 3200 12792 3206 12844
rect 3970 12792 3976 12844
rect 4028 12832 4034 12844
rect 4338 12841 4344 12844
rect 4065 12835 4123 12841
rect 4065 12832 4077 12835
rect 4028 12804 4077 12832
rect 4028 12792 4034 12804
rect 4065 12801 4077 12804
rect 4111 12801 4123 12835
rect 4332 12832 4344 12841
rect 4299 12804 4344 12832
rect 4065 12795 4123 12801
rect 4332 12795 4344 12804
rect 4396 12832 4402 12844
rect 4798 12832 4804 12844
rect 4396 12804 4804 12832
rect 4338 12792 4344 12795
rect 4396 12792 4402 12804
rect 4798 12792 4804 12804
rect 4856 12792 4862 12844
rect 5074 12724 5080 12776
rect 5132 12764 5138 12776
rect 6564 12773 6592 12872
rect 6816 12835 6874 12841
rect 6816 12801 6828 12835
rect 6862 12832 6874 12835
rect 6862 12804 8432 12832
rect 6862 12801 6874 12804
rect 6816 12795 6874 12801
rect 6549 12767 6607 12773
rect 6549 12764 6561 12767
rect 5132 12736 6561 12764
rect 5132 12724 5138 12736
rect 6549 12733 6561 12736
rect 6595 12733 6607 12767
rect 6549 12727 6607 12733
rect 8404 12705 8432 12804
rect 8570 12792 8576 12844
rect 8628 12792 8634 12844
rect 9784 12841 9812 12872
rect 9858 12860 9864 12872
rect 9916 12900 9922 12912
rect 11422 12900 11428 12912
rect 9916 12872 11428 12900
rect 9916 12860 9922 12872
rect 11422 12860 11428 12872
rect 11480 12860 11486 12912
rect 13440 12903 13498 12909
rect 13440 12869 13452 12903
rect 13486 12900 13498 12903
rect 15028 12900 15056 12931
rect 20806 12928 20812 12940
rect 20864 12928 20870 12980
rect 22186 12968 22192 12980
rect 21008 12940 22192 12968
rect 13486 12872 15056 12900
rect 17957 12903 18015 12909
rect 13486 12869 13498 12872
rect 13440 12863 13498 12869
rect 17957 12869 17969 12903
rect 18003 12900 18015 12903
rect 18003 12872 19274 12900
rect 18003 12869 18015 12872
rect 17957 12863 18015 12869
rect 10042 12841 10048 12844
rect 9769 12835 9827 12841
rect 9769 12801 9781 12835
rect 9815 12801 9827 12835
rect 9769 12795 9827 12801
rect 10036 12795 10048 12841
rect 10042 12792 10048 12795
rect 10100 12792 10106 12844
rect 11146 12792 11152 12844
rect 11204 12832 11210 12844
rect 12069 12835 12127 12841
rect 12069 12832 12081 12835
rect 11204 12804 12081 12832
rect 11204 12792 11210 12804
rect 12069 12801 12081 12804
rect 12115 12801 12127 12835
rect 12069 12795 12127 12801
rect 13814 12792 13820 12844
rect 13872 12832 13878 12844
rect 15197 12835 15255 12841
rect 15197 12832 15209 12835
rect 13872 12804 15209 12832
rect 13872 12792 13878 12804
rect 15197 12801 15209 12804
rect 15243 12801 15255 12835
rect 15197 12795 15255 12801
rect 17218 12792 17224 12844
rect 17276 12832 17282 12844
rect 17865 12835 17923 12841
rect 17865 12832 17877 12835
rect 17276 12804 17877 12832
rect 17276 12792 17282 12804
rect 17865 12801 17877 12804
rect 17911 12801 17923 12835
rect 17865 12795 17923 12801
rect 12342 12724 12348 12776
rect 12400 12724 12406 12776
rect 13170 12724 13176 12776
rect 13228 12724 13234 12776
rect 17880 12764 17908 12795
rect 18138 12792 18144 12844
rect 18196 12832 18202 12844
rect 18506 12832 18512 12844
rect 18196 12804 18512 12832
rect 18196 12792 18202 12804
rect 18506 12792 18512 12804
rect 18564 12792 18570 12844
rect 20898 12792 20904 12844
rect 20956 12792 20962 12844
rect 21008 12841 21036 12940
rect 22186 12928 22192 12940
rect 22244 12928 22250 12980
rect 22373 12971 22431 12977
rect 22373 12937 22385 12971
rect 22419 12968 22431 12971
rect 22462 12968 22468 12980
rect 22419 12940 22468 12968
rect 22419 12937 22431 12940
rect 22373 12931 22431 12937
rect 22462 12928 22468 12940
rect 22520 12928 22526 12980
rect 27154 12928 27160 12980
rect 27212 12968 27218 12980
rect 27341 12971 27399 12977
rect 27341 12968 27353 12971
rect 27212 12940 27353 12968
rect 27212 12928 27218 12940
rect 27341 12937 27353 12940
rect 27387 12937 27399 12971
rect 27341 12931 27399 12937
rect 31389 12971 31447 12977
rect 31389 12937 31401 12971
rect 31435 12968 31447 12971
rect 31938 12968 31944 12980
rect 31435 12940 31944 12968
rect 31435 12937 31447 12940
rect 31389 12931 31447 12937
rect 31938 12928 31944 12940
rect 31996 12928 32002 12980
rect 33042 12928 33048 12980
rect 33100 12968 33106 12980
rect 33613 12971 33671 12977
rect 33613 12968 33625 12971
rect 33100 12940 33625 12968
rect 33100 12928 33106 12940
rect 33613 12937 33625 12940
rect 33659 12937 33671 12971
rect 33613 12931 33671 12937
rect 33781 12971 33839 12977
rect 33781 12937 33793 12971
rect 33827 12937 33839 12971
rect 37461 12971 37519 12977
rect 37461 12968 37473 12971
rect 33781 12931 33839 12937
rect 35084 12940 37473 12968
rect 24872 12872 31432 12900
rect 20993 12835 21051 12841
rect 20993 12801 21005 12835
rect 21039 12801 21051 12835
rect 20993 12795 21051 12801
rect 21082 12792 21088 12844
rect 21140 12792 21146 12844
rect 21223 12835 21281 12841
rect 21223 12832 21235 12835
rect 21218 12801 21235 12832
rect 21269 12801 21281 12835
rect 21218 12795 21281 12801
rect 17954 12764 17960 12776
rect 17880 12736 17960 12764
rect 17954 12724 17960 12736
rect 18012 12724 18018 12776
rect 18785 12767 18843 12773
rect 18785 12733 18797 12767
rect 18831 12764 18843 12767
rect 20717 12767 20775 12773
rect 20717 12764 20729 12767
rect 18831 12736 20729 12764
rect 18831 12733 18843 12736
rect 18785 12727 18843 12733
rect 20717 12733 20729 12736
rect 20763 12733 20775 12767
rect 20717 12727 20775 12733
rect 20806 12724 20812 12776
rect 20864 12764 20870 12776
rect 21218 12764 21246 12795
rect 22002 12792 22008 12844
rect 22060 12792 22066 12844
rect 24872 12841 24900 12872
rect 24857 12835 24915 12841
rect 24857 12801 24869 12835
rect 24903 12801 24915 12835
rect 24857 12795 24915 12801
rect 25222 12792 25228 12844
rect 25280 12832 25286 12844
rect 25869 12835 25927 12841
rect 25869 12832 25881 12835
rect 25280 12804 25881 12832
rect 25280 12792 25286 12804
rect 25869 12801 25881 12804
rect 25915 12801 25927 12835
rect 25869 12795 25927 12801
rect 25958 12792 25964 12844
rect 26016 12832 26022 12844
rect 26053 12835 26111 12841
rect 26053 12832 26065 12835
rect 26016 12804 26065 12832
rect 26016 12792 26022 12804
rect 26053 12801 26065 12804
rect 26099 12801 26111 12835
rect 26053 12795 26111 12801
rect 26237 12835 26295 12841
rect 26237 12801 26249 12835
rect 26283 12832 26295 12835
rect 27249 12835 27307 12841
rect 27249 12832 27261 12835
rect 26283 12804 27261 12832
rect 26283 12801 26295 12804
rect 26237 12795 26295 12801
rect 27249 12801 27261 12804
rect 27295 12801 27307 12835
rect 27249 12795 27307 12801
rect 29178 12792 29184 12844
rect 29236 12792 29242 12844
rect 29454 12841 29460 12844
rect 29448 12795 29460 12841
rect 29454 12792 29460 12795
rect 29512 12792 29518 12844
rect 20864 12736 21246 12764
rect 21361 12767 21419 12773
rect 20864 12724 20870 12736
rect 21361 12733 21373 12767
rect 21407 12764 21419 12767
rect 21450 12764 21456 12776
rect 21407 12736 21456 12764
rect 21407 12733 21419 12736
rect 21361 12727 21419 12733
rect 8389 12699 8447 12705
rect 8389 12665 8401 12699
rect 8435 12665 8447 12699
rect 21266 12696 21272 12708
rect 8389 12659 8447 12665
rect 20548 12668 21272 12696
rect 2774 12588 2780 12640
rect 2832 12628 2838 12640
rect 2961 12631 3019 12637
rect 2961 12628 2973 12631
rect 2832 12600 2973 12628
rect 2832 12588 2838 12600
rect 2961 12597 2973 12600
rect 3007 12597 3019 12631
rect 2961 12591 3019 12597
rect 7742 12588 7748 12640
rect 7800 12628 7806 12640
rect 7929 12631 7987 12637
rect 7929 12628 7941 12631
rect 7800 12600 7941 12628
rect 7800 12588 7806 12600
rect 7929 12597 7941 12600
rect 7975 12597 7987 12631
rect 7929 12591 7987 12597
rect 11146 12588 11152 12640
rect 11204 12588 11210 12640
rect 14090 12588 14096 12640
rect 14148 12628 14154 12640
rect 14366 12628 14372 12640
rect 14148 12600 14372 12628
rect 14148 12588 14154 12600
rect 14366 12588 14372 12600
rect 14424 12628 14430 12640
rect 20548 12628 20576 12668
rect 21266 12656 21272 12668
rect 21324 12656 21330 12708
rect 14424 12600 20576 12628
rect 14424 12588 14430 12600
rect 20622 12588 20628 12640
rect 20680 12628 20686 12640
rect 21376 12628 21404 12727
rect 21450 12724 21456 12736
rect 21508 12724 21514 12776
rect 22097 12767 22155 12773
rect 22097 12733 22109 12767
rect 22143 12733 22155 12767
rect 22097 12727 22155 12733
rect 21542 12656 21548 12708
rect 21600 12696 21606 12708
rect 22112 12696 22140 12727
rect 22186 12724 22192 12776
rect 22244 12764 22250 12776
rect 24670 12764 24676 12776
rect 22244 12736 24676 12764
rect 22244 12724 22250 12736
rect 24670 12724 24676 12736
rect 24728 12764 24734 12776
rect 24949 12767 25007 12773
rect 24949 12764 24961 12767
rect 24728 12736 24961 12764
rect 24728 12724 24734 12736
rect 24949 12733 24961 12736
rect 24995 12733 25007 12767
rect 31404 12764 31432 12872
rect 31478 12860 31484 12912
rect 31536 12860 31542 12912
rect 32309 12903 32367 12909
rect 32309 12869 32321 12903
rect 32355 12900 32367 12903
rect 33226 12900 33232 12912
rect 32355 12872 33232 12900
rect 32355 12869 32367 12872
rect 32309 12863 32367 12869
rect 33226 12860 33232 12872
rect 33284 12860 33290 12912
rect 33410 12860 33416 12912
rect 33468 12860 33474 12912
rect 33796 12900 33824 12931
rect 34425 12903 34483 12909
rect 34425 12900 34437 12903
rect 33796 12872 34437 12900
rect 34425 12869 34437 12872
rect 34471 12869 34483 12903
rect 34425 12863 34483 12869
rect 31570 12792 31576 12844
rect 31628 12792 31634 12844
rect 31757 12835 31815 12841
rect 31757 12801 31769 12835
rect 31803 12832 31815 12835
rect 32582 12832 32588 12844
rect 31803 12804 32588 12832
rect 31803 12801 31815 12804
rect 31757 12795 31815 12801
rect 32582 12792 32588 12804
rect 32640 12792 32646 12844
rect 32674 12792 32680 12844
rect 32732 12792 32738 12844
rect 32769 12835 32827 12841
rect 32769 12801 32781 12835
rect 32815 12832 32827 12835
rect 35084 12832 35112 12940
rect 37461 12937 37473 12940
rect 37507 12937 37519 12971
rect 37461 12931 37519 12937
rect 37550 12928 37556 12980
rect 37608 12968 37614 12980
rect 38381 12971 38439 12977
rect 38381 12968 38393 12971
rect 37608 12940 38393 12968
rect 37608 12928 37614 12940
rect 38381 12937 38393 12940
rect 38427 12937 38439 12971
rect 40034 12968 40040 12980
rect 38381 12931 38439 12937
rect 38580 12940 40040 12968
rect 36170 12900 36176 12912
rect 35452 12872 36176 12900
rect 35452 12841 35480 12872
rect 36170 12860 36176 12872
rect 36228 12860 36234 12912
rect 36354 12860 36360 12912
rect 36412 12900 36418 12912
rect 38580 12900 38608 12940
rect 40034 12928 40040 12940
rect 40092 12928 40098 12980
rect 40221 12971 40279 12977
rect 40221 12937 40233 12971
rect 40267 12968 40279 12971
rect 40310 12968 40316 12980
rect 40267 12940 40316 12968
rect 40267 12937 40279 12940
rect 40221 12931 40279 12937
rect 40310 12928 40316 12940
rect 40368 12928 40374 12980
rect 40405 12971 40463 12977
rect 40405 12937 40417 12971
rect 40451 12968 40463 12971
rect 40494 12968 40500 12980
rect 40451 12940 40500 12968
rect 40451 12937 40463 12940
rect 40405 12931 40463 12937
rect 40494 12928 40500 12940
rect 40552 12928 40558 12980
rect 41046 12928 41052 12980
rect 41104 12968 41110 12980
rect 41233 12971 41291 12977
rect 41233 12968 41245 12971
rect 41104 12940 41245 12968
rect 41104 12928 41110 12940
rect 41233 12937 41245 12940
rect 41279 12937 41291 12971
rect 41601 12971 41659 12977
rect 41601 12968 41613 12971
rect 41233 12931 41291 12937
rect 41386 12940 41613 12968
rect 39758 12900 39764 12912
rect 36412 12872 38608 12900
rect 36412 12860 36418 12872
rect 32815 12804 35112 12832
rect 35437 12835 35495 12841
rect 32815 12801 32827 12804
rect 32769 12795 32827 12801
rect 35437 12801 35449 12835
rect 35483 12801 35495 12835
rect 35437 12795 35495 12801
rect 35618 12792 35624 12844
rect 35676 12792 35682 12844
rect 35710 12792 35716 12844
rect 35768 12832 35774 12844
rect 36081 12835 36139 12841
rect 36081 12832 36093 12835
rect 35768 12804 36093 12832
rect 35768 12792 35774 12804
rect 36081 12801 36093 12804
rect 36127 12801 36139 12835
rect 36081 12795 36139 12801
rect 36262 12792 36268 12844
rect 36320 12792 36326 12844
rect 36446 12792 36452 12844
rect 36504 12792 36510 12844
rect 36630 12792 36636 12844
rect 36688 12792 36694 12844
rect 37642 12792 37648 12844
rect 37700 12792 37706 12844
rect 37829 12835 37887 12841
rect 37829 12801 37841 12835
rect 37875 12801 37887 12835
rect 37829 12795 37887 12801
rect 32490 12764 32496 12776
rect 31404 12736 32496 12764
rect 24949 12727 25007 12733
rect 32490 12724 32496 12736
rect 32548 12724 32554 12776
rect 35529 12767 35587 12773
rect 35529 12733 35541 12767
rect 35575 12764 35587 12767
rect 36357 12767 36415 12773
rect 36357 12764 36369 12767
rect 35575 12736 36369 12764
rect 35575 12733 35587 12736
rect 35529 12727 35587 12733
rect 36357 12733 36369 12736
rect 36403 12733 36415 12767
rect 36357 12727 36415 12733
rect 21600 12668 22140 12696
rect 21600 12656 21606 12668
rect 22278 12656 22284 12708
rect 22336 12696 22342 12708
rect 23106 12696 23112 12708
rect 22336 12668 23112 12696
rect 22336 12656 22342 12668
rect 23106 12656 23112 12668
rect 23164 12656 23170 12708
rect 31205 12699 31263 12705
rect 31205 12665 31217 12699
rect 31251 12696 31263 12699
rect 32122 12696 32128 12708
rect 31251 12668 32128 12696
rect 31251 12665 31263 12668
rect 31205 12659 31263 12665
rect 32122 12656 32128 12668
rect 32180 12656 32186 12708
rect 33502 12656 33508 12708
rect 33560 12696 33566 12708
rect 34609 12699 34667 12705
rect 33560 12668 33732 12696
rect 33560 12656 33566 12668
rect 22094 12628 22100 12640
rect 20680 12600 22100 12628
rect 20680 12588 20686 12600
rect 22094 12588 22100 12600
rect 22152 12588 22158 12640
rect 22189 12631 22247 12637
rect 22189 12597 22201 12631
rect 22235 12628 22247 12631
rect 22646 12628 22652 12640
rect 22235 12600 22652 12628
rect 22235 12597 22247 12600
rect 22189 12591 22247 12597
rect 22646 12588 22652 12600
rect 22704 12588 22710 12640
rect 30558 12588 30564 12640
rect 30616 12588 30622 12640
rect 31938 12588 31944 12640
rect 31996 12628 32002 12640
rect 32953 12631 33011 12637
rect 32953 12628 32965 12631
rect 31996 12600 32965 12628
rect 31996 12588 32002 12600
rect 32953 12597 32965 12600
rect 32999 12628 33011 12631
rect 33597 12631 33655 12637
rect 33597 12628 33609 12631
rect 32999 12600 33609 12628
rect 32999 12597 33011 12600
rect 32953 12591 33011 12597
rect 33597 12597 33609 12600
rect 33643 12597 33655 12631
rect 33704 12628 33732 12668
rect 34609 12665 34621 12699
rect 34655 12696 34667 12699
rect 36078 12696 36084 12708
rect 34655 12668 36084 12696
rect 34655 12665 34667 12668
rect 34609 12659 34667 12665
rect 36078 12656 36084 12668
rect 36136 12656 36142 12708
rect 37844 12696 37872 12795
rect 37918 12792 37924 12844
rect 37976 12832 37982 12844
rect 38580 12841 38608 12872
rect 38856 12872 39764 12900
rect 38565 12835 38623 12841
rect 37976 12804 38424 12832
rect 37976 12792 37982 12804
rect 38396 12764 38424 12804
rect 38565 12801 38577 12835
rect 38611 12801 38623 12835
rect 38565 12795 38623 12801
rect 38654 12792 38660 12844
rect 38712 12832 38718 12844
rect 38856 12841 38884 12872
rect 39758 12860 39764 12872
rect 39816 12900 39822 12912
rect 40129 12903 40187 12909
rect 40129 12900 40141 12903
rect 39816 12872 40141 12900
rect 39816 12860 39822 12872
rect 40129 12869 40141 12872
rect 40175 12869 40187 12903
rect 40129 12863 40187 12869
rect 38749 12835 38807 12841
rect 38749 12832 38761 12835
rect 38712 12804 38761 12832
rect 38712 12792 38718 12804
rect 38749 12801 38761 12804
rect 38795 12801 38807 12835
rect 38749 12795 38807 12801
rect 38841 12835 38899 12841
rect 38841 12801 38853 12835
rect 38887 12801 38899 12835
rect 38841 12795 38899 12801
rect 39301 12835 39359 12841
rect 39301 12801 39313 12835
rect 39347 12801 39359 12835
rect 39301 12795 39359 12801
rect 39485 12835 39543 12841
rect 39485 12801 39497 12835
rect 39531 12801 39543 12835
rect 39485 12795 39543 12801
rect 40037 12835 40095 12841
rect 40037 12801 40049 12835
rect 40083 12801 40095 12835
rect 41386 12832 41414 12940
rect 41601 12937 41613 12940
rect 41647 12968 41659 12971
rect 42058 12968 42064 12980
rect 41647 12940 42064 12968
rect 41647 12937 41659 12940
rect 41601 12931 41659 12937
rect 42058 12928 42064 12940
rect 42116 12928 42122 12980
rect 40037 12795 40095 12801
rect 40420 12804 41414 12832
rect 39316 12764 39344 12795
rect 38396 12736 39344 12764
rect 39390 12724 39396 12776
rect 39448 12724 39454 12776
rect 38562 12696 38568 12708
rect 36188 12668 37504 12696
rect 37844 12668 38568 12696
rect 36188 12628 36216 12668
rect 33704 12600 36216 12628
rect 36817 12631 36875 12637
rect 33597 12591 33655 12597
rect 36817 12597 36829 12631
rect 36863 12628 36875 12631
rect 37366 12628 37372 12640
rect 36863 12600 37372 12628
rect 36863 12597 36875 12600
rect 36817 12591 36875 12597
rect 37366 12588 37372 12600
rect 37424 12588 37430 12640
rect 37476 12628 37504 12668
rect 38562 12656 38568 12668
rect 38620 12696 38626 12708
rect 39500 12696 39528 12795
rect 38620 12668 39528 12696
rect 38620 12656 38626 12668
rect 40052 12628 40080 12795
rect 40126 12724 40132 12776
rect 40184 12764 40190 12776
rect 40420 12773 40448 12804
rect 41506 12792 41512 12844
rect 41564 12832 41570 12844
rect 42334 12832 42340 12844
rect 41564 12804 42340 12832
rect 41564 12792 41570 12804
rect 42334 12792 42340 12804
rect 42392 12792 42398 12844
rect 40405 12767 40463 12773
rect 40405 12764 40417 12767
rect 40184 12736 40417 12764
rect 40184 12724 40190 12736
rect 40405 12733 40417 12736
rect 40451 12733 40463 12767
rect 40405 12727 40463 12733
rect 41417 12767 41475 12773
rect 41417 12733 41429 12767
rect 41463 12733 41475 12767
rect 41417 12727 41475 12733
rect 37476 12600 40080 12628
rect 40126 12588 40132 12640
rect 40184 12628 40190 12640
rect 40954 12628 40960 12640
rect 40184 12600 40960 12628
rect 40184 12588 40190 12600
rect 40954 12588 40960 12600
rect 41012 12628 41018 12640
rect 41432 12628 41460 12727
rect 41690 12724 41696 12776
rect 41748 12764 41754 12776
rect 41785 12767 41843 12773
rect 41785 12764 41797 12767
rect 41748 12736 41797 12764
rect 41748 12724 41754 12736
rect 41785 12733 41797 12736
rect 41831 12733 41843 12767
rect 41785 12727 41843 12733
rect 41874 12724 41880 12776
rect 41932 12724 41938 12776
rect 41598 12628 41604 12640
rect 41012 12600 41604 12628
rect 41012 12588 41018 12600
rect 41598 12588 41604 12600
rect 41656 12588 41662 12640
rect 44361 12631 44419 12637
rect 44361 12597 44373 12631
rect 44407 12628 44419 12631
rect 45002 12628 45008 12640
rect 44407 12600 45008 12628
rect 44407 12597 44419 12600
rect 44361 12591 44419 12597
rect 45002 12588 45008 12600
rect 45060 12588 45066 12640
rect 1104 12538 44896 12560
rect 1104 12486 6423 12538
rect 6475 12486 6487 12538
rect 6539 12486 6551 12538
rect 6603 12486 6615 12538
rect 6667 12486 6679 12538
rect 6731 12486 17370 12538
rect 17422 12486 17434 12538
rect 17486 12486 17498 12538
rect 17550 12486 17562 12538
rect 17614 12486 17626 12538
rect 17678 12486 28317 12538
rect 28369 12486 28381 12538
rect 28433 12486 28445 12538
rect 28497 12486 28509 12538
rect 28561 12486 28573 12538
rect 28625 12486 39264 12538
rect 39316 12486 39328 12538
rect 39380 12486 39392 12538
rect 39444 12486 39456 12538
rect 39508 12486 39520 12538
rect 39572 12486 44896 12538
rect 1104 12464 44896 12486
rect 2958 12384 2964 12436
rect 3016 12384 3022 12436
rect 7374 12384 7380 12436
rect 7432 12384 7438 12436
rect 10042 12384 10048 12436
rect 10100 12424 10106 12436
rect 10137 12427 10195 12433
rect 10137 12424 10149 12427
rect 10100 12396 10149 12424
rect 10100 12384 10106 12396
rect 10137 12393 10149 12396
rect 10183 12393 10195 12427
rect 10137 12387 10195 12393
rect 11054 12384 11060 12436
rect 11112 12424 11118 12436
rect 11112 12396 11744 12424
rect 11112 12384 11118 12396
rect 11716 12356 11744 12396
rect 11790 12384 11796 12436
rect 11848 12424 11854 12436
rect 12161 12427 12219 12433
rect 12161 12424 12173 12427
rect 11848 12396 12173 12424
rect 11848 12384 11854 12396
rect 12161 12393 12173 12396
rect 12207 12393 12219 12427
rect 12161 12387 12219 12393
rect 12989 12427 13047 12433
rect 12989 12393 13001 12427
rect 13035 12424 13047 12427
rect 13814 12424 13820 12436
rect 13035 12396 13820 12424
rect 13035 12393 13047 12396
rect 12989 12387 13047 12393
rect 13814 12384 13820 12396
rect 13872 12384 13878 12436
rect 20714 12384 20720 12436
rect 20772 12424 20778 12436
rect 21177 12427 21235 12433
rect 21177 12424 21189 12427
rect 20772 12396 21189 12424
rect 20772 12384 20778 12396
rect 21177 12393 21189 12396
rect 21223 12424 21235 12427
rect 21910 12424 21916 12436
rect 21223 12396 21916 12424
rect 21223 12393 21235 12396
rect 21177 12387 21235 12393
rect 21910 12384 21916 12396
rect 21968 12384 21974 12436
rect 25866 12424 25872 12436
rect 22020 12396 25872 12424
rect 11716 12328 11836 12356
rect 4893 12291 4951 12297
rect 4893 12257 4905 12291
rect 4939 12288 4951 12291
rect 8021 12291 8079 12297
rect 4939 12260 5580 12288
rect 4939 12257 4951 12260
rect 4893 12251 4951 12257
rect 3145 12223 3203 12229
rect 3145 12189 3157 12223
rect 3191 12220 3203 12223
rect 3418 12220 3424 12232
rect 3191 12192 3424 12220
rect 3191 12189 3203 12192
rect 3145 12183 3203 12189
rect 3418 12180 3424 12192
rect 3476 12180 3482 12232
rect 5074 12180 5080 12232
rect 5132 12220 5138 12232
rect 5445 12223 5503 12229
rect 5445 12220 5457 12223
rect 5132 12192 5457 12220
rect 5132 12180 5138 12192
rect 5445 12189 5457 12192
rect 5491 12189 5503 12223
rect 5552 12220 5580 12260
rect 8021 12257 8033 12291
rect 8067 12288 8079 12291
rect 9674 12288 9680 12300
rect 8067 12260 9680 12288
rect 8067 12257 8079 12260
rect 8021 12251 8079 12257
rect 9674 12248 9680 12260
rect 9732 12248 9738 12300
rect 11808 12288 11836 12328
rect 12342 12316 12348 12368
rect 12400 12356 12406 12368
rect 12400 12328 15240 12356
rect 12400 12316 12406 12328
rect 15212 12297 15240 12328
rect 20898 12316 20904 12368
rect 20956 12356 20962 12368
rect 20956 12328 21864 12356
rect 20956 12316 20962 12328
rect 13633 12291 13691 12297
rect 13633 12288 13645 12291
rect 11808 12260 13645 12288
rect 13633 12257 13645 12260
rect 13679 12288 13691 12291
rect 15197 12291 15255 12297
rect 13679 12260 15148 12288
rect 13679 12257 13691 12260
rect 13633 12251 13691 12257
rect 7558 12220 7564 12232
rect 5552 12192 7564 12220
rect 5445 12183 5503 12189
rect 7558 12180 7564 12192
rect 7616 12180 7622 12232
rect 7742 12180 7748 12232
rect 7800 12180 7806 12232
rect 10318 12180 10324 12232
rect 10376 12180 10382 12232
rect 10781 12223 10839 12229
rect 10781 12189 10793 12223
rect 10827 12220 10839 12223
rect 11422 12220 11428 12232
rect 10827 12192 11428 12220
rect 10827 12189 10839 12192
rect 10781 12183 10839 12189
rect 11422 12180 11428 12192
rect 11480 12180 11486 12232
rect 14550 12180 14556 12232
rect 14608 12220 14614 12232
rect 15013 12223 15071 12229
rect 15013 12220 15025 12223
rect 14608 12192 15025 12220
rect 14608 12180 14614 12192
rect 15013 12189 15025 12192
rect 15059 12189 15071 12223
rect 15120 12220 15148 12260
rect 15197 12257 15209 12291
rect 15243 12288 15255 12291
rect 17218 12288 17224 12300
rect 15243 12260 17224 12288
rect 15243 12257 15255 12260
rect 15197 12251 15255 12257
rect 17218 12248 17224 12260
rect 17276 12248 17282 12300
rect 18506 12248 18512 12300
rect 18564 12288 18570 12300
rect 19429 12291 19487 12297
rect 19429 12288 19441 12291
rect 18564 12260 19441 12288
rect 18564 12248 18570 12260
rect 19429 12257 19441 12260
rect 19475 12257 19487 12291
rect 19429 12251 19487 12257
rect 19705 12291 19763 12297
rect 19705 12257 19717 12291
rect 19751 12288 19763 12291
rect 21637 12291 21695 12297
rect 21637 12288 21649 12291
rect 19751 12260 21649 12288
rect 19751 12257 19763 12260
rect 19705 12251 19763 12257
rect 21637 12257 21649 12260
rect 21683 12257 21695 12291
rect 21637 12251 21695 12257
rect 21836 12232 21864 12328
rect 17494 12220 17500 12232
rect 15120 12192 17500 12220
rect 15013 12183 15071 12189
rect 17494 12180 17500 12192
rect 17552 12180 17558 12232
rect 17954 12180 17960 12232
rect 18012 12220 18018 12232
rect 18690 12220 18696 12232
rect 18012 12192 18696 12220
rect 18012 12180 18018 12192
rect 18690 12180 18696 12192
rect 18748 12180 18754 12232
rect 21818 12180 21824 12232
rect 21876 12180 21882 12232
rect 22020 12229 22048 12396
rect 22094 12248 22100 12300
rect 22152 12288 22158 12300
rect 22281 12291 22339 12297
rect 22281 12288 22293 12291
rect 22152 12260 22293 12288
rect 22152 12248 22158 12260
rect 22281 12257 22293 12260
rect 22327 12257 22339 12291
rect 22281 12251 22339 12257
rect 22756 12229 22784 12396
rect 25866 12384 25872 12396
rect 25924 12384 25930 12436
rect 26878 12384 26884 12436
rect 26936 12384 26942 12436
rect 31202 12384 31208 12436
rect 31260 12424 31266 12436
rect 32953 12427 33011 12433
rect 32953 12424 32965 12427
rect 31260 12396 32965 12424
rect 31260 12384 31266 12396
rect 32953 12393 32965 12396
rect 32999 12424 33011 12427
rect 33318 12424 33324 12436
rect 32999 12396 33324 12424
rect 32999 12393 33011 12396
rect 32953 12387 33011 12393
rect 33318 12384 33324 12396
rect 33376 12384 33382 12436
rect 35342 12384 35348 12436
rect 35400 12424 35406 12436
rect 35437 12427 35495 12433
rect 35437 12424 35449 12427
rect 35400 12396 35449 12424
rect 35400 12384 35406 12396
rect 35437 12393 35449 12396
rect 35483 12393 35495 12427
rect 35437 12387 35495 12393
rect 35526 12384 35532 12436
rect 35584 12424 35590 12436
rect 35584 12396 36216 12424
rect 35584 12384 35590 12396
rect 29546 12316 29552 12368
rect 29604 12356 29610 12368
rect 31021 12359 31079 12365
rect 31021 12356 31033 12359
rect 29604 12328 31033 12356
rect 29604 12316 29610 12328
rect 31021 12325 31033 12328
rect 31067 12325 31079 12359
rect 31021 12319 31079 12325
rect 31754 12316 31760 12368
rect 31812 12356 31818 12368
rect 33042 12356 33048 12368
rect 31812 12328 33048 12356
rect 31812 12316 31818 12328
rect 24578 12248 24584 12300
rect 24636 12288 24642 12300
rect 24854 12288 24860 12300
rect 24636 12260 24860 12288
rect 24636 12248 24642 12260
rect 24854 12248 24860 12260
rect 24912 12288 24918 12300
rect 26510 12288 26516 12300
rect 24912 12260 26516 12288
rect 24912 12248 24918 12260
rect 26510 12248 26516 12260
rect 26568 12248 26574 12300
rect 28902 12248 28908 12300
rect 28960 12288 28966 12300
rect 30009 12291 30067 12297
rect 30009 12288 30021 12291
rect 28960 12260 30021 12288
rect 28960 12248 28966 12260
rect 30009 12257 30021 12260
rect 30055 12257 30067 12291
rect 32122 12288 32128 12300
rect 30009 12251 30067 12257
rect 31772 12260 32128 12288
rect 31772 12232 31800 12260
rect 32122 12248 32128 12260
rect 32180 12248 32186 12300
rect 22005 12223 22063 12229
rect 22005 12189 22017 12223
rect 22051 12189 22063 12223
rect 22005 12183 22063 12189
rect 22741 12223 22799 12229
rect 22741 12189 22753 12223
rect 22787 12189 22799 12223
rect 23017 12223 23075 12229
rect 23017 12220 23029 12223
rect 22741 12183 22799 12189
rect 22848 12192 23029 12220
rect 5712 12155 5770 12161
rect 5712 12121 5724 12155
rect 5758 12152 5770 12155
rect 5994 12152 6000 12164
rect 5758 12124 6000 12152
rect 5758 12121 5770 12124
rect 5712 12115 5770 12121
rect 5994 12112 6000 12124
rect 6052 12112 6058 12164
rect 8202 12152 8208 12164
rect 6748 12124 8208 12152
rect 4246 12044 4252 12096
rect 4304 12044 4310 12096
rect 4614 12044 4620 12096
rect 4672 12044 4678 12096
rect 4709 12087 4767 12093
rect 4709 12053 4721 12087
rect 4755 12084 4767 12087
rect 6748 12084 6776 12124
rect 8202 12112 8208 12124
rect 8260 12112 8266 12164
rect 11048 12155 11106 12161
rect 11048 12121 11060 12155
rect 11094 12152 11106 12155
rect 12434 12152 12440 12164
rect 11094 12124 12440 12152
rect 11094 12121 11106 12124
rect 11048 12115 11106 12121
rect 12434 12112 12440 12124
rect 12492 12112 12498 12164
rect 19812 12124 20194 12152
rect 4755 12056 6776 12084
rect 6825 12087 6883 12093
rect 4755 12053 4767 12056
rect 4709 12047 4767 12053
rect 6825 12053 6837 12087
rect 6871 12084 6883 12087
rect 7374 12084 7380 12096
rect 6871 12056 7380 12084
rect 6871 12053 6883 12056
rect 6825 12047 6883 12053
rect 7374 12044 7380 12056
rect 7432 12044 7438 12096
rect 7837 12087 7895 12093
rect 7837 12053 7849 12087
rect 7883 12084 7895 12087
rect 11146 12084 11152 12096
rect 7883 12056 11152 12084
rect 7883 12053 7895 12056
rect 7837 12047 7895 12053
rect 11146 12044 11152 12056
rect 11204 12044 11210 12096
rect 13354 12044 13360 12096
rect 13412 12044 13418 12096
rect 13449 12087 13507 12093
rect 13449 12053 13461 12087
rect 13495 12084 13507 12087
rect 14645 12087 14703 12093
rect 14645 12084 14657 12087
rect 13495 12056 14657 12084
rect 13495 12053 13507 12056
rect 13449 12047 13507 12053
rect 14645 12053 14657 12056
rect 14691 12053 14703 12087
rect 14645 12047 14703 12053
rect 15105 12087 15163 12093
rect 15105 12053 15117 12087
rect 15151 12084 15163 12087
rect 17126 12084 17132 12096
rect 15151 12056 17132 12084
rect 15151 12053 15163 12056
rect 15105 12047 15163 12053
rect 17126 12044 17132 12056
rect 17184 12044 17190 12096
rect 18785 12087 18843 12093
rect 18785 12053 18797 12087
rect 18831 12084 18843 12087
rect 19812 12084 19840 12124
rect 21910 12112 21916 12164
rect 21968 12112 21974 12164
rect 22094 12112 22100 12164
rect 22152 12161 22158 12164
rect 22152 12155 22181 12161
rect 22169 12121 22181 12155
rect 22848 12152 22876 12192
rect 23017 12189 23029 12192
rect 23063 12189 23075 12223
rect 23017 12183 23075 12189
rect 23106 12180 23112 12232
rect 23164 12180 23170 12232
rect 26142 12180 26148 12232
rect 26200 12220 26206 12232
rect 26789 12223 26847 12229
rect 26789 12220 26801 12223
rect 26200 12192 26801 12220
rect 26200 12180 26206 12192
rect 26789 12189 26801 12192
rect 26835 12189 26847 12223
rect 26789 12183 26847 12189
rect 29730 12180 29736 12232
rect 29788 12180 29794 12232
rect 31297 12223 31355 12229
rect 31297 12220 31309 12223
rect 30392 12192 31309 12220
rect 22152 12115 22181 12121
rect 22572 12124 22876 12152
rect 22925 12155 22983 12161
rect 22152 12112 22158 12115
rect 18831 12056 19840 12084
rect 18831 12053 18843 12056
rect 18785 12047 18843 12053
rect 21450 12044 21456 12096
rect 21508 12084 21514 12096
rect 22572 12084 22600 12124
rect 22925 12121 22937 12155
rect 22971 12121 22983 12155
rect 24857 12155 24915 12161
rect 24857 12152 24869 12155
rect 22925 12115 22983 12121
rect 23308 12124 24869 12152
rect 21508 12056 22600 12084
rect 21508 12044 21514 12056
rect 22738 12044 22744 12096
rect 22796 12084 22802 12096
rect 22940 12084 22968 12115
rect 23308 12093 23336 12124
rect 24857 12121 24869 12124
rect 24903 12121 24915 12155
rect 24857 12115 24915 12121
rect 25498 12112 25504 12164
rect 25556 12112 25562 12164
rect 29638 12112 29644 12164
rect 29696 12152 29702 12164
rect 30392 12152 30420 12192
rect 31297 12189 31309 12192
rect 31343 12189 31355 12223
rect 31297 12183 31355 12189
rect 29696 12124 30420 12152
rect 29696 12112 29702 12124
rect 30926 12112 30932 12164
rect 30984 12152 30990 12164
rect 31021 12155 31079 12161
rect 31021 12152 31033 12155
rect 30984 12124 31033 12152
rect 30984 12112 30990 12124
rect 31021 12121 31033 12124
rect 31067 12121 31079 12155
rect 31021 12115 31079 12121
rect 22796 12056 22968 12084
rect 23293 12087 23351 12093
rect 22796 12044 22802 12056
rect 23293 12053 23305 12087
rect 23339 12053 23351 12087
rect 23293 12047 23351 12053
rect 25130 12044 25136 12096
rect 25188 12084 25194 12096
rect 26329 12087 26387 12093
rect 26329 12084 26341 12087
rect 25188 12056 26341 12084
rect 25188 12044 25194 12056
rect 26329 12053 26341 12056
rect 26375 12053 26387 12087
rect 26329 12047 26387 12053
rect 31202 12044 31208 12096
rect 31260 12044 31266 12096
rect 31312 12084 31340 12183
rect 31754 12180 31760 12232
rect 31812 12180 31818 12232
rect 31938 12180 31944 12232
rect 31996 12180 32002 12232
rect 32033 12223 32091 12229
rect 32033 12189 32045 12223
rect 32079 12220 32091 12223
rect 32232 12220 32260 12328
rect 33042 12316 33048 12328
rect 33100 12316 33106 12368
rect 35250 12316 35256 12368
rect 35308 12356 35314 12368
rect 35802 12356 35808 12368
rect 35308 12328 35808 12356
rect 35308 12316 35314 12328
rect 35802 12316 35808 12328
rect 35860 12356 35866 12368
rect 35860 12328 36124 12356
rect 35860 12316 35866 12328
rect 32490 12248 32496 12300
rect 32548 12288 32554 12300
rect 35986 12288 35992 12300
rect 32548 12260 35992 12288
rect 32548 12248 32554 12260
rect 32079 12192 32260 12220
rect 32309 12223 32367 12229
rect 32079 12189 32091 12192
rect 32033 12183 32091 12189
rect 32309 12189 32321 12223
rect 32355 12220 32367 12223
rect 33226 12220 33232 12232
rect 32355 12192 33232 12220
rect 32355 12189 32367 12192
rect 32309 12183 32367 12189
rect 32122 12112 32128 12164
rect 32180 12112 32186 12164
rect 32324 12084 32352 12183
rect 33226 12180 33232 12192
rect 33284 12180 33290 12232
rect 34072 12229 34100 12260
rect 35986 12248 35992 12260
rect 36044 12248 36050 12300
rect 36096 12297 36124 12328
rect 36081 12291 36139 12297
rect 36081 12257 36093 12291
rect 36127 12257 36139 12291
rect 36188 12288 36216 12396
rect 36262 12384 36268 12436
rect 36320 12424 36326 12436
rect 36449 12427 36507 12433
rect 36449 12424 36461 12427
rect 36320 12396 36461 12424
rect 36320 12384 36326 12396
rect 36449 12393 36461 12396
rect 36495 12393 36507 12427
rect 36449 12387 36507 12393
rect 36909 12427 36967 12433
rect 36909 12393 36921 12427
rect 36955 12424 36967 12427
rect 37918 12424 37924 12436
rect 36955 12396 37924 12424
rect 36955 12393 36967 12396
rect 36909 12387 36967 12393
rect 37918 12384 37924 12396
rect 37976 12384 37982 12436
rect 38120 12396 40632 12424
rect 38010 12356 38016 12368
rect 37200 12328 38016 12356
rect 37200 12288 37228 12328
rect 38010 12316 38016 12328
rect 38068 12316 38074 12368
rect 38120 12288 38148 12396
rect 38654 12316 38660 12368
rect 38712 12356 38718 12368
rect 39206 12356 39212 12368
rect 38712 12328 39212 12356
rect 38712 12316 38718 12328
rect 39206 12316 39212 12328
rect 39264 12316 39270 12368
rect 40218 12316 40224 12368
rect 40276 12356 40282 12368
rect 40276 12328 40540 12356
rect 40276 12316 40282 12328
rect 40034 12288 40040 12300
rect 36188 12260 37228 12288
rect 36081 12251 36139 12257
rect 34057 12223 34115 12229
rect 34057 12189 34069 12223
rect 34103 12189 34115 12223
rect 34057 12183 34115 12189
rect 35176 12192 36032 12220
rect 32766 12112 32772 12164
rect 32824 12112 32830 12164
rect 32985 12155 33043 12161
rect 32985 12121 32997 12155
rect 33031 12152 33043 12155
rect 35176 12152 35204 12192
rect 33031 12124 35204 12152
rect 33031 12121 33043 12124
rect 32985 12115 33043 12121
rect 35250 12112 35256 12164
rect 35308 12112 35314 12164
rect 35469 12155 35527 12161
rect 35469 12121 35481 12155
rect 35515 12152 35527 12155
rect 35710 12152 35716 12164
rect 35515 12124 35716 12152
rect 35515 12121 35527 12124
rect 35469 12115 35527 12121
rect 35710 12112 35716 12124
rect 35768 12112 35774 12164
rect 31312 12056 32352 12084
rect 33134 12044 33140 12096
rect 33192 12044 33198 12096
rect 34241 12087 34299 12093
rect 34241 12053 34253 12087
rect 34287 12084 34299 12087
rect 35158 12084 35164 12096
rect 34287 12056 35164 12084
rect 34287 12053 34299 12056
rect 34241 12047 34299 12053
rect 35158 12044 35164 12056
rect 35216 12044 35222 12096
rect 35618 12044 35624 12096
rect 35676 12044 35682 12096
rect 36004 12084 36032 12192
rect 36096 12152 36124 12251
rect 36170 12180 36176 12232
rect 36228 12220 36234 12232
rect 36265 12223 36323 12229
rect 36265 12220 36277 12223
rect 36228 12192 36277 12220
rect 36228 12180 36234 12192
rect 36265 12189 36277 12192
rect 36311 12220 36323 12223
rect 36630 12220 36636 12232
rect 36311 12192 36636 12220
rect 36311 12189 36323 12192
rect 36265 12183 36323 12189
rect 36630 12180 36636 12192
rect 36688 12180 36694 12232
rect 37200 12229 37228 12260
rect 37476 12260 38148 12288
rect 38948 12260 40040 12288
rect 37185 12223 37243 12229
rect 37185 12189 37197 12223
rect 37231 12189 37243 12223
rect 37185 12183 37243 12189
rect 37274 12180 37280 12232
rect 37332 12180 37338 12232
rect 37366 12180 37372 12232
rect 37424 12180 37430 12232
rect 37476 12152 37504 12260
rect 37553 12223 37611 12229
rect 37553 12189 37565 12223
rect 37599 12220 37611 12223
rect 37918 12220 37924 12232
rect 37599 12192 37924 12220
rect 37599 12189 37611 12192
rect 37553 12183 37611 12189
rect 37918 12180 37924 12192
rect 37976 12180 37982 12232
rect 38013 12223 38071 12229
rect 38013 12189 38025 12223
rect 38059 12189 38071 12223
rect 38013 12183 38071 12189
rect 36096 12124 37504 12152
rect 37734 12112 37740 12164
rect 37792 12152 37798 12164
rect 38028 12152 38056 12183
rect 38102 12180 38108 12232
rect 38160 12220 38166 12232
rect 38197 12223 38255 12229
rect 38197 12220 38209 12223
rect 38160 12192 38209 12220
rect 38160 12180 38166 12192
rect 38197 12189 38209 12192
rect 38243 12220 38255 12223
rect 38746 12220 38752 12232
rect 38243 12192 38752 12220
rect 38243 12189 38255 12192
rect 38197 12183 38255 12189
rect 38746 12180 38752 12192
rect 38804 12180 38810 12232
rect 38948 12229 38976 12260
rect 40034 12248 40040 12260
rect 40092 12288 40098 12300
rect 40402 12288 40408 12300
rect 40092 12260 40408 12288
rect 40092 12248 40098 12260
rect 40402 12248 40408 12260
rect 40460 12248 40466 12300
rect 40512 12297 40540 12328
rect 40497 12291 40555 12297
rect 40497 12257 40509 12291
rect 40543 12257 40555 12291
rect 40604 12288 40632 12396
rect 40706 12291 40764 12297
rect 40706 12288 40718 12291
rect 40604 12260 40718 12288
rect 40497 12251 40555 12257
rect 40706 12257 40718 12260
rect 40752 12257 40764 12291
rect 41690 12288 41696 12300
rect 40706 12251 40764 12257
rect 40880 12260 41696 12288
rect 38841 12223 38899 12229
rect 38841 12189 38853 12223
rect 38887 12189 38899 12223
rect 38841 12183 38899 12189
rect 38933 12223 38991 12229
rect 38933 12189 38945 12223
rect 38979 12189 38991 12223
rect 38933 12183 38991 12189
rect 38654 12152 38660 12164
rect 37792 12124 38660 12152
rect 37792 12112 37798 12124
rect 38654 12112 38660 12124
rect 38712 12112 38718 12164
rect 38856 12152 38884 12183
rect 39114 12180 39120 12232
rect 39172 12180 39178 12232
rect 39206 12180 39212 12232
rect 39264 12180 39270 12232
rect 39301 12223 39359 12229
rect 39301 12189 39313 12223
rect 39347 12189 39359 12223
rect 39301 12183 39359 12189
rect 40221 12223 40279 12229
rect 40221 12189 40233 12223
rect 40267 12189 40279 12223
rect 40880 12220 40908 12260
rect 41690 12248 41696 12260
rect 41748 12248 41754 12300
rect 40221 12183 40279 12189
rect 40696 12192 40908 12220
rect 39022 12152 39028 12164
rect 38856 12124 39028 12152
rect 39022 12112 39028 12124
rect 39080 12112 39086 12164
rect 39316 12152 39344 12183
rect 39132 12124 39344 12152
rect 39132 12096 39160 12124
rect 38102 12084 38108 12096
rect 36004 12056 38108 12084
rect 38102 12044 38108 12056
rect 38160 12044 38166 12096
rect 38378 12044 38384 12096
rect 38436 12044 38442 12096
rect 38838 12044 38844 12096
rect 38896 12044 38902 12096
rect 39114 12044 39120 12096
rect 39172 12044 39178 12096
rect 40236 12084 40264 12183
rect 40310 12112 40316 12164
rect 40368 12152 40374 12164
rect 40589 12155 40647 12161
rect 40589 12152 40601 12155
rect 40368 12124 40601 12152
rect 40368 12112 40374 12124
rect 40589 12121 40601 12124
rect 40635 12152 40647 12155
rect 40696 12152 40724 12192
rect 41414 12180 41420 12232
rect 41472 12220 41478 12232
rect 41785 12223 41843 12229
rect 41785 12220 41797 12223
rect 41472 12192 41797 12220
rect 41472 12180 41478 12192
rect 41785 12189 41797 12192
rect 41831 12189 41843 12223
rect 41785 12183 41843 12189
rect 41966 12180 41972 12232
rect 42024 12220 42030 12232
rect 42061 12223 42119 12229
rect 42061 12220 42073 12223
rect 42024 12192 42073 12220
rect 42024 12180 42030 12192
rect 42061 12189 42073 12192
rect 42107 12189 42119 12223
rect 42061 12183 42119 12189
rect 42242 12180 42248 12232
rect 42300 12180 42306 12232
rect 41506 12152 41512 12164
rect 40635 12124 40724 12152
rect 40788 12124 41512 12152
rect 40635 12121 40647 12124
rect 40589 12115 40647 12121
rect 40788 12084 40816 12124
rect 41506 12112 41512 12124
rect 41564 12112 41570 12164
rect 40236 12056 40816 12084
rect 40862 12044 40868 12096
rect 40920 12044 40926 12096
rect 41601 12087 41659 12093
rect 41601 12053 41613 12087
rect 41647 12084 41659 12087
rect 41690 12084 41696 12096
rect 41647 12056 41696 12084
rect 41647 12053 41659 12056
rect 41601 12047 41659 12053
rect 41690 12044 41696 12056
rect 41748 12044 41754 12096
rect 1104 11994 45051 12016
rect 1104 11942 11896 11994
rect 11948 11942 11960 11994
rect 12012 11942 12024 11994
rect 12076 11942 12088 11994
rect 12140 11942 12152 11994
rect 12204 11942 22843 11994
rect 22895 11942 22907 11994
rect 22959 11942 22971 11994
rect 23023 11942 23035 11994
rect 23087 11942 23099 11994
rect 23151 11942 33790 11994
rect 33842 11942 33854 11994
rect 33906 11942 33918 11994
rect 33970 11942 33982 11994
rect 34034 11942 34046 11994
rect 34098 11942 44737 11994
rect 44789 11942 44801 11994
rect 44853 11942 44865 11994
rect 44917 11942 44929 11994
rect 44981 11942 44993 11994
rect 45045 11942 45051 11994
rect 1104 11920 45051 11942
rect 3973 11883 4031 11889
rect 3973 11849 3985 11883
rect 4019 11880 4031 11883
rect 5997 11883 6055 11889
rect 4019 11852 5212 11880
rect 4019 11849 4031 11852
rect 3973 11843 4031 11849
rect 4522 11812 4528 11824
rect 3436 11784 4528 11812
rect 3436 11753 3464 11784
rect 4522 11772 4528 11784
rect 4580 11772 4586 11824
rect 5074 11812 5080 11824
rect 4632 11784 5080 11812
rect 3421 11747 3479 11753
rect 3421 11713 3433 11747
rect 3467 11713 3479 11747
rect 3421 11707 3479 11713
rect 4157 11747 4215 11753
rect 4157 11713 4169 11747
rect 4203 11744 4215 11747
rect 4246 11744 4252 11756
rect 4203 11716 4252 11744
rect 4203 11713 4215 11716
rect 4157 11707 4215 11713
rect 4246 11704 4252 11716
rect 4304 11704 4310 11756
rect 4632 11685 4660 11784
rect 5074 11772 5080 11784
rect 5132 11772 5138 11824
rect 4884 11747 4942 11753
rect 4884 11713 4896 11747
rect 4930 11744 4942 11747
rect 5184 11744 5212 11852
rect 5997 11849 6009 11883
rect 6043 11849 6055 11883
rect 5997 11843 6055 11849
rect 4930 11716 5212 11744
rect 6012 11744 6040 11843
rect 7374 11840 7380 11892
rect 7432 11840 7438 11892
rect 7469 11883 7527 11889
rect 7469 11849 7481 11883
rect 7515 11880 7527 11883
rect 7742 11880 7748 11892
rect 7515 11852 7748 11880
rect 7515 11849 7527 11852
rect 7469 11843 7527 11849
rect 7742 11840 7748 11852
rect 7800 11840 7806 11892
rect 8202 11840 8208 11892
rect 8260 11840 8266 11892
rect 13354 11840 13360 11892
rect 13412 11880 13418 11892
rect 14553 11883 14611 11889
rect 14553 11880 14565 11883
rect 13412 11852 14565 11880
rect 13412 11840 13418 11852
rect 14553 11849 14565 11852
rect 14599 11849 14611 11883
rect 14553 11843 14611 11849
rect 15013 11883 15071 11889
rect 15013 11849 15025 11883
rect 15059 11849 15071 11883
rect 15013 11843 15071 11849
rect 19705 11883 19763 11889
rect 19705 11849 19717 11883
rect 19751 11849 19763 11883
rect 19705 11843 19763 11849
rect 7392 11812 7420 11840
rect 8665 11815 8723 11821
rect 8665 11812 8677 11815
rect 7392 11784 8677 11812
rect 8665 11781 8677 11784
rect 8711 11781 8723 11815
rect 10778 11812 10784 11824
rect 8665 11775 8723 11781
rect 10244 11784 10784 11812
rect 8573 11747 8631 11753
rect 8573 11744 8585 11747
rect 6012 11716 8585 11744
rect 4930 11713 4942 11716
rect 4884 11707 4942 11713
rect 8573 11713 8585 11716
rect 8619 11744 8631 11747
rect 10244 11744 10272 11784
rect 10778 11772 10784 11784
rect 10836 11772 10842 11824
rect 13440 11815 13498 11821
rect 13440 11781 13452 11815
rect 13486 11812 13498 11815
rect 15028 11812 15056 11843
rect 13486 11784 15056 11812
rect 13486 11781 13498 11784
rect 13440 11775 13498 11781
rect 8619 11716 10272 11744
rect 8619 11713 8631 11716
rect 8573 11707 8631 11713
rect 10318 11704 10324 11756
rect 10376 11704 10382 11756
rect 12894 11704 12900 11756
rect 12952 11744 12958 11756
rect 13170 11744 13176 11756
rect 12952 11716 13176 11744
rect 12952 11704 12958 11716
rect 13170 11704 13176 11716
rect 13228 11704 13234 11756
rect 14642 11704 14648 11756
rect 14700 11744 14706 11756
rect 15197 11747 15255 11753
rect 15197 11744 15209 11747
rect 14700 11716 15209 11744
rect 14700 11704 14706 11716
rect 15197 11713 15209 11716
rect 15243 11713 15255 11747
rect 15197 11707 15255 11713
rect 16390 11704 16396 11756
rect 16448 11744 16454 11756
rect 17221 11747 17279 11753
rect 17221 11744 17233 11747
rect 16448 11716 17233 11744
rect 16448 11704 16454 11716
rect 17221 11713 17233 11716
rect 17267 11713 17279 11747
rect 17221 11707 17279 11713
rect 19245 11747 19303 11753
rect 19245 11713 19257 11747
rect 19291 11744 19303 11747
rect 19720 11744 19748 11843
rect 19978 11840 19984 11892
rect 20036 11880 20042 11892
rect 20073 11883 20131 11889
rect 20073 11880 20085 11883
rect 20036 11852 20085 11880
rect 20036 11840 20042 11852
rect 20073 11849 20085 11852
rect 20119 11849 20131 11883
rect 20073 11843 20131 11849
rect 22738 11840 22744 11892
rect 22796 11880 22802 11892
rect 22925 11883 22983 11889
rect 22925 11880 22937 11883
rect 22796 11852 22937 11880
rect 22796 11840 22802 11852
rect 22925 11849 22937 11852
rect 22971 11849 22983 11883
rect 22925 11843 22983 11849
rect 25866 11840 25872 11892
rect 25924 11880 25930 11892
rect 26605 11883 26663 11889
rect 26605 11880 26617 11883
rect 25924 11852 26617 11880
rect 25924 11840 25930 11852
rect 26605 11849 26617 11852
rect 26651 11849 26663 11883
rect 26605 11843 26663 11849
rect 29365 11883 29423 11889
rect 29365 11849 29377 11883
rect 29411 11880 29423 11883
rect 29454 11880 29460 11892
rect 29411 11852 29460 11880
rect 29411 11849 29423 11852
rect 29365 11843 29423 11849
rect 29454 11840 29460 11852
rect 29512 11840 29518 11892
rect 29730 11840 29736 11892
rect 29788 11880 29794 11892
rect 32677 11883 32735 11889
rect 32677 11880 32689 11883
rect 29788 11852 32689 11880
rect 29788 11840 29794 11852
rect 32677 11849 32689 11852
rect 32723 11849 32735 11883
rect 32677 11843 32735 11849
rect 33502 11840 33508 11892
rect 33560 11840 33566 11892
rect 35434 11840 35440 11892
rect 35492 11880 35498 11892
rect 36538 11880 36544 11892
rect 35492 11852 36544 11880
rect 35492 11840 35498 11852
rect 36538 11840 36544 11852
rect 36596 11840 36602 11892
rect 36630 11840 36636 11892
rect 36688 11880 36694 11892
rect 37550 11880 37556 11892
rect 36688 11852 37556 11880
rect 36688 11840 36694 11852
rect 37550 11840 37556 11852
rect 37608 11840 37614 11892
rect 37642 11840 37648 11892
rect 37700 11880 37706 11892
rect 37829 11883 37887 11889
rect 37829 11880 37841 11883
rect 37700 11852 37841 11880
rect 37700 11840 37706 11852
rect 37829 11849 37841 11852
rect 37875 11849 37887 11883
rect 37829 11843 37887 11849
rect 38102 11840 38108 11892
rect 38160 11840 38166 11892
rect 38562 11840 38568 11892
rect 38620 11840 38626 11892
rect 38930 11840 38936 11892
rect 38988 11840 38994 11892
rect 41414 11840 41420 11892
rect 41472 11840 41478 11892
rect 20165 11815 20223 11821
rect 20165 11781 20177 11815
rect 20211 11812 20223 11815
rect 20211 11784 21496 11812
rect 20211 11781 20223 11784
rect 20165 11775 20223 11781
rect 21468 11756 21496 11784
rect 21910 11772 21916 11824
rect 21968 11812 21974 11824
rect 25038 11812 25044 11824
rect 21968 11784 25044 11812
rect 21968 11772 21974 11784
rect 19291 11716 19748 11744
rect 19291 11713 19303 11716
rect 19245 11707 19303 11713
rect 20990 11704 20996 11756
rect 21048 11744 21054 11756
rect 21361 11747 21419 11753
rect 21361 11744 21373 11747
rect 21048 11716 21373 11744
rect 21048 11704 21054 11716
rect 21361 11713 21373 11716
rect 21407 11713 21419 11747
rect 21361 11707 21419 11713
rect 21450 11704 21456 11756
rect 21508 11704 21514 11756
rect 22094 11704 22100 11756
rect 22152 11704 22158 11756
rect 22189 11747 22247 11753
rect 22189 11713 22201 11747
rect 22235 11744 22247 11747
rect 22278 11744 22284 11756
rect 22235 11716 22284 11744
rect 22235 11713 22247 11716
rect 22189 11707 22247 11713
rect 22278 11704 22284 11716
rect 22336 11704 22342 11756
rect 22830 11704 22836 11756
rect 22888 11704 22894 11756
rect 23032 11753 23060 11784
rect 25038 11772 25044 11784
rect 25096 11772 25102 11824
rect 25130 11772 25136 11824
rect 25188 11772 25194 11824
rect 28813 11815 28871 11821
rect 28813 11781 28825 11815
rect 28859 11812 28871 11815
rect 30650 11812 30656 11824
rect 28859 11784 30656 11812
rect 28859 11781 28871 11784
rect 28813 11775 28871 11781
rect 23017 11747 23075 11753
rect 23017 11713 23029 11747
rect 23063 11713 23075 11747
rect 23017 11707 23075 11713
rect 26142 11704 26148 11756
rect 26200 11744 26206 11756
rect 28629 11747 28687 11753
rect 26200 11716 26266 11744
rect 26200 11704 26206 11716
rect 28629 11713 28641 11747
rect 28675 11713 28687 11747
rect 28629 11707 28687 11713
rect 28905 11747 28963 11753
rect 28905 11713 28917 11747
rect 28951 11713 28963 11747
rect 28905 11707 28963 11713
rect 4617 11679 4675 11685
rect 4617 11676 4629 11679
rect 4172 11648 4629 11676
rect 4172 11620 4200 11648
rect 4617 11645 4629 11648
rect 4663 11645 4675 11679
rect 4617 11639 4675 11645
rect 7653 11679 7711 11685
rect 7653 11645 7665 11679
rect 7699 11676 7711 11679
rect 8849 11679 8907 11685
rect 8849 11676 8861 11679
rect 7699 11648 8861 11676
rect 7699 11645 7711 11648
rect 7653 11639 7711 11645
rect 8849 11645 8861 11648
rect 8895 11676 8907 11679
rect 9674 11676 9680 11688
rect 8895 11648 9680 11676
rect 8895 11645 8907 11648
rect 8849 11639 8907 11645
rect 9674 11636 9680 11648
rect 9732 11676 9738 11688
rect 10870 11676 10876 11688
rect 9732 11648 10876 11676
rect 9732 11636 9738 11648
rect 10870 11636 10876 11648
rect 10928 11636 10934 11688
rect 17034 11636 17040 11688
rect 17092 11676 17098 11688
rect 17313 11679 17371 11685
rect 17313 11676 17325 11679
rect 17092 11648 17325 11676
rect 17092 11636 17098 11648
rect 17313 11645 17325 11648
rect 17359 11645 17371 11679
rect 17313 11639 17371 11645
rect 17494 11636 17500 11688
rect 17552 11636 17558 11688
rect 20254 11636 20260 11688
rect 20312 11676 20318 11688
rect 20622 11676 20628 11688
rect 20312 11648 20628 11676
rect 20312 11636 20318 11648
rect 20622 11636 20628 11648
rect 20680 11676 20686 11688
rect 21177 11679 21235 11685
rect 21177 11676 21189 11679
rect 20680 11648 21189 11676
rect 20680 11636 20686 11648
rect 21177 11645 21189 11648
rect 21223 11645 21235 11679
rect 21177 11639 21235 11645
rect 24854 11636 24860 11688
rect 24912 11636 24918 11688
rect 4154 11568 4160 11620
rect 4212 11568 4218 11620
rect 17512 11608 17540 11636
rect 24762 11608 24768 11620
rect 17512 11580 24768 11608
rect 24762 11568 24768 11580
rect 24820 11568 24826 11620
rect 28644 11608 28672 11707
rect 28920 11676 28948 11707
rect 29546 11704 29552 11756
rect 29604 11704 29610 11756
rect 29638 11676 29644 11688
rect 28920 11648 29644 11676
rect 29638 11636 29644 11648
rect 29696 11676 29702 11688
rect 29840 11685 29868 11784
rect 30650 11772 30656 11784
rect 30708 11812 30714 11824
rect 31202 11812 31208 11824
rect 30708 11784 31208 11812
rect 30708 11772 30714 11784
rect 31202 11772 31208 11784
rect 31260 11772 31266 11824
rect 32122 11772 32128 11824
rect 32180 11812 32186 11824
rect 32180 11784 32628 11812
rect 32180 11772 32186 11784
rect 30552 11747 30610 11753
rect 30552 11713 30564 11747
rect 30598 11744 30610 11747
rect 31846 11744 31852 11756
rect 30598 11716 31852 11744
rect 30598 11713 30610 11716
rect 30552 11707 30610 11713
rect 31846 11704 31852 11716
rect 31904 11704 31910 11756
rect 31938 11704 31944 11756
rect 31996 11744 32002 11756
rect 32493 11747 32551 11753
rect 32493 11744 32505 11747
rect 31996 11716 32505 11744
rect 31996 11704 32002 11716
rect 32493 11713 32505 11716
rect 32539 11713 32551 11747
rect 32600 11744 32628 11784
rect 32766 11772 32772 11824
rect 32824 11812 32830 11824
rect 33137 11815 33195 11821
rect 33137 11812 33149 11815
rect 32824 11784 33149 11812
rect 32824 11772 32830 11784
rect 33137 11781 33149 11784
rect 33183 11781 33195 11815
rect 33353 11815 33411 11821
rect 33353 11812 33365 11815
rect 33137 11775 33195 11781
rect 33244 11784 33365 11812
rect 33244 11744 33272 11784
rect 33353 11781 33365 11784
rect 33399 11812 33411 11815
rect 35618 11812 35624 11824
rect 33399 11784 35624 11812
rect 33399 11781 33411 11784
rect 33353 11775 33411 11781
rect 35618 11772 35624 11784
rect 35676 11772 35682 11824
rect 35710 11772 35716 11824
rect 35768 11812 35774 11824
rect 36449 11815 36507 11821
rect 36449 11812 36461 11815
rect 35768 11784 36461 11812
rect 35768 11772 35774 11784
rect 36449 11781 36461 11784
rect 36495 11812 36507 11815
rect 36495 11784 36952 11812
rect 36495 11781 36507 11784
rect 36449 11775 36507 11781
rect 32600 11716 33272 11744
rect 34232 11747 34290 11753
rect 32493 11707 32551 11713
rect 34232 11713 34244 11747
rect 34278 11744 34290 11747
rect 35250 11744 35256 11756
rect 34278 11716 35256 11744
rect 34278 11713 34290 11716
rect 34232 11707 34290 11713
rect 35250 11704 35256 11716
rect 35308 11704 35314 11756
rect 35802 11704 35808 11756
rect 35860 11704 35866 11756
rect 36078 11704 36084 11756
rect 36136 11744 36142 11756
rect 36630 11744 36636 11756
rect 36136 11716 36636 11744
rect 36136 11704 36142 11716
rect 36630 11704 36636 11716
rect 36688 11704 36694 11756
rect 36924 11744 36952 11784
rect 37734 11772 37740 11824
rect 37792 11772 37798 11824
rect 37946 11815 38004 11821
rect 37946 11781 37958 11815
rect 37992 11812 38004 11815
rect 40862 11812 40868 11824
rect 37992 11784 40868 11812
rect 37992 11781 38004 11784
rect 37946 11775 38004 11781
rect 40862 11772 40868 11784
rect 40920 11772 40926 11824
rect 41782 11772 41788 11824
rect 41840 11812 41846 11824
rect 42242 11812 42248 11824
rect 41840 11784 42248 11812
rect 41840 11772 41846 11784
rect 42242 11772 42248 11784
rect 42300 11812 42306 11824
rect 42794 11812 42800 11824
rect 42300 11784 42800 11812
rect 42300 11772 42306 11784
rect 42794 11772 42800 11784
rect 42852 11772 42858 11824
rect 38378 11744 38384 11756
rect 36924 11716 38384 11744
rect 38378 11704 38384 11716
rect 38436 11704 38442 11756
rect 38838 11704 38844 11756
rect 38896 11704 38902 11756
rect 39025 11747 39083 11753
rect 39025 11713 39037 11747
rect 39071 11744 39083 11747
rect 40773 11747 40831 11753
rect 39071 11716 40264 11744
rect 39071 11713 39083 11716
rect 39025 11707 39083 11713
rect 29733 11679 29791 11685
rect 29733 11676 29745 11679
rect 29696 11648 29745 11676
rect 29696 11636 29702 11648
rect 29733 11645 29745 11648
rect 29779 11645 29791 11679
rect 29733 11639 29791 11645
rect 29825 11679 29883 11685
rect 29825 11645 29837 11679
rect 29871 11645 29883 11679
rect 29825 11639 29883 11645
rect 30282 11636 30288 11688
rect 30340 11636 30346 11688
rect 31754 11636 31760 11688
rect 31812 11676 31818 11688
rect 32309 11679 32367 11685
rect 32309 11676 32321 11679
rect 31812 11648 32321 11676
rect 31812 11636 31818 11648
rect 32309 11645 32321 11648
rect 32355 11645 32367 11679
rect 32309 11639 32367 11645
rect 33502 11636 33508 11688
rect 33560 11676 33566 11688
rect 33686 11676 33692 11688
rect 33560 11648 33692 11676
rect 33560 11636 33566 11648
rect 33686 11636 33692 11648
rect 33744 11676 33750 11688
rect 33965 11679 34023 11685
rect 33965 11676 33977 11679
rect 33744 11648 33977 11676
rect 33744 11636 33750 11648
rect 33965 11645 33977 11648
rect 34011 11645 34023 11679
rect 33965 11639 34023 11645
rect 35345 11611 35403 11617
rect 28644 11580 30328 11608
rect 3237 11543 3295 11549
rect 3237 11509 3249 11543
rect 3283 11540 3295 11543
rect 3970 11540 3976 11552
rect 3283 11512 3976 11540
rect 3283 11509 3295 11512
rect 3237 11503 3295 11509
rect 3970 11500 3976 11512
rect 4028 11500 4034 11552
rect 4062 11500 4068 11552
rect 4120 11540 4126 11552
rect 5626 11540 5632 11552
rect 4120 11512 5632 11540
rect 4120 11500 4126 11512
rect 5626 11500 5632 11512
rect 5684 11500 5690 11552
rect 7009 11543 7067 11549
rect 7009 11509 7021 11543
rect 7055 11540 7067 11543
rect 7190 11540 7196 11552
rect 7055 11512 7196 11540
rect 7055 11509 7067 11512
rect 7009 11503 7067 11509
rect 7190 11500 7196 11512
rect 7248 11500 7254 11552
rect 10137 11543 10195 11549
rect 10137 11509 10149 11543
rect 10183 11540 10195 11543
rect 10226 11540 10232 11552
rect 10183 11512 10232 11540
rect 10183 11509 10195 11512
rect 10137 11503 10195 11509
rect 10226 11500 10232 11512
rect 10284 11500 10290 11552
rect 16850 11500 16856 11552
rect 16908 11500 16914 11552
rect 19061 11543 19119 11549
rect 19061 11509 19073 11543
rect 19107 11540 19119 11543
rect 19702 11540 19708 11552
rect 19107 11512 19708 11540
rect 19107 11509 19119 11512
rect 19061 11503 19119 11509
rect 19702 11500 19708 11512
rect 19760 11500 19766 11552
rect 20990 11500 20996 11552
rect 21048 11500 21054 11552
rect 22373 11543 22431 11549
rect 22373 11509 22385 11543
rect 22419 11540 22431 11543
rect 22646 11540 22652 11552
rect 22419 11512 22652 11540
rect 22419 11509 22431 11512
rect 22373 11503 22431 11509
rect 22646 11500 22652 11512
rect 22704 11500 22710 11552
rect 28629 11543 28687 11549
rect 28629 11509 28641 11543
rect 28675 11540 28687 11543
rect 29638 11540 29644 11552
rect 28675 11512 29644 11540
rect 28675 11509 28687 11512
rect 28629 11503 28687 11509
rect 29638 11500 29644 11512
rect 29696 11500 29702 11552
rect 30300 11540 30328 11580
rect 35345 11577 35357 11611
rect 35391 11608 35403 11611
rect 35820 11608 35848 11704
rect 35986 11636 35992 11688
rect 36044 11676 36050 11688
rect 36817 11679 36875 11685
rect 36817 11676 36829 11679
rect 36044 11648 36829 11676
rect 36044 11636 36050 11648
rect 36817 11645 36829 11648
rect 36863 11645 36875 11679
rect 36817 11639 36875 11645
rect 37461 11679 37519 11685
rect 37461 11645 37473 11679
rect 37507 11645 37519 11679
rect 37461 11639 37519 11645
rect 35391 11580 35848 11608
rect 35391 11577 35403 11580
rect 35345 11571 35403 11577
rect 36538 11568 36544 11620
rect 36596 11608 36602 11620
rect 37476 11608 37504 11639
rect 37550 11636 37556 11688
rect 37608 11676 37614 11688
rect 38102 11676 38108 11688
rect 37608 11648 38108 11676
rect 37608 11636 37614 11648
rect 38102 11636 38108 11648
rect 38160 11636 38166 11688
rect 39206 11636 39212 11688
rect 39264 11636 39270 11688
rect 39301 11679 39359 11685
rect 39301 11645 39313 11679
rect 39347 11645 39359 11679
rect 40236 11676 40264 11716
rect 40773 11713 40785 11747
rect 40819 11744 40831 11747
rect 41506 11744 41512 11756
rect 40819 11716 41512 11744
rect 40819 11713 40831 11716
rect 40773 11707 40831 11713
rect 41506 11704 41512 11716
rect 41564 11704 41570 11756
rect 41598 11704 41604 11756
rect 41656 11704 41662 11756
rect 41877 11747 41935 11753
rect 41877 11713 41889 11747
rect 41923 11744 41935 11747
rect 41966 11744 41972 11756
rect 41923 11716 41972 11744
rect 41923 11713 41935 11716
rect 41877 11707 41935 11713
rect 41966 11704 41972 11716
rect 42024 11704 42030 11756
rect 43162 11676 43168 11688
rect 40236 11648 43168 11676
rect 39301 11639 39359 11645
rect 37642 11608 37648 11620
rect 36596 11580 37648 11608
rect 36596 11568 36602 11580
rect 37642 11568 37648 11580
rect 37700 11608 37706 11620
rect 38286 11608 38292 11620
rect 37700 11580 38292 11608
rect 37700 11568 37706 11580
rect 38286 11568 38292 11580
rect 38344 11568 38350 11620
rect 39316 11608 39344 11639
rect 43162 11636 43168 11648
rect 43220 11636 43226 11688
rect 40034 11608 40040 11620
rect 39316 11580 40040 11608
rect 40034 11568 40040 11580
rect 40092 11608 40098 11620
rect 40865 11611 40923 11617
rect 40865 11608 40877 11611
rect 40092 11580 40877 11608
rect 40092 11568 40098 11580
rect 40865 11577 40877 11580
rect 40911 11577 40923 11611
rect 40865 11571 40923 11577
rect 31665 11543 31723 11549
rect 31665 11540 31677 11543
rect 30300 11512 31677 11540
rect 31665 11509 31677 11512
rect 31711 11540 31723 11543
rect 31754 11540 31760 11552
rect 31711 11512 31760 11540
rect 31711 11509 31723 11512
rect 31665 11503 31723 11509
rect 31754 11500 31760 11512
rect 31812 11540 31818 11552
rect 32766 11540 32772 11552
rect 31812 11512 32772 11540
rect 31812 11500 31818 11512
rect 32766 11500 32772 11512
rect 32824 11500 32830 11552
rect 33318 11500 33324 11552
rect 33376 11500 33382 11552
rect 35894 11500 35900 11552
rect 35952 11500 35958 11552
rect 36722 11500 36728 11552
rect 36780 11500 36786 11552
rect 36909 11543 36967 11549
rect 36909 11509 36921 11543
rect 36955 11540 36967 11543
rect 37550 11540 37556 11552
rect 36955 11512 37556 11540
rect 36955 11509 36967 11512
rect 36909 11503 36967 11509
rect 37550 11500 37556 11512
rect 37608 11500 37614 11552
rect 1104 11450 44896 11472
rect 1104 11398 6423 11450
rect 6475 11398 6487 11450
rect 6539 11398 6551 11450
rect 6603 11398 6615 11450
rect 6667 11398 6679 11450
rect 6731 11398 17370 11450
rect 17422 11398 17434 11450
rect 17486 11398 17498 11450
rect 17550 11398 17562 11450
rect 17614 11398 17626 11450
rect 17678 11398 28317 11450
rect 28369 11398 28381 11450
rect 28433 11398 28445 11450
rect 28497 11398 28509 11450
rect 28561 11398 28573 11450
rect 28625 11398 39264 11450
rect 39316 11398 39328 11450
rect 39380 11398 39392 11450
rect 39444 11398 39456 11450
rect 39508 11398 39520 11450
rect 39572 11398 44896 11450
rect 1104 11376 44896 11398
rect 3418 11296 3424 11348
rect 3476 11296 3482 11348
rect 5534 11296 5540 11348
rect 5592 11296 5598 11348
rect 5994 11296 6000 11348
rect 6052 11296 6058 11348
rect 13648 11308 13860 11336
rect 6733 11271 6791 11277
rect 6733 11237 6745 11271
rect 6779 11237 6791 11271
rect 6733 11231 6791 11237
rect 3970 11160 3976 11212
rect 4028 11200 4034 11212
rect 4028 11172 4292 11200
rect 4028 11160 4034 11172
rect 3142 11092 3148 11144
rect 3200 11092 3206 11144
rect 3234 11092 3240 11144
rect 3292 11092 3298 11144
rect 4154 11092 4160 11144
rect 4212 11092 4218 11144
rect 4264 11132 4292 11172
rect 4413 11135 4471 11141
rect 4413 11132 4425 11135
rect 4264 11104 4425 11132
rect 4413 11101 4425 11104
rect 4459 11101 4471 11135
rect 4413 11095 4471 11101
rect 6181 11135 6239 11141
rect 6181 11101 6193 11135
rect 6227 11132 6239 11135
rect 6748 11132 6776 11231
rect 7190 11160 7196 11212
rect 7248 11160 7254 11212
rect 7377 11203 7435 11209
rect 7377 11169 7389 11203
rect 7423 11200 7435 11203
rect 7558 11200 7564 11212
rect 7423 11172 7564 11200
rect 7423 11169 7435 11172
rect 7377 11163 7435 11169
rect 7558 11160 7564 11172
rect 7616 11160 7622 11212
rect 9858 11160 9864 11212
rect 9916 11200 9922 11212
rect 9953 11203 10011 11209
rect 9953 11200 9965 11203
rect 9916 11172 9965 11200
rect 9916 11160 9922 11172
rect 9953 11169 9965 11172
rect 9999 11169 10011 11203
rect 9953 11163 10011 11169
rect 11422 11160 11428 11212
rect 11480 11200 11486 11212
rect 12345 11203 12403 11209
rect 12345 11200 12357 11203
rect 11480 11172 12357 11200
rect 11480 11160 11486 11172
rect 12345 11169 12357 11172
rect 12391 11169 12403 11203
rect 12345 11163 12403 11169
rect 6227 11104 6776 11132
rect 6227 11101 6239 11104
rect 6181 11095 6239 11101
rect 7926 11092 7932 11144
rect 7984 11092 7990 11144
rect 10226 11141 10232 11144
rect 10220 11132 10232 11141
rect 10187 11104 10232 11132
rect 10220 11095 10232 11104
rect 10226 11092 10232 11095
rect 10284 11092 10290 11144
rect 12612 11135 12670 11141
rect 12612 11101 12624 11135
rect 12658 11132 12670 11135
rect 13648 11132 13676 11308
rect 13725 11271 13783 11277
rect 13725 11237 13737 11271
rect 13771 11237 13783 11271
rect 13832 11268 13860 11308
rect 14642 11296 14648 11348
rect 14700 11296 14706 11348
rect 14752 11308 16712 11336
rect 14752 11268 14780 11308
rect 13832 11240 14780 11268
rect 16684 11268 16712 11308
rect 17126 11296 17132 11348
rect 17184 11296 17190 11348
rect 17862 11296 17868 11348
rect 17920 11336 17926 11348
rect 21177 11339 21235 11345
rect 17920 11308 20760 11336
rect 17920 11296 17926 11308
rect 17880 11268 17908 11296
rect 16684 11240 17908 11268
rect 20732 11268 20760 11308
rect 21177 11305 21189 11339
rect 21223 11336 21235 11339
rect 21450 11336 21456 11348
rect 21223 11308 21456 11336
rect 21223 11305 21235 11308
rect 21177 11299 21235 11305
rect 21450 11296 21456 11308
rect 21508 11296 21514 11348
rect 21818 11296 21824 11348
rect 21876 11336 21882 11348
rect 21876 11308 22876 11336
rect 21876 11296 21882 11308
rect 22848 11280 22876 11308
rect 25498 11296 25504 11348
rect 25556 11296 25562 11348
rect 26142 11296 26148 11348
rect 26200 11296 26206 11348
rect 29638 11296 29644 11348
rect 29696 11336 29702 11348
rect 29696 11308 31754 11336
rect 29696 11296 29702 11308
rect 20732 11240 22094 11268
rect 13725 11231 13783 11237
rect 13740 11200 13768 11231
rect 13740 11172 14504 11200
rect 12658 11104 13676 11132
rect 12658 11101 12670 11104
rect 12612 11095 12670 11101
rect 14366 11092 14372 11144
rect 14424 11092 14430 11144
rect 14476 11141 14504 11172
rect 19702 11160 19708 11212
rect 19760 11160 19766 11212
rect 14461 11135 14519 11141
rect 14461 11101 14473 11135
rect 14507 11101 14519 11135
rect 14461 11095 14519 11101
rect 15749 11135 15807 11141
rect 15749 11101 15761 11135
rect 15795 11132 15807 11135
rect 16758 11132 16764 11144
rect 15795 11104 16764 11132
rect 15795 11101 15807 11104
rect 15749 11095 15807 11101
rect 7101 11067 7159 11073
rect 7101 11033 7113 11067
rect 7147 11064 7159 11067
rect 8294 11064 8300 11076
rect 7147 11036 8300 11064
rect 7147 11033 7159 11036
rect 7101 11027 7159 11033
rect 8294 11024 8300 11036
rect 8352 11024 8358 11076
rect 10870 11024 10876 11076
rect 10928 11064 10934 11076
rect 12342 11064 12348 11076
rect 10928 11036 12348 11064
rect 10928 11024 10934 11036
rect 12342 11024 12348 11036
rect 12400 11024 12406 11076
rect 12894 11024 12900 11076
rect 12952 11064 12958 11076
rect 15764 11064 15792 11095
rect 16758 11092 16764 11104
rect 16816 11132 16822 11144
rect 18506 11132 18512 11144
rect 16816 11104 18512 11132
rect 16816 11092 16822 11104
rect 18506 11092 18512 11104
rect 18564 11132 18570 11144
rect 19429 11135 19487 11141
rect 19429 11132 19441 11135
rect 18564 11104 19441 11132
rect 18564 11092 18570 11104
rect 19429 11101 19441 11104
rect 19475 11101 19487 11135
rect 19429 11095 19487 11101
rect 20806 11092 20812 11144
rect 20864 11092 20870 11144
rect 12952 11036 15792 11064
rect 12952 11024 12958 11036
rect 15838 11024 15844 11076
rect 15896 11064 15902 11076
rect 15994 11067 16052 11073
rect 15994 11064 16006 11067
rect 15896 11036 16006 11064
rect 15896 11024 15902 11036
rect 15994 11033 16006 11036
rect 16040 11033 16052 11067
rect 22066 11064 22094 11240
rect 22830 11228 22836 11280
rect 22888 11268 22894 11280
rect 28902 11268 28908 11280
rect 22888 11240 28908 11268
rect 22888 11228 22894 11240
rect 22646 11092 22652 11144
rect 22704 11092 22710 11144
rect 24596 11141 24624 11240
rect 28902 11228 28908 11240
rect 28960 11228 28966 11280
rect 31726 11268 31754 11308
rect 31846 11296 31852 11348
rect 31904 11336 31910 11348
rect 32585 11339 32643 11345
rect 32585 11336 32597 11339
rect 31904 11308 32597 11336
rect 31904 11296 31910 11308
rect 32585 11305 32597 11308
rect 32631 11305 32643 11339
rect 32585 11299 32643 11305
rect 33226 11296 33232 11348
rect 33284 11336 33290 11348
rect 35161 11339 35219 11345
rect 35161 11336 35173 11339
rect 33284 11308 35173 11336
rect 33284 11296 33290 11308
rect 35161 11305 35173 11308
rect 35207 11305 35219 11339
rect 35161 11299 35219 11305
rect 35250 11296 35256 11348
rect 35308 11296 35314 11348
rect 36722 11296 36728 11348
rect 36780 11336 36786 11348
rect 39209 11339 39267 11345
rect 39209 11336 39221 11339
rect 36780 11308 39221 11336
rect 36780 11296 36786 11308
rect 39209 11305 39221 11308
rect 39255 11305 39267 11339
rect 39209 11299 39267 11305
rect 32677 11271 32735 11277
rect 32677 11268 32689 11271
rect 31726 11240 32689 11268
rect 32677 11237 32689 11240
rect 32723 11237 32735 11271
rect 32677 11231 32735 11237
rect 36446 11228 36452 11280
rect 36504 11268 36510 11280
rect 37369 11271 37427 11277
rect 37369 11268 37381 11271
rect 36504 11240 37381 11268
rect 36504 11228 36510 11240
rect 37369 11237 37381 11240
rect 37415 11237 37427 11271
rect 38378 11268 38384 11280
rect 37369 11231 37427 11237
rect 37568 11240 38384 11268
rect 24762 11160 24768 11212
rect 24820 11160 24826 11212
rect 25038 11160 25044 11212
rect 25096 11200 25102 11212
rect 33134 11200 33140 11212
rect 25096 11172 33140 11200
rect 25096 11160 25102 11172
rect 33134 11160 33140 11172
rect 33192 11160 33198 11212
rect 35894 11200 35900 11212
rect 35084 11172 35900 11200
rect 24581 11135 24639 11141
rect 24581 11101 24593 11135
rect 24627 11101 24639 11135
rect 24581 11095 24639 11101
rect 24670 11092 24676 11144
rect 24728 11092 24734 11144
rect 24949 11135 25007 11141
rect 24949 11101 24961 11135
rect 24995 11132 25007 11135
rect 25314 11132 25320 11144
rect 24995 11104 25320 11132
rect 24995 11101 25007 11104
rect 24949 11095 25007 11101
rect 25314 11092 25320 11104
rect 25372 11092 25378 11144
rect 25406 11092 25412 11144
rect 25464 11092 25470 11144
rect 25498 11092 25504 11144
rect 25556 11132 25562 11144
rect 26050 11132 26056 11144
rect 25556 11104 26056 11132
rect 25556 11092 25562 11104
rect 26050 11092 26056 11104
rect 26108 11092 26114 11144
rect 29178 11092 29184 11144
rect 29236 11132 29242 11144
rect 29730 11132 29736 11144
rect 29236 11104 29736 11132
rect 29236 11092 29242 11104
rect 29730 11092 29736 11104
rect 29788 11132 29794 11144
rect 30282 11132 30288 11144
rect 29788 11104 30288 11132
rect 29788 11092 29794 11104
rect 30282 11092 30288 11104
rect 30340 11092 30346 11144
rect 30650 11092 30656 11144
rect 30708 11092 30714 11144
rect 32079 11135 32137 11141
rect 32079 11101 32091 11135
rect 32125 11132 32137 11135
rect 32490 11132 32496 11144
rect 32125 11104 32496 11132
rect 32125 11101 32137 11104
rect 32079 11095 32137 11101
rect 32490 11092 32496 11104
rect 32548 11092 32554 11144
rect 32582 11092 32588 11144
rect 32640 11092 32646 11144
rect 32674 11092 32680 11144
rect 32732 11132 32738 11144
rect 32861 11135 32919 11141
rect 32861 11132 32873 11135
rect 32732 11104 32873 11132
rect 32732 11092 32738 11104
rect 32861 11101 32873 11104
rect 32907 11132 32919 11135
rect 34974 11132 34980 11144
rect 32907 11104 34980 11132
rect 32907 11101 32919 11104
rect 32861 11095 32919 11101
rect 34974 11092 34980 11104
rect 35032 11092 35038 11144
rect 35084 11141 35112 11172
rect 35894 11160 35900 11172
rect 35952 11160 35958 11212
rect 37568 11200 37596 11240
rect 38378 11228 38384 11240
rect 38436 11228 38442 11280
rect 38470 11228 38476 11280
rect 38528 11268 38534 11280
rect 39114 11268 39120 11280
rect 38528 11240 39120 11268
rect 38528 11228 38534 11240
rect 39114 11228 39120 11240
rect 39172 11268 39178 11280
rect 39172 11240 39896 11268
rect 39172 11228 39178 11240
rect 38746 11200 38752 11212
rect 37476 11172 37596 11200
rect 38212 11172 38752 11200
rect 35069 11135 35127 11141
rect 35069 11101 35081 11135
rect 35115 11101 35127 11135
rect 35069 11095 35127 11101
rect 35158 11092 35164 11144
rect 35216 11132 35222 11144
rect 35253 11135 35311 11141
rect 35253 11132 35265 11135
rect 35216 11104 35265 11132
rect 35216 11092 35222 11104
rect 35253 11101 35265 11104
rect 35299 11132 35311 11135
rect 35986 11132 35992 11144
rect 35299 11104 35992 11132
rect 35299 11101 35311 11104
rect 35253 11095 35311 11101
rect 35986 11092 35992 11104
rect 36044 11092 36050 11144
rect 36538 11092 36544 11144
rect 36596 11092 36602 11144
rect 36817 11135 36875 11141
rect 36817 11101 36829 11135
rect 36863 11132 36875 11135
rect 37277 11135 37335 11141
rect 37277 11132 37289 11135
rect 36863 11104 37289 11132
rect 36863 11101 36875 11104
rect 36817 11095 36875 11101
rect 37277 11101 37289 11104
rect 37323 11132 37335 11135
rect 37476 11132 37504 11172
rect 37323 11104 37504 11132
rect 37553 11135 37611 11141
rect 37323 11101 37335 11104
rect 37277 11095 37335 11101
rect 37553 11101 37565 11135
rect 37599 11132 37611 11135
rect 37642 11132 37648 11144
rect 37599 11104 37648 11132
rect 37599 11101 37611 11104
rect 37553 11095 37611 11101
rect 37642 11092 37648 11104
rect 37700 11092 37706 11144
rect 38010 11092 38016 11144
rect 38068 11092 38074 11144
rect 38212 11141 38240 11172
rect 38746 11160 38752 11172
rect 38804 11160 38810 11212
rect 38930 11160 38936 11212
rect 38988 11200 38994 11212
rect 38988 11172 39436 11200
rect 38988 11160 38994 11172
rect 38197 11135 38255 11141
rect 38197 11101 38209 11135
rect 38243 11101 38255 11135
rect 38197 11095 38255 11101
rect 38286 11092 38292 11144
rect 38344 11092 38350 11144
rect 38381 11135 38439 11141
rect 38381 11101 38393 11135
rect 38427 11132 38439 11135
rect 38470 11132 38476 11144
rect 38427 11104 38476 11132
rect 38427 11101 38439 11104
rect 38381 11095 38439 11101
rect 38470 11092 38476 11104
rect 38528 11092 38534 11144
rect 38565 11135 38623 11141
rect 38565 11101 38577 11135
rect 38611 11132 38623 11135
rect 38654 11132 38660 11144
rect 38611 11104 38660 11132
rect 38611 11101 38623 11104
rect 38565 11095 38623 11101
rect 38654 11092 38660 11104
rect 38712 11132 38718 11144
rect 38838 11132 38844 11144
rect 38712 11104 38844 11132
rect 38712 11092 38718 11104
rect 38838 11092 38844 11104
rect 38896 11132 38902 11144
rect 39408 11141 39436 11172
rect 39209 11135 39267 11141
rect 39209 11132 39221 11135
rect 38896 11104 39221 11132
rect 38896 11092 38902 11104
rect 39209 11101 39221 11104
rect 39255 11101 39267 11135
rect 39209 11095 39267 11101
rect 39393 11135 39451 11141
rect 39393 11101 39405 11135
rect 39439 11101 39451 11135
rect 39393 11095 39451 11101
rect 39485 11135 39543 11141
rect 39485 11101 39497 11135
rect 39531 11132 39543 11135
rect 39758 11132 39764 11144
rect 39531 11104 39764 11132
rect 39531 11101 39543 11104
rect 39485 11095 39543 11101
rect 26234 11064 26240 11076
rect 22066 11036 26240 11064
rect 15994 11027 16052 11033
rect 26234 11024 26240 11036
rect 26292 11024 26298 11076
rect 32398 11064 32404 11076
rect 31694 11036 32404 11064
rect 32398 11024 32404 11036
rect 32456 11024 32462 11076
rect 34885 11067 34943 11073
rect 34885 11033 34897 11067
rect 34931 11064 34943 11067
rect 36446 11064 36452 11076
rect 34931 11036 36452 11064
rect 34931 11033 34943 11036
rect 34885 11027 34943 11033
rect 36446 11024 36452 11036
rect 36504 11024 36510 11076
rect 36630 11024 36636 11076
rect 36688 11064 36694 11076
rect 36725 11067 36783 11073
rect 36725 11064 36737 11067
rect 36688 11036 36737 11064
rect 36688 11024 36694 11036
rect 36725 11033 36737 11036
rect 36771 11064 36783 11067
rect 37461 11067 37519 11073
rect 37461 11064 37473 11067
rect 36771 11036 37473 11064
rect 36771 11033 36783 11036
rect 36725 11027 36783 11033
rect 37461 11033 37473 11036
rect 37507 11064 37519 11067
rect 37507 11036 37872 11064
rect 37507 11033 37519 11036
rect 37461 11027 37519 11033
rect 8573 10999 8631 11005
rect 8573 10965 8585 10999
rect 8619 10996 8631 10999
rect 9582 10996 9588 11008
rect 8619 10968 9588 10996
rect 8619 10965 8631 10968
rect 8573 10959 8631 10965
rect 9582 10956 9588 10968
rect 9640 10956 9646 11008
rect 11330 10956 11336 11008
rect 11388 10956 11394 11008
rect 17218 10956 17224 11008
rect 17276 10996 17282 11008
rect 21082 10996 21088 11008
rect 17276 10968 21088 10996
rect 17276 10956 17282 10968
rect 21082 10956 21088 10968
rect 21140 10956 21146 11008
rect 22465 10999 22523 11005
rect 22465 10965 22477 10999
rect 22511 10996 22523 10999
rect 23198 10996 23204 11008
rect 22511 10968 23204 10996
rect 22511 10965 22523 10968
rect 22465 10959 22523 10965
rect 23198 10956 23204 10968
rect 23256 10956 23262 11008
rect 24857 10999 24915 11005
rect 24857 10965 24869 10999
rect 24903 10996 24915 10999
rect 24946 10996 24952 11008
rect 24903 10968 24952 10996
rect 24903 10965 24915 10968
rect 24857 10959 24915 10965
rect 24946 10956 24952 10968
rect 25004 10956 25010 11008
rect 25222 10956 25228 11008
rect 25280 10996 25286 11008
rect 26050 10996 26056 11008
rect 25280 10968 26056 10996
rect 25280 10956 25286 10968
rect 26050 10956 26056 10968
rect 26108 10956 26114 11008
rect 30926 10956 30932 11008
rect 30984 10996 30990 11008
rect 32674 10996 32680 11008
rect 30984 10968 32680 10996
rect 30984 10956 30990 10968
rect 32674 10956 32680 10968
rect 32732 10956 32738 11008
rect 36354 10956 36360 11008
rect 36412 10956 36418 11008
rect 37844 10996 37872 11036
rect 37918 11024 37924 11076
rect 37976 11064 37982 11076
rect 38749 11067 38807 11073
rect 38749 11064 38761 11067
rect 37976 11036 38761 11064
rect 37976 11024 37982 11036
rect 38749 11033 38761 11036
rect 38795 11033 38807 11067
rect 39500 11064 39528 11095
rect 39758 11092 39764 11104
rect 39816 11092 39822 11144
rect 38749 11027 38807 11033
rect 38856 11036 39528 11064
rect 39868 11064 39896 11240
rect 40586 11160 40592 11212
rect 40644 11200 40650 11212
rect 41417 11203 41475 11209
rect 41417 11200 41429 11203
rect 40644 11172 41429 11200
rect 40644 11160 40650 11172
rect 41417 11169 41429 11172
rect 41463 11169 41475 11203
rect 41417 11163 41475 11169
rect 41690 11141 41696 11144
rect 41684 11132 41696 11141
rect 41651 11104 41696 11132
rect 41684 11095 41696 11104
rect 41690 11092 41696 11095
rect 41748 11092 41754 11144
rect 44361 11135 44419 11141
rect 44361 11101 44373 11135
rect 44407 11132 44419 11135
rect 45002 11132 45008 11144
rect 44407 11104 45008 11132
rect 44407 11101 44419 11104
rect 44361 11095 44419 11101
rect 45002 11092 45008 11104
rect 45060 11092 45066 11144
rect 42886 11064 42892 11076
rect 39868 11036 42892 11064
rect 38856 10996 38884 11036
rect 42886 11024 42892 11036
rect 42944 11024 42950 11076
rect 37844 10968 38884 10996
rect 42794 10956 42800 11008
rect 42852 10956 42858 11008
rect 1104 10906 45051 10928
rect 1104 10854 11896 10906
rect 11948 10854 11960 10906
rect 12012 10854 12024 10906
rect 12076 10854 12088 10906
rect 12140 10854 12152 10906
rect 12204 10854 22843 10906
rect 22895 10854 22907 10906
rect 22959 10854 22971 10906
rect 23023 10854 23035 10906
rect 23087 10854 23099 10906
rect 23151 10854 33790 10906
rect 33842 10854 33854 10906
rect 33906 10854 33918 10906
rect 33970 10854 33982 10906
rect 34034 10854 34046 10906
rect 34098 10854 44737 10906
rect 44789 10854 44801 10906
rect 44853 10854 44865 10906
rect 44917 10854 44929 10906
rect 44981 10854 44993 10906
rect 45045 10854 45051 10906
rect 1104 10832 45051 10854
rect 2317 10795 2375 10801
rect 2317 10761 2329 10795
rect 2363 10792 2375 10795
rect 2363 10764 2774 10792
rect 2363 10761 2375 10764
rect 2317 10755 2375 10761
rect 2746 10724 2774 10764
rect 4614 10752 4620 10804
rect 4672 10792 4678 10804
rect 5353 10795 5411 10801
rect 5353 10792 5365 10795
rect 4672 10764 5365 10792
rect 4672 10752 4678 10764
rect 5353 10761 5365 10764
rect 5399 10761 5411 10795
rect 5353 10755 5411 10761
rect 8294 10752 8300 10804
rect 8352 10752 8358 10804
rect 9585 10795 9643 10801
rect 9585 10761 9597 10795
rect 9631 10792 9643 10795
rect 10321 10795 10379 10801
rect 10321 10792 10333 10795
rect 9631 10764 10333 10792
rect 9631 10761 9643 10764
rect 9585 10755 9643 10761
rect 10321 10761 10333 10764
rect 10367 10761 10379 10795
rect 10321 10755 10379 10761
rect 10778 10752 10784 10804
rect 10836 10752 10842 10804
rect 13081 10795 13139 10801
rect 13081 10761 13093 10795
rect 13127 10792 13139 10795
rect 14001 10795 14059 10801
rect 14001 10792 14013 10795
rect 13127 10764 14013 10792
rect 13127 10761 13139 10764
rect 13081 10755 13139 10761
rect 14001 10761 14013 10764
rect 14047 10761 14059 10795
rect 14001 10755 14059 10761
rect 15473 10795 15531 10801
rect 15473 10761 15485 10795
rect 15519 10792 15531 10795
rect 15838 10792 15844 10804
rect 15519 10764 15844 10792
rect 15519 10761 15531 10764
rect 15473 10755 15531 10761
rect 15838 10752 15844 10764
rect 15896 10752 15902 10804
rect 16117 10795 16175 10801
rect 16117 10761 16129 10795
rect 16163 10792 16175 10795
rect 16574 10792 16580 10804
rect 16163 10764 16580 10792
rect 16163 10761 16175 10764
rect 16117 10755 16175 10761
rect 16574 10752 16580 10764
rect 16632 10752 16638 10804
rect 16945 10795 17003 10801
rect 16945 10761 16957 10795
rect 16991 10792 17003 10795
rect 17034 10792 17040 10804
rect 16991 10764 17040 10792
rect 16991 10761 17003 10764
rect 16945 10755 17003 10761
rect 17034 10752 17040 10764
rect 17092 10752 17098 10804
rect 17126 10752 17132 10804
rect 17184 10792 17190 10804
rect 17313 10795 17371 10801
rect 17313 10792 17325 10795
rect 17184 10764 17325 10792
rect 17184 10752 17190 10764
rect 17313 10761 17325 10764
rect 17359 10761 17371 10795
rect 17313 10755 17371 10761
rect 18690 10752 18696 10804
rect 18748 10792 18754 10804
rect 18748 10764 20760 10792
rect 18748 10752 18754 10764
rect 3142 10724 3148 10736
rect 2746 10696 3148 10724
rect 3142 10684 3148 10696
rect 3200 10724 3206 10736
rect 6086 10724 6092 10736
rect 3200 10696 6092 10724
rect 3200 10684 3206 10696
rect 6086 10684 6092 10696
rect 6144 10684 6150 10736
rect 9858 10724 9864 10736
rect 6932 10696 9864 10724
rect 1946 10616 1952 10668
rect 2004 10656 2010 10668
rect 2133 10659 2191 10665
rect 2133 10656 2145 10659
rect 2004 10628 2145 10656
rect 2004 10616 2010 10628
rect 2133 10625 2145 10628
rect 2179 10625 2191 10659
rect 2133 10619 2191 10625
rect 3973 10659 4031 10665
rect 3973 10625 3985 10659
rect 4019 10656 4031 10659
rect 4062 10656 4068 10668
rect 4019 10628 4068 10656
rect 4019 10625 4031 10628
rect 3973 10619 4031 10625
rect 4062 10616 4068 10628
rect 4120 10616 4126 10668
rect 4246 10665 4252 10668
rect 4240 10619 4252 10665
rect 4246 10616 4252 10619
rect 4304 10616 4310 10668
rect 6932 10665 6960 10696
rect 9858 10684 9864 10696
rect 9916 10684 9922 10736
rect 10689 10727 10747 10733
rect 10689 10693 10701 10727
rect 10735 10724 10747 10727
rect 11330 10724 11336 10736
rect 10735 10696 11336 10724
rect 10735 10693 10747 10696
rect 10689 10687 10747 10693
rect 11330 10684 11336 10696
rect 11388 10724 11394 10736
rect 11946 10727 12004 10733
rect 11946 10724 11958 10727
rect 11388 10696 11958 10724
rect 11388 10684 11394 10696
rect 11946 10693 11958 10696
rect 11992 10693 12004 10727
rect 16850 10724 16856 10736
rect 11946 10687 12004 10693
rect 15672 10696 16856 10724
rect 6917 10659 6975 10665
rect 6917 10625 6929 10659
rect 6963 10625 6975 10659
rect 6917 10619 6975 10625
rect 7184 10659 7242 10665
rect 7184 10625 7196 10659
rect 7230 10656 7242 10659
rect 8386 10656 8392 10668
rect 7230 10628 8392 10656
rect 7230 10625 7242 10628
rect 7184 10619 7242 10625
rect 8386 10616 8392 10628
rect 8444 10616 8450 10668
rect 9493 10659 9551 10665
rect 9493 10625 9505 10659
rect 9539 10656 9551 10659
rect 10962 10656 10968 10668
rect 9539 10628 10968 10656
rect 9539 10625 9551 10628
rect 9493 10619 9551 10625
rect 10962 10616 10968 10628
rect 11020 10616 11026 10668
rect 11422 10616 11428 10668
rect 11480 10656 11486 10668
rect 11701 10659 11759 10665
rect 11701 10656 11713 10659
rect 11480 10628 11713 10656
rect 11480 10616 11486 10628
rect 11701 10625 11713 10628
rect 11747 10625 11759 10659
rect 11701 10619 11759 10625
rect 13906 10616 13912 10668
rect 13964 10616 13970 10668
rect 13998 10616 14004 10668
rect 14056 10656 14062 10668
rect 15672 10665 15700 10696
rect 16850 10684 16856 10696
rect 16908 10684 16914 10736
rect 20254 10684 20260 10736
rect 20312 10684 20318 10736
rect 15013 10659 15071 10665
rect 15013 10656 15025 10659
rect 14056 10628 15025 10656
rect 14056 10616 14062 10628
rect 15013 10625 15025 10628
rect 15059 10625 15071 10659
rect 15013 10619 15071 10625
rect 15657 10659 15715 10665
rect 15657 10625 15669 10659
rect 15703 10625 15715 10659
rect 15657 10619 15715 10625
rect 16298 10616 16304 10668
rect 16356 10616 16362 10668
rect 17218 10616 17224 10668
rect 17276 10656 17282 10668
rect 18877 10659 18935 10665
rect 17276 10628 17540 10656
rect 17276 10616 17282 10628
rect 2961 10591 3019 10597
rect 2961 10557 2973 10591
rect 3007 10557 3019 10591
rect 2961 10551 3019 10557
rect 9769 10591 9827 10597
rect 9769 10557 9781 10591
rect 9815 10588 9827 10591
rect 9815 10560 10824 10588
rect 9815 10557 9827 10560
rect 9769 10551 9827 10557
rect 2976 10520 3004 10551
rect 9125 10523 9183 10529
rect 2976 10492 4016 10520
rect 3142 10412 3148 10464
rect 3200 10452 3206 10464
rect 3513 10455 3571 10461
rect 3513 10452 3525 10455
rect 3200 10424 3525 10452
rect 3200 10412 3206 10424
rect 3513 10421 3525 10424
rect 3559 10421 3571 10455
rect 3988 10452 4016 10492
rect 9125 10489 9137 10523
rect 9171 10520 9183 10523
rect 10318 10520 10324 10532
rect 9171 10492 10324 10520
rect 9171 10489 9183 10492
rect 9125 10483 9183 10489
rect 10318 10480 10324 10492
rect 10376 10480 10382 10532
rect 10796 10520 10824 10560
rect 10870 10548 10876 10600
rect 10928 10548 10934 10600
rect 14090 10548 14096 10600
rect 14148 10548 14154 10600
rect 17512 10597 17540 10628
rect 18877 10625 18889 10659
rect 18923 10656 18935 10659
rect 19426 10656 19432 10668
rect 18923 10628 19432 10656
rect 18923 10625 18935 10628
rect 18877 10619 18935 10625
rect 19426 10616 19432 10628
rect 19484 10616 19490 10668
rect 20073 10659 20131 10665
rect 20073 10625 20085 10659
rect 20119 10656 20131 10659
rect 20162 10656 20168 10668
rect 20119 10628 20168 10656
rect 20119 10625 20131 10628
rect 20073 10619 20131 10625
rect 20162 10616 20168 10628
rect 20220 10616 20226 10668
rect 20732 10665 20760 10764
rect 20806 10752 20812 10804
rect 20864 10752 20870 10804
rect 21082 10752 21088 10804
rect 21140 10792 21146 10804
rect 22646 10792 22652 10804
rect 21140 10764 22652 10792
rect 21140 10752 21146 10764
rect 22646 10752 22652 10764
rect 22704 10752 22710 10804
rect 25222 10792 25228 10804
rect 22756 10764 25228 10792
rect 22756 10724 22784 10764
rect 25222 10752 25228 10764
rect 25280 10752 25286 10804
rect 25314 10752 25320 10804
rect 25372 10792 25378 10804
rect 26142 10792 26148 10804
rect 25372 10764 26148 10792
rect 25372 10752 25378 10764
rect 26142 10752 26148 10764
rect 26200 10752 26206 10804
rect 27341 10795 27399 10801
rect 27341 10761 27353 10795
rect 27387 10792 27399 10795
rect 27430 10792 27436 10804
rect 27387 10764 27436 10792
rect 27387 10761 27399 10764
rect 27341 10755 27399 10761
rect 27430 10752 27436 10764
rect 27488 10752 27494 10804
rect 30650 10752 30656 10804
rect 30708 10792 30714 10804
rect 30837 10795 30895 10801
rect 30837 10792 30849 10795
rect 30708 10764 30849 10792
rect 30708 10752 30714 10764
rect 30837 10761 30849 10764
rect 30883 10761 30895 10795
rect 30837 10755 30895 10761
rect 30926 10752 30932 10804
rect 30984 10792 30990 10804
rect 31205 10795 31263 10801
rect 31205 10792 31217 10795
rect 30984 10764 31217 10792
rect 30984 10752 30990 10764
rect 31205 10761 31217 10764
rect 31251 10761 31263 10795
rect 31205 10755 31263 10761
rect 32398 10752 32404 10804
rect 32456 10752 32462 10804
rect 36357 10795 36415 10801
rect 36357 10761 36369 10795
rect 36403 10792 36415 10795
rect 36446 10792 36452 10804
rect 36403 10764 36452 10792
rect 36403 10761 36415 10764
rect 36357 10755 36415 10761
rect 36446 10752 36452 10764
rect 36504 10752 36510 10804
rect 38838 10752 38844 10804
rect 38896 10752 38902 10804
rect 39022 10752 39028 10804
rect 39080 10792 39086 10804
rect 39761 10795 39819 10801
rect 39761 10792 39773 10795
rect 39080 10764 39773 10792
rect 39080 10752 39086 10764
rect 39761 10761 39773 10764
rect 39807 10761 39819 10795
rect 39761 10755 39819 10761
rect 43162 10752 43168 10804
rect 43220 10752 43226 10804
rect 22664 10696 22784 10724
rect 23109 10727 23167 10733
rect 20717 10659 20775 10665
rect 20717 10625 20729 10659
rect 20763 10656 20775 10659
rect 22097 10659 22155 10665
rect 22097 10656 22109 10659
rect 20763 10628 22109 10656
rect 20763 10625 20775 10628
rect 20717 10619 20775 10625
rect 22097 10625 22109 10628
rect 22143 10656 22155 10659
rect 22664 10656 22692 10696
rect 23109 10693 23121 10727
rect 23155 10724 23167 10727
rect 23198 10724 23204 10736
rect 23155 10696 23204 10724
rect 23155 10693 23167 10696
rect 23109 10687 23167 10693
rect 23198 10684 23204 10696
rect 23256 10684 23262 10736
rect 24670 10724 24676 10736
rect 24334 10696 24676 10724
rect 24670 10684 24676 10696
rect 24728 10684 24734 10736
rect 24762 10684 24768 10736
rect 24820 10724 24826 10736
rect 25501 10727 25559 10733
rect 25501 10724 25513 10727
rect 24820 10696 25513 10724
rect 24820 10684 24826 10696
rect 25501 10693 25513 10696
rect 25547 10693 25559 10727
rect 25501 10687 25559 10693
rect 25774 10684 25780 10736
rect 25832 10724 25838 10736
rect 33781 10727 33839 10733
rect 33781 10724 33793 10727
rect 25832 10696 26280 10724
rect 25832 10684 25838 10696
rect 22143 10628 22692 10656
rect 25409 10659 25467 10665
rect 22143 10625 22155 10628
rect 22097 10619 22155 10625
rect 25409 10625 25421 10659
rect 25455 10656 25467 10659
rect 25792 10656 25820 10684
rect 25455 10628 25820 10656
rect 25455 10625 25467 10628
rect 25409 10619 25467 10625
rect 26050 10616 26056 10668
rect 26108 10616 26114 10668
rect 26252 10665 26280 10696
rect 28736 10696 33793 10724
rect 28736 10668 28764 10696
rect 33781 10693 33793 10696
rect 33827 10693 33839 10727
rect 33781 10687 33839 10693
rect 38654 10684 38660 10736
rect 38712 10724 38718 10736
rect 39301 10727 39359 10733
rect 39301 10724 39313 10727
rect 38712 10696 39313 10724
rect 38712 10684 38718 10696
rect 39301 10693 39313 10696
rect 39347 10724 39359 10727
rect 44450 10724 44456 10736
rect 39347 10696 44456 10724
rect 39347 10693 39359 10696
rect 39301 10687 39359 10693
rect 44450 10684 44456 10696
rect 44508 10684 44514 10736
rect 26237 10659 26295 10665
rect 26237 10625 26249 10659
rect 26283 10625 26295 10659
rect 26237 10619 26295 10625
rect 27246 10616 27252 10668
rect 27304 10656 27310 10668
rect 27614 10656 27620 10668
rect 27304 10628 27620 10656
rect 27304 10616 27310 10628
rect 27614 10616 27620 10628
rect 27672 10616 27678 10668
rect 28629 10659 28687 10665
rect 28629 10625 28641 10659
rect 28675 10656 28687 10659
rect 28718 10656 28724 10668
rect 28675 10628 28724 10656
rect 28675 10625 28687 10628
rect 28629 10619 28687 10625
rect 28718 10616 28724 10628
rect 28776 10616 28782 10668
rect 31021 10659 31079 10665
rect 31021 10625 31033 10659
rect 31067 10625 31079 10659
rect 31021 10619 31079 10625
rect 17405 10591 17463 10597
rect 17405 10557 17417 10591
rect 17451 10557 17463 10591
rect 17405 10551 17463 10557
rect 17497 10591 17555 10597
rect 17497 10557 17509 10591
rect 17543 10557 17555 10591
rect 17497 10551 17555 10557
rect 11054 10520 11060 10532
rect 10796 10492 11060 10520
rect 11054 10480 11060 10492
rect 11112 10480 11118 10532
rect 13541 10523 13599 10529
rect 13541 10489 13553 10523
rect 13587 10520 13599 10523
rect 14182 10520 14188 10532
rect 13587 10492 14188 10520
rect 13587 10489 13599 10492
rect 13541 10483 13599 10489
rect 14182 10480 14188 10492
rect 14240 10480 14246 10532
rect 17420 10520 17448 10551
rect 21174 10548 21180 10600
rect 21232 10588 21238 10600
rect 22554 10588 22560 10600
rect 21232 10560 22560 10588
rect 21232 10548 21238 10560
rect 22554 10548 22560 10560
rect 22612 10588 22618 10600
rect 22833 10591 22891 10597
rect 22833 10588 22845 10591
rect 22612 10560 22845 10588
rect 22612 10548 22618 10560
rect 22833 10557 22845 10560
rect 22879 10557 22891 10591
rect 22833 10551 22891 10557
rect 24578 10548 24584 10600
rect 24636 10588 24642 10600
rect 24857 10591 24915 10597
rect 24857 10588 24869 10591
rect 24636 10560 24869 10588
rect 24636 10548 24642 10560
rect 24857 10557 24869 10560
rect 24903 10588 24915 10591
rect 31036 10588 31064 10619
rect 31294 10616 31300 10668
rect 31352 10616 31358 10668
rect 32309 10659 32367 10665
rect 32309 10625 32321 10659
rect 32355 10625 32367 10659
rect 32309 10619 32367 10625
rect 24903 10560 31064 10588
rect 24903 10557 24915 10560
rect 24857 10551 24915 10557
rect 17420 10492 22968 10520
rect 4614 10452 4620 10464
rect 3988 10424 4620 10452
rect 3513 10415 3571 10421
rect 4614 10412 4620 10424
rect 4672 10412 4678 10464
rect 14829 10455 14887 10461
rect 14829 10421 14841 10455
rect 14875 10452 14887 10455
rect 15194 10452 15200 10464
rect 14875 10424 15200 10452
rect 14875 10421 14887 10424
rect 14829 10415 14887 10421
rect 15194 10412 15200 10424
rect 15252 10412 15258 10464
rect 18690 10412 18696 10464
rect 18748 10412 18754 10464
rect 22186 10412 22192 10464
rect 22244 10412 22250 10464
rect 22940 10452 22968 10492
rect 25406 10480 25412 10532
rect 25464 10520 25470 10532
rect 32324 10520 32352 10619
rect 35986 10616 35992 10668
rect 36044 10616 36050 10668
rect 36814 10616 36820 10668
rect 36872 10656 36878 10668
rect 37461 10659 37519 10665
rect 37461 10656 37473 10659
rect 36872 10628 37473 10656
rect 36872 10616 36878 10628
rect 37461 10625 37473 10628
rect 37507 10625 37519 10659
rect 37461 10619 37519 10625
rect 37550 10616 37556 10668
rect 37608 10656 37614 10668
rect 37717 10659 37775 10665
rect 37717 10656 37729 10659
rect 37608 10628 37729 10656
rect 37608 10616 37614 10628
rect 37717 10625 37729 10628
rect 37763 10625 37775 10659
rect 37717 10619 37775 10625
rect 42794 10616 42800 10668
rect 42852 10616 42858 10668
rect 42889 10591 42947 10597
rect 42889 10557 42901 10591
rect 42935 10588 42947 10591
rect 44266 10588 44272 10600
rect 42935 10560 44272 10588
rect 42935 10557 42947 10560
rect 42889 10551 42947 10557
rect 44266 10548 44272 10560
rect 44324 10548 44330 10600
rect 32858 10520 32864 10532
rect 25464 10492 32864 10520
rect 25464 10480 25470 10492
rect 32858 10480 32864 10492
rect 32916 10480 32922 10532
rect 38470 10480 38476 10532
rect 38528 10520 38534 10532
rect 39577 10523 39635 10529
rect 39577 10520 39589 10523
rect 38528 10492 39589 10520
rect 38528 10480 38534 10492
rect 39577 10489 39589 10492
rect 39623 10489 39635 10523
rect 39577 10483 39635 10489
rect 25314 10452 25320 10464
rect 22940 10424 25320 10452
rect 25314 10412 25320 10424
rect 25372 10412 25378 10464
rect 29730 10412 29736 10464
rect 29788 10452 29794 10464
rect 29917 10455 29975 10461
rect 29917 10452 29929 10455
rect 29788 10424 29929 10452
rect 29788 10412 29794 10424
rect 29917 10421 29929 10424
rect 29963 10421 29975 10455
rect 29917 10415 29975 10421
rect 33502 10412 33508 10464
rect 33560 10452 33566 10464
rect 35069 10455 35127 10461
rect 35069 10452 35081 10455
rect 33560 10424 35081 10452
rect 33560 10412 33566 10424
rect 35069 10421 35081 10424
rect 35115 10452 35127 10455
rect 36262 10452 36268 10464
rect 35115 10424 36268 10452
rect 35115 10421 35127 10424
rect 35069 10415 35127 10421
rect 36262 10412 36268 10424
rect 36320 10412 36326 10464
rect 36354 10412 36360 10464
rect 36412 10412 36418 10464
rect 36541 10455 36599 10461
rect 36541 10421 36553 10455
rect 36587 10452 36599 10455
rect 36906 10452 36912 10464
rect 36587 10424 36912 10452
rect 36587 10421 36599 10424
rect 36541 10415 36599 10421
rect 36906 10412 36912 10424
rect 36964 10412 36970 10464
rect 1104 10362 44896 10384
rect 1104 10310 6423 10362
rect 6475 10310 6487 10362
rect 6539 10310 6551 10362
rect 6603 10310 6615 10362
rect 6667 10310 6679 10362
rect 6731 10310 17370 10362
rect 17422 10310 17434 10362
rect 17486 10310 17498 10362
rect 17550 10310 17562 10362
rect 17614 10310 17626 10362
rect 17678 10310 28317 10362
rect 28369 10310 28381 10362
rect 28433 10310 28445 10362
rect 28497 10310 28509 10362
rect 28561 10310 28573 10362
rect 28625 10310 39264 10362
rect 39316 10310 39328 10362
rect 39380 10310 39392 10362
rect 39444 10310 39456 10362
rect 39508 10310 39520 10362
rect 39572 10310 44896 10362
rect 1104 10288 44896 10310
rect 934 10208 940 10260
rect 992 10248 998 10260
rect 1765 10251 1823 10257
rect 1765 10248 1777 10251
rect 992 10220 1777 10248
rect 992 10208 998 10220
rect 1765 10217 1777 10220
rect 1811 10217 1823 10251
rect 1765 10211 1823 10217
rect 7926 10208 7932 10260
rect 7984 10208 7990 10260
rect 8386 10208 8392 10260
rect 8444 10208 8450 10260
rect 11422 10208 11428 10260
rect 11480 10248 11486 10260
rect 11701 10251 11759 10257
rect 11701 10248 11713 10251
rect 11480 10220 11713 10248
rect 11480 10208 11486 10220
rect 11701 10217 11713 10220
rect 11747 10217 11759 10251
rect 24578 10248 24584 10260
rect 11701 10211 11759 10217
rect 12406 10220 24584 10248
rect 8478 10140 8484 10192
rect 8536 10180 8542 10192
rect 10594 10180 10600 10192
rect 8536 10152 10600 10180
rect 8536 10140 8542 10152
rect 3142 10072 3148 10124
rect 3200 10072 3206 10124
rect 3237 10115 3295 10121
rect 3237 10081 3249 10115
rect 3283 10112 3295 10115
rect 3418 10112 3424 10124
rect 3283 10084 3424 10112
rect 3283 10081 3295 10084
rect 3237 10075 3295 10081
rect 3418 10072 3424 10084
rect 3476 10072 3482 10124
rect 9582 10072 9588 10124
rect 9640 10072 9646 10124
rect 9784 10121 9812 10152
rect 10594 10140 10600 10152
rect 10652 10180 10658 10192
rect 12406 10180 12434 10220
rect 24578 10208 24584 10220
rect 24636 10208 24642 10260
rect 24670 10208 24676 10260
rect 24728 10208 24734 10260
rect 32033 10251 32091 10257
rect 32033 10217 32045 10251
rect 32079 10248 32091 10251
rect 38010 10248 38016 10260
rect 32079 10220 38016 10248
rect 32079 10217 32091 10220
rect 32033 10211 32091 10217
rect 38010 10208 38016 10220
rect 38068 10208 38074 10260
rect 38197 10251 38255 10257
rect 38197 10217 38209 10251
rect 38243 10248 38255 10251
rect 38286 10248 38292 10260
rect 38243 10220 38292 10248
rect 38243 10217 38255 10220
rect 38197 10211 38255 10217
rect 38286 10208 38292 10220
rect 38344 10208 38350 10260
rect 38746 10208 38752 10260
rect 38804 10208 38810 10260
rect 42886 10208 42892 10260
rect 42944 10208 42950 10260
rect 10652 10152 12434 10180
rect 13725 10183 13783 10189
rect 10652 10140 10658 10152
rect 13725 10149 13737 10183
rect 13771 10180 13783 10183
rect 13998 10180 14004 10192
rect 13771 10152 14004 10180
rect 13771 10149 13783 10152
rect 13725 10143 13783 10149
rect 13998 10140 14004 10152
rect 14056 10140 14062 10192
rect 14921 10183 14979 10189
rect 14921 10149 14933 10183
rect 14967 10180 14979 10183
rect 16298 10180 16304 10192
rect 14967 10152 16304 10180
rect 14967 10149 14979 10152
rect 14921 10143 14979 10149
rect 16298 10140 16304 10152
rect 16356 10140 16362 10192
rect 16758 10140 16764 10192
rect 16816 10180 16822 10192
rect 17129 10183 17187 10189
rect 17129 10180 17141 10183
rect 16816 10152 17141 10180
rect 16816 10140 16822 10152
rect 17129 10149 17141 10152
rect 17175 10180 17187 10183
rect 17175 10152 19334 10180
rect 17175 10149 17187 10152
rect 17129 10143 17187 10149
rect 9769 10115 9827 10121
rect 9769 10081 9781 10115
rect 9815 10081 9827 10115
rect 9769 10075 9827 10081
rect 12406 10084 13492 10112
rect 1581 10047 1639 10053
rect 1581 10013 1593 10047
rect 1627 10044 1639 10047
rect 2774 10044 2780 10056
rect 1627 10016 2780 10044
rect 1627 10013 1639 10016
rect 1581 10007 1639 10013
rect 2774 10004 2780 10016
rect 2832 10004 2838 10056
rect 3326 10004 3332 10056
rect 3384 10044 3390 10056
rect 4525 10047 4583 10053
rect 4525 10044 4537 10047
rect 3384 10016 4537 10044
rect 3384 10004 3390 10016
rect 4525 10013 4537 10016
rect 4571 10013 4583 10047
rect 4525 10007 4583 10013
rect 4614 10004 4620 10056
rect 4672 10044 4678 10056
rect 4781 10047 4839 10053
rect 4781 10044 4793 10047
rect 4672 10016 4793 10044
rect 4672 10004 4678 10016
rect 4781 10013 4793 10016
rect 4827 10013 4839 10047
rect 4781 10007 4839 10013
rect 6549 10047 6607 10053
rect 6549 10013 6561 10047
rect 6595 10044 6607 10047
rect 7190 10044 7196 10056
rect 6595 10016 7196 10044
rect 6595 10013 6607 10016
rect 6549 10007 6607 10013
rect 7190 10004 7196 10016
rect 7248 10004 7254 10056
rect 8570 10004 8576 10056
rect 8628 10004 8634 10056
rect 6794 9979 6852 9985
rect 6794 9976 6806 9979
rect 5920 9948 6806 9976
rect 5920 9920 5948 9948
rect 6794 9945 6806 9948
rect 6840 9945 6852 9979
rect 6794 9939 6852 9945
rect 10410 9936 10416 9988
rect 10468 9976 10474 9988
rect 12406 9976 12434 10084
rect 13357 10047 13415 10053
rect 13357 10044 13369 10047
rect 10468 9948 12434 9976
rect 13280 10016 13369 10044
rect 10468 9936 10474 9948
rect 2222 9868 2228 9920
rect 2280 9908 2286 9920
rect 2685 9911 2743 9917
rect 2685 9908 2697 9911
rect 2280 9880 2697 9908
rect 2280 9868 2286 9880
rect 2685 9877 2697 9880
rect 2731 9877 2743 9911
rect 2685 9871 2743 9877
rect 3053 9911 3111 9917
rect 3053 9877 3065 9911
rect 3099 9908 3111 9911
rect 4338 9908 4344 9920
rect 3099 9880 4344 9908
rect 3099 9877 3111 9880
rect 3053 9871 3111 9877
rect 4338 9868 4344 9880
rect 4396 9868 4402 9920
rect 5902 9868 5908 9920
rect 5960 9868 5966 9920
rect 9125 9911 9183 9917
rect 9125 9877 9137 9911
rect 9171 9908 9183 9911
rect 9306 9908 9312 9920
rect 9171 9880 9312 9908
rect 9171 9877 9183 9880
rect 9125 9871 9183 9877
rect 9306 9868 9312 9880
rect 9364 9868 9370 9920
rect 9493 9911 9551 9917
rect 9493 9877 9505 9911
rect 9539 9908 9551 9911
rect 10042 9908 10048 9920
rect 9539 9880 10048 9908
rect 9539 9877 9551 9880
rect 9493 9871 9551 9877
rect 10042 9868 10048 9880
rect 10100 9868 10106 9920
rect 13280 9908 13308 10016
rect 13357 10013 13369 10016
rect 13403 10013 13415 10047
rect 13357 10007 13415 10013
rect 13464 9976 13492 10084
rect 13630 10072 13636 10124
rect 13688 10112 13694 10124
rect 13688 10084 14780 10112
rect 13688 10072 13694 10084
rect 13541 10047 13599 10053
rect 13541 10013 13553 10047
rect 13587 10044 13599 10047
rect 14274 10044 14280 10056
rect 13587 10016 14280 10044
rect 13587 10013 13599 10016
rect 13541 10007 13599 10013
rect 14274 10004 14280 10016
rect 14332 10004 14338 10056
rect 14642 10004 14648 10056
rect 14700 10004 14706 10056
rect 14752 10053 14780 10084
rect 18414 10072 18420 10124
rect 18472 10112 18478 10124
rect 18509 10115 18567 10121
rect 18509 10112 18521 10115
rect 18472 10084 18521 10112
rect 18472 10072 18478 10084
rect 18509 10081 18521 10084
rect 18555 10081 18567 10115
rect 18509 10075 18567 10081
rect 18693 10115 18751 10121
rect 18693 10081 18705 10115
rect 18739 10112 18751 10115
rect 19150 10112 19156 10124
rect 18739 10084 19156 10112
rect 18739 10081 18751 10084
rect 18693 10075 18751 10081
rect 19150 10072 19156 10084
rect 19208 10072 19214 10124
rect 19306 10112 19334 10152
rect 22738 10140 22744 10192
rect 22796 10180 22802 10192
rect 22925 10183 22983 10189
rect 22925 10180 22937 10183
rect 22796 10152 22937 10180
rect 22796 10140 22802 10152
rect 22925 10149 22937 10152
rect 22971 10149 22983 10183
rect 24946 10180 24952 10192
rect 22925 10143 22983 10149
rect 23492 10152 24952 10180
rect 21453 10115 21511 10121
rect 19306 10084 21128 10112
rect 14737 10047 14795 10053
rect 14737 10013 14749 10047
rect 14783 10013 14795 10047
rect 14737 10007 14795 10013
rect 17954 10004 17960 10056
rect 18012 10044 18018 10056
rect 19429 10047 19487 10053
rect 19429 10044 19441 10047
rect 18012 10016 19441 10044
rect 18012 10004 18018 10016
rect 19429 10013 19441 10016
rect 19475 10044 19487 10047
rect 21100 10044 21128 10084
rect 21453 10081 21465 10115
rect 21499 10112 21511 10115
rect 23492 10112 23520 10152
rect 24946 10140 24952 10152
rect 25004 10140 25010 10192
rect 21499 10084 23520 10112
rect 21499 10081 21511 10084
rect 21453 10075 21511 10081
rect 24854 10072 24860 10124
rect 24912 10112 24918 10124
rect 25685 10115 25743 10121
rect 25685 10112 25697 10115
rect 24912 10084 25697 10112
rect 24912 10072 24918 10084
rect 25685 10081 25697 10084
rect 25731 10081 25743 10115
rect 25685 10075 25743 10081
rect 31846 10072 31852 10124
rect 31904 10072 31910 10124
rect 36262 10072 36268 10124
rect 36320 10112 36326 10124
rect 36814 10112 36820 10124
rect 36320 10084 36820 10112
rect 36320 10072 36326 10084
rect 36814 10072 36820 10084
rect 36872 10072 36878 10124
rect 21174 10044 21180 10056
rect 19475 10016 19656 10044
rect 21100 10016 21180 10044
rect 19475 10013 19487 10016
rect 19429 10007 19487 10013
rect 15654 9976 15660 9988
rect 13464 9948 15660 9976
rect 15654 9936 15660 9948
rect 15712 9936 15718 9988
rect 13814 9908 13820 9920
rect 13280 9880 13820 9908
rect 13814 9868 13820 9880
rect 13872 9908 13878 9920
rect 14366 9908 14372 9920
rect 13872 9880 14372 9908
rect 13872 9868 13878 9880
rect 14366 9868 14372 9880
rect 14424 9908 14430 9920
rect 14642 9908 14648 9920
rect 14424 9880 14648 9908
rect 14424 9868 14430 9880
rect 14642 9868 14648 9880
rect 14700 9868 14706 9920
rect 18046 9868 18052 9920
rect 18104 9868 18110 9920
rect 18414 9868 18420 9920
rect 18472 9868 18478 9920
rect 19518 9868 19524 9920
rect 19576 9868 19582 9920
rect 19628 9908 19656 10016
rect 21174 10004 21180 10016
rect 21232 10004 21238 10056
rect 23569 10047 23627 10053
rect 23569 10013 23581 10047
rect 23615 10044 23627 10047
rect 24581 10047 24639 10053
rect 24581 10044 24593 10047
rect 23615 10016 24593 10044
rect 23615 10013 23627 10016
rect 23569 10007 23627 10013
rect 24581 10013 24593 10016
rect 24627 10044 24639 10047
rect 25498 10044 25504 10056
rect 24627 10016 25504 10044
rect 24627 10013 24639 10016
rect 24581 10007 24639 10013
rect 22186 9936 22192 9988
rect 22244 9936 22250 9988
rect 23584 9976 23612 10007
rect 25498 10004 25504 10016
rect 25556 10004 25562 10056
rect 28994 10004 29000 10056
rect 29052 10044 29058 10056
rect 29730 10044 29736 10056
rect 29052 10016 29736 10044
rect 29052 10004 29058 10016
rect 29730 10004 29736 10016
rect 29788 10004 29794 10056
rect 29822 10004 29828 10056
rect 29880 10044 29886 10056
rect 29989 10047 30047 10053
rect 29989 10044 30001 10047
rect 29880 10016 30001 10044
rect 29880 10004 29886 10016
rect 29989 10013 30001 10016
rect 30035 10044 30047 10047
rect 30926 10044 30932 10056
rect 30035 10016 30932 10044
rect 30035 10013 30047 10016
rect 29989 10007 30047 10013
rect 30926 10004 30932 10016
rect 30984 10004 30990 10056
rect 31754 10004 31760 10056
rect 31812 10004 31818 10056
rect 32674 10004 32680 10056
rect 32732 10004 32738 10056
rect 32766 10004 32772 10056
rect 32824 10004 32830 10056
rect 38654 10004 38660 10056
rect 38712 10004 38718 10056
rect 42797 10047 42855 10053
rect 42797 10013 42809 10047
rect 42843 10044 42855 10047
rect 43438 10044 43444 10056
rect 42843 10016 43444 10044
rect 42843 10013 42855 10016
rect 42797 10007 42855 10013
rect 43438 10004 43444 10016
rect 43496 10004 43502 10056
rect 22756 9948 23612 9976
rect 25952 9979 26010 9985
rect 22756 9908 22784 9948
rect 25952 9945 25964 9979
rect 25998 9976 26010 9979
rect 26418 9976 26424 9988
rect 25998 9948 26424 9976
rect 25998 9945 26010 9948
rect 25952 9939 26010 9945
rect 26418 9936 26424 9948
rect 26476 9936 26482 9988
rect 36722 9936 36728 9988
rect 36780 9976 36786 9988
rect 37062 9979 37120 9985
rect 37062 9976 37074 9979
rect 36780 9948 37074 9976
rect 36780 9936 36786 9948
rect 37062 9945 37074 9948
rect 37108 9945 37120 9979
rect 37062 9939 37120 9945
rect 19628 9880 22784 9908
rect 23566 9868 23572 9920
rect 23624 9908 23630 9920
rect 23661 9911 23719 9917
rect 23661 9908 23673 9911
rect 23624 9880 23673 9908
rect 23624 9868 23630 9880
rect 23661 9877 23673 9880
rect 23707 9877 23719 9911
rect 23661 9871 23719 9877
rect 25314 9868 25320 9920
rect 25372 9908 25378 9920
rect 27065 9911 27123 9917
rect 27065 9908 27077 9911
rect 25372 9880 27077 9908
rect 25372 9868 25378 9880
rect 27065 9877 27077 9880
rect 27111 9877 27123 9911
rect 27065 9871 27123 9877
rect 30650 9868 30656 9920
rect 30708 9908 30714 9920
rect 31113 9911 31171 9917
rect 31113 9908 31125 9911
rect 30708 9880 31125 9908
rect 30708 9868 30714 9880
rect 31113 9877 31125 9880
rect 31159 9877 31171 9911
rect 31113 9871 31171 9877
rect 32490 9868 32496 9920
rect 32548 9908 32554 9920
rect 32953 9911 33011 9917
rect 32953 9908 32965 9911
rect 32548 9880 32965 9908
rect 32548 9868 32554 9880
rect 32953 9877 32965 9880
rect 32999 9877 33011 9911
rect 32953 9871 33011 9877
rect 1104 9818 45051 9840
rect 1104 9766 11896 9818
rect 11948 9766 11960 9818
rect 12012 9766 12024 9818
rect 12076 9766 12088 9818
rect 12140 9766 12152 9818
rect 12204 9766 22843 9818
rect 22895 9766 22907 9818
rect 22959 9766 22971 9818
rect 23023 9766 23035 9818
rect 23087 9766 23099 9818
rect 23151 9766 33790 9818
rect 33842 9766 33854 9818
rect 33906 9766 33918 9818
rect 33970 9766 33982 9818
rect 34034 9766 34046 9818
rect 34098 9766 44737 9818
rect 44789 9766 44801 9818
rect 44853 9766 44865 9818
rect 44917 9766 44929 9818
rect 44981 9766 44993 9818
rect 45045 9766 45051 9818
rect 1104 9744 45051 9766
rect 4614 9664 4620 9716
rect 4672 9704 4678 9716
rect 4709 9707 4767 9713
rect 4709 9704 4721 9707
rect 4672 9676 4721 9704
rect 4672 9664 4678 9676
rect 4709 9673 4721 9676
rect 4755 9673 4767 9707
rect 4709 9667 4767 9673
rect 6086 9664 6092 9716
rect 6144 9704 6150 9716
rect 13814 9704 13820 9716
rect 6144 9676 13820 9704
rect 6144 9664 6150 9676
rect 13814 9664 13820 9676
rect 13872 9664 13878 9716
rect 14274 9664 14280 9716
rect 14332 9664 14338 9716
rect 22646 9664 22652 9716
rect 22704 9704 22710 9716
rect 25130 9704 25136 9716
rect 22704 9676 25136 9704
rect 22704 9664 22710 9676
rect 2884 9608 5488 9636
rect 2222 9528 2228 9580
rect 2280 9528 2286 9580
rect 2884 9577 2912 9608
rect 2869 9571 2927 9577
rect 2869 9537 2881 9571
rect 2915 9537 2927 9571
rect 2869 9531 2927 9537
rect 3326 9528 3332 9580
rect 3384 9528 3390 9580
rect 3596 9571 3654 9577
rect 3596 9537 3608 9571
rect 3642 9568 3654 9571
rect 3642 9540 5304 9568
rect 3642 9537 3654 9540
rect 3596 9531 3654 9537
rect 4522 9392 4528 9444
rect 4580 9432 4586 9444
rect 5169 9435 5227 9441
rect 5169 9432 5181 9435
rect 4580 9404 5181 9432
rect 4580 9392 4586 9404
rect 5169 9401 5181 9404
rect 5215 9401 5227 9435
rect 5276 9432 5304 9540
rect 5460 9500 5488 9608
rect 5534 9596 5540 9648
rect 5592 9596 5598 9648
rect 9122 9636 9128 9648
rect 7208 9608 9128 9636
rect 7208 9580 7236 9608
rect 9122 9596 9128 9608
rect 9180 9596 9186 9648
rect 15194 9645 15200 9648
rect 15188 9636 15200 9645
rect 12912 9608 14964 9636
rect 15155 9608 15200 9636
rect 12912 9580 12940 9608
rect 5629 9571 5687 9577
rect 5629 9537 5641 9571
rect 5675 9568 5687 9571
rect 6270 9568 6276 9580
rect 5675 9540 6276 9568
rect 5675 9537 5687 9540
rect 5629 9531 5687 9537
rect 6270 9528 6276 9540
rect 6328 9528 6334 9580
rect 7190 9528 7196 9580
rect 7248 9528 7254 9580
rect 7460 9571 7518 9577
rect 7460 9537 7472 9571
rect 7506 9568 7518 9571
rect 7926 9568 7932 9580
rect 7506 9540 7932 9568
rect 7506 9537 7518 9540
rect 7460 9531 7518 9537
rect 7926 9528 7932 9540
rect 7984 9528 7990 9580
rect 9677 9571 9735 9577
rect 9677 9537 9689 9571
rect 9723 9568 9735 9571
rect 9766 9568 9772 9580
rect 9723 9540 9772 9568
rect 9723 9537 9735 9540
rect 9677 9531 9735 9537
rect 9766 9528 9772 9540
rect 9824 9528 9830 9580
rect 9944 9571 10002 9577
rect 9944 9537 9956 9571
rect 9990 9568 10002 9571
rect 11606 9568 11612 9580
rect 9990 9540 11612 9568
rect 9990 9537 10002 9540
rect 9944 9531 10002 9537
rect 11606 9528 11612 9540
rect 11664 9528 11670 9580
rect 11885 9571 11943 9577
rect 11885 9537 11897 9571
rect 11931 9537 11943 9571
rect 11885 9531 11943 9537
rect 5534 9500 5540 9512
rect 5460 9472 5540 9500
rect 5534 9460 5540 9472
rect 5592 9460 5598 9512
rect 5810 9460 5816 9512
rect 5868 9460 5874 9512
rect 10686 9460 10692 9512
rect 10744 9500 10750 9512
rect 11900 9500 11928 9531
rect 12894 9528 12900 9580
rect 12952 9528 12958 9580
rect 13170 9577 13176 9580
rect 13164 9568 13176 9577
rect 13131 9540 13176 9568
rect 13164 9531 13176 9540
rect 13170 9528 13176 9531
rect 13228 9528 13234 9580
rect 14936 9577 14964 9608
rect 15188 9599 15200 9608
rect 15194 9596 15200 9599
rect 15252 9596 15258 9648
rect 18046 9636 18052 9648
rect 17144 9608 18052 9636
rect 17144 9577 17172 9608
rect 18046 9596 18052 9608
rect 18104 9596 18110 9648
rect 19518 9596 19524 9648
rect 19576 9596 19582 9648
rect 22738 9596 22744 9648
rect 22796 9636 22802 9648
rect 22833 9639 22891 9645
rect 22833 9636 22845 9639
rect 22796 9608 22845 9636
rect 22796 9596 22802 9608
rect 22833 9605 22845 9608
rect 22879 9605 22891 9639
rect 22833 9599 22891 9605
rect 23566 9596 23572 9648
rect 23624 9596 23630 9648
rect 24596 9645 24624 9676
rect 25130 9664 25136 9676
rect 25188 9664 25194 9716
rect 26418 9664 26424 9716
rect 26476 9664 26482 9716
rect 31294 9664 31300 9716
rect 31352 9704 31358 9716
rect 31665 9707 31723 9713
rect 31665 9704 31677 9707
rect 31352 9676 31677 9704
rect 31352 9664 31358 9676
rect 31665 9673 31677 9676
rect 31711 9673 31723 9707
rect 31665 9667 31723 9673
rect 36722 9664 36728 9716
rect 36780 9664 36786 9716
rect 24581 9639 24639 9645
rect 24581 9605 24593 9639
rect 24627 9605 24639 9639
rect 24581 9599 24639 9605
rect 25314 9596 25320 9648
rect 25372 9636 25378 9648
rect 26145 9639 26203 9645
rect 26145 9636 26157 9639
rect 25372 9608 26157 9636
rect 25372 9596 25378 9608
rect 26145 9605 26157 9608
rect 26191 9605 26203 9639
rect 28994 9636 29000 9648
rect 26145 9599 26203 9605
rect 28460 9608 29000 9636
rect 14921 9571 14979 9577
rect 14921 9537 14933 9571
rect 14967 9537 14979 9571
rect 14921 9531 14979 9537
rect 17129 9571 17187 9577
rect 17129 9537 17141 9571
rect 17175 9537 17187 9571
rect 17129 9531 17187 9537
rect 17589 9571 17647 9577
rect 17589 9537 17601 9571
rect 17635 9568 17647 9571
rect 17954 9568 17960 9580
rect 17635 9540 17960 9568
rect 17635 9537 17647 9540
rect 17589 9531 17647 9537
rect 17954 9528 17960 9540
rect 18012 9528 18018 9580
rect 18601 9571 18659 9577
rect 18601 9537 18613 9571
rect 18647 9568 18659 9571
rect 18690 9568 18696 9580
rect 18647 9540 18696 9568
rect 18647 9537 18659 9540
rect 18601 9531 18659 9537
rect 18690 9528 18696 9540
rect 18748 9528 18754 9580
rect 22554 9528 22560 9580
rect 22612 9528 22618 9580
rect 25409 9571 25467 9577
rect 25409 9537 25421 9571
rect 25455 9568 25467 9571
rect 25590 9568 25596 9580
rect 25455 9540 25596 9568
rect 25455 9537 25467 9540
rect 25409 9531 25467 9537
rect 25590 9528 25596 9540
rect 25648 9528 25654 9580
rect 25774 9528 25780 9580
rect 25832 9568 25838 9580
rect 25869 9571 25927 9577
rect 25869 9568 25881 9571
rect 25832 9540 25881 9568
rect 25832 9528 25838 9540
rect 25869 9537 25881 9540
rect 25915 9537 25927 9571
rect 25869 9531 25927 9537
rect 26053 9571 26111 9577
rect 26053 9537 26065 9571
rect 26099 9537 26111 9571
rect 26053 9531 26111 9537
rect 10744 9472 11928 9500
rect 10744 9460 10750 9472
rect 16758 9460 16764 9512
rect 16816 9500 16822 9512
rect 18233 9503 18291 9509
rect 18233 9500 18245 9503
rect 16816 9472 18245 9500
rect 16816 9460 16822 9472
rect 18233 9469 18245 9472
rect 18279 9469 18291 9503
rect 18233 9463 18291 9469
rect 6914 9432 6920 9444
rect 5276 9404 6920 9432
rect 5169 9395 5227 9401
rect 6914 9392 6920 9404
rect 6972 9392 6978 9444
rect 10962 9392 10968 9444
rect 11020 9432 11026 9444
rect 11057 9435 11115 9441
rect 11057 9432 11069 9435
rect 11020 9404 11069 9432
rect 11020 9392 11026 9404
rect 11057 9401 11069 9404
rect 11103 9401 11115 9435
rect 11057 9395 11115 9401
rect 16301 9435 16359 9441
rect 16301 9401 16313 9435
rect 16347 9432 16359 9435
rect 16390 9432 16396 9444
rect 16347 9404 16396 9432
rect 16347 9401 16359 9404
rect 16301 9395 16359 9401
rect 16390 9392 16396 9404
rect 16448 9392 16454 9444
rect 2038 9324 2044 9376
rect 2096 9324 2102 9376
rect 2685 9367 2743 9373
rect 2685 9333 2697 9367
rect 2731 9364 2743 9367
rect 4246 9364 4252 9376
rect 2731 9336 4252 9364
rect 2731 9333 2743 9336
rect 2685 9327 2743 9333
rect 4246 9324 4252 9336
rect 4304 9324 4310 9376
rect 8294 9324 8300 9376
rect 8352 9364 8358 9376
rect 8573 9367 8631 9373
rect 8573 9364 8585 9367
rect 8352 9336 8585 9364
rect 8352 9324 8358 9336
rect 8573 9333 8585 9336
rect 8619 9333 8631 9367
rect 8573 9327 8631 9333
rect 10318 9324 10324 9376
rect 10376 9364 10382 9376
rect 11701 9367 11759 9373
rect 11701 9364 11713 9367
rect 10376 9336 11713 9364
rect 10376 9324 10382 9336
rect 11701 9333 11713 9336
rect 11747 9333 11759 9367
rect 11701 9327 11759 9333
rect 16942 9324 16948 9376
rect 17000 9324 17006 9376
rect 17681 9367 17739 9373
rect 17681 9333 17693 9367
rect 17727 9364 17739 9367
rect 17770 9364 17776 9376
rect 17727 9336 17776 9364
rect 17727 9333 17739 9336
rect 17681 9327 17739 9333
rect 17770 9324 17776 9336
rect 17828 9324 17834 9376
rect 20027 9367 20085 9373
rect 20027 9333 20039 9367
rect 20073 9364 20085 9367
rect 20714 9364 20720 9376
rect 20073 9336 20720 9364
rect 20073 9333 20085 9336
rect 20027 9327 20085 9333
rect 20714 9324 20720 9336
rect 20772 9324 20778 9376
rect 25038 9324 25044 9376
rect 25096 9364 25102 9376
rect 25225 9367 25283 9373
rect 25225 9364 25237 9367
rect 25096 9336 25237 9364
rect 25096 9324 25102 9336
rect 25225 9333 25237 9336
rect 25271 9333 25283 9367
rect 26068 9364 26096 9531
rect 26234 9528 26240 9580
rect 26292 9528 26298 9580
rect 28460 9577 28488 9608
rect 28994 9596 29000 9608
rect 29052 9596 29058 9648
rect 29178 9596 29184 9648
rect 29236 9596 29242 9648
rect 30650 9596 30656 9648
rect 30708 9596 30714 9648
rect 32766 9636 32772 9648
rect 31726 9608 32772 9636
rect 28445 9571 28503 9577
rect 28445 9537 28457 9571
rect 28491 9537 28503 9571
rect 31573 9571 31631 9577
rect 31573 9568 31585 9571
rect 28445 9531 28503 9537
rect 30208 9540 31585 9568
rect 27614 9460 27620 9512
rect 27672 9500 27678 9512
rect 30208 9509 30236 9540
rect 31573 9537 31585 9540
rect 31619 9568 31631 9571
rect 31726 9568 31754 9608
rect 32766 9596 32772 9608
rect 32824 9596 32830 9648
rect 33502 9636 33508 9648
rect 32968 9608 33508 9636
rect 31619 9540 31754 9568
rect 31619 9537 31631 9540
rect 31573 9531 31631 9537
rect 32490 9528 32496 9580
rect 32548 9528 32554 9580
rect 32968 9577 32996 9608
rect 33502 9596 33508 9608
rect 33560 9596 33566 9648
rect 33686 9596 33692 9648
rect 33744 9596 33750 9648
rect 44082 9636 44088 9648
rect 35636 9608 44088 9636
rect 32953 9571 33011 9577
rect 32953 9537 32965 9571
rect 32999 9537 33011 9571
rect 35636 9568 35664 9608
rect 44082 9596 44088 9608
rect 44140 9596 44146 9648
rect 32953 9531 33011 9537
rect 34900 9540 35664 9568
rect 35805 9571 35863 9577
rect 28721 9503 28779 9509
rect 28721 9500 28733 9503
rect 27672 9472 28733 9500
rect 27672 9460 27678 9472
rect 28721 9469 28733 9472
rect 28767 9469 28779 9503
rect 28721 9463 28779 9469
rect 30193 9503 30251 9509
rect 30193 9469 30205 9503
rect 30239 9469 30251 9503
rect 33229 9503 33287 9509
rect 33229 9500 33241 9503
rect 30193 9463 30251 9469
rect 32324 9472 33241 9500
rect 30926 9392 30932 9444
rect 30984 9392 30990 9444
rect 32324 9441 32352 9472
rect 33229 9469 33241 9472
rect 33275 9500 33287 9503
rect 34900 9500 34928 9540
rect 35805 9537 35817 9571
rect 35851 9568 35863 9571
rect 36354 9568 36360 9580
rect 35851 9540 36360 9568
rect 35851 9537 35863 9540
rect 35805 9531 35863 9537
rect 36354 9528 36360 9540
rect 36412 9528 36418 9580
rect 36906 9528 36912 9580
rect 36964 9528 36970 9580
rect 37734 9528 37740 9580
rect 37792 9528 37798 9580
rect 33275 9472 34928 9500
rect 33275 9469 33287 9472
rect 33229 9463 33287 9469
rect 34974 9460 34980 9512
rect 35032 9460 35038 9512
rect 35897 9503 35955 9509
rect 35897 9500 35909 9503
rect 35084 9472 35909 9500
rect 32309 9435 32367 9441
rect 32309 9401 32321 9435
rect 32355 9401 32367 9435
rect 35084 9432 35112 9472
rect 35897 9469 35909 9472
rect 35943 9469 35955 9503
rect 35897 9463 35955 9469
rect 35989 9503 36047 9509
rect 35989 9469 36001 9503
rect 36035 9469 36047 9503
rect 35989 9463 36047 9469
rect 32309 9395 32367 9401
rect 34256 9404 35112 9432
rect 29822 9364 29828 9376
rect 26068 9336 29828 9364
rect 25225 9327 25283 9333
rect 29822 9324 29828 9336
rect 29880 9324 29886 9376
rect 31113 9367 31171 9373
rect 31113 9333 31125 9367
rect 31159 9364 31171 9367
rect 31662 9364 31668 9376
rect 31159 9336 31668 9364
rect 31159 9333 31171 9336
rect 31113 9327 31171 9333
rect 31662 9324 31668 9336
rect 31720 9324 31726 9376
rect 32950 9324 32956 9376
rect 33008 9364 33014 9376
rect 34256 9364 34284 9404
rect 35710 9392 35716 9444
rect 35768 9432 35774 9444
rect 36004 9432 36032 9463
rect 35768 9404 36032 9432
rect 35768 9392 35774 9404
rect 33008 9336 34284 9364
rect 33008 9324 33014 9336
rect 34330 9324 34336 9376
rect 34388 9364 34394 9376
rect 35437 9367 35495 9373
rect 35437 9364 35449 9367
rect 34388 9336 35449 9364
rect 34388 9324 34394 9336
rect 35437 9333 35449 9336
rect 35483 9333 35495 9367
rect 35437 9327 35495 9333
rect 37550 9324 37556 9376
rect 37608 9324 37614 9376
rect 1104 9274 44896 9296
rect 1104 9222 6423 9274
rect 6475 9222 6487 9274
rect 6539 9222 6551 9274
rect 6603 9222 6615 9274
rect 6667 9222 6679 9274
rect 6731 9222 17370 9274
rect 17422 9222 17434 9274
rect 17486 9222 17498 9274
rect 17550 9222 17562 9274
rect 17614 9222 17626 9274
rect 17678 9222 28317 9274
rect 28369 9222 28381 9274
rect 28433 9222 28445 9274
rect 28497 9222 28509 9274
rect 28561 9222 28573 9274
rect 28625 9222 39264 9274
rect 39316 9222 39328 9274
rect 39380 9222 39392 9274
rect 39444 9222 39456 9274
rect 39508 9222 39520 9274
rect 39572 9222 44896 9274
rect 1104 9200 44896 9222
rect 7837 9163 7895 9169
rect 7837 9129 7849 9163
rect 7883 9160 7895 9163
rect 10686 9160 10692 9172
rect 7883 9132 10692 9160
rect 7883 9129 7895 9132
rect 7837 9123 7895 9129
rect 10686 9120 10692 9132
rect 10744 9120 10750 9172
rect 11606 9120 11612 9172
rect 11664 9120 11670 9172
rect 13906 9120 13912 9172
rect 13964 9160 13970 9172
rect 14277 9163 14335 9169
rect 14277 9160 14289 9163
rect 13964 9132 14289 9160
rect 13964 9120 13970 9132
rect 14277 9129 14289 9132
rect 14323 9129 14335 9163
rect 14277 9123 14335 9129
rect 16114 9120 16120 9172
rect 16172 9160 16178 9172
rect 17954 9160 17960 9172
rect 16172 9132 17960 9160
rect 16172 9120 16178 9132
rect 17954 9120 17960 9132
rect 18012 9120 18018 9172
rect 18414 9120 18420 9172
rect 18472 9160 18478 9172
rect 18831 9163 18889 9169
rect 18831 9160 18843 9163
rect 18472 9132 18843 9160
rect 18472 9120 18478 9132
rect 18831 9129 18843 9132
rect 18877 9160 18889 9163
rect 19058 9160 19064 9172
rect 18877 9132 19064 9160
rect 18877 9129 18889 9132
rect 18831 9123 18889 9129
rect 19058 9120 19064 9132
rect 19116 9120 19122 9172
rect 19426 9120 19432 9172
rect 19484 9120 19490 9172
rect 32950 9160 32956 9172
rect 20824 9132 32956 9160
rect 2685 9095 2743 9101
rect 2685 9061 2697 9095
rect 2731 9061 2743 9095
rect 13630 9092 13636 9104
rect 2685 9055 2743 9061
rect 11164 9064 13636 9092
rect 2225 8959 2283 8965
rect 2225 8925 2237 8959
rect 2271 8956 2283 8959
rect 2700 8956 2728 9055
rect 3329 9027 3387 9033
rect 3329 8993 3341 9027
rect 3375 9024 3387 9027
rect 3418 9024 3424 9036
rect 3375 8996 3424 9024
rect 3375 8993 3387 8996
rect 3329 8987 3387 8993
rect 3418 8984 3424 8996
rect 3476 9024 3482 9036
rect 5810 9024 5816 9036
rect 3476 8996 5816 9024
rect 3476 8984 3482 8996
rect 5810 8984 5816 8996
rect 5868 9024 5874 9036
rect 8478 9024 8484 9036
rect 5868 8996 8484 9024
rect 5868 8984 5874 8996
rect 8478 8984 8484 8996
rect 8536 8984 8542 9036
rect 9766 8984 9772 9036
rect 9824 8984 9830 9036
rect 2271 8928 2728 8956
rect 4065 8959 4123 8965
rect 2271 8925 2283 8928
rect 2225 8919 2283 8925
rect 4065 8925 4077 8959
rect 4111 8956 4123 8959
rect 5350 8956 5356 8968
rect 4111 8928 5356 8956
rect 4111 8925 4123 8928
rect 4065 8919 4123 8925
rect 5350 8916 5356 8928
rect 5408 8916 5414 8968
rect 5626 8916 5632 8968
rect 5684 8916 5690 8968
rect 8202 8916 8208 8968
rect 8260 8956 8266 8968
rect 8297 8959 8355 8965
rect 8297 8956 8309 8959
rect 8260 8928 8309 8956
rect 8260 8916 8266 8928
rect 8297 8925 8309 8928
rect 8343 8925 8355 8959
rect 8297 8919 8355 8925
rect 9306 8916 9312 8968
rect 9364 8916 9370 8968
rect 10036 8959 10094 8965
rect 10036 8925 10048 8959
rect 10082 8956 10094 8959
rect 10318 8956 10324 8968
rect 10082 8928 10324 8956
rect 10082 8925 10094 8928
rect 10036 8919 10094 8925
rect 10318 8916 10324 8928
rect 10376 8916 10382 8968
rect 3053 8891 3111 8897
rect 3053 8857 3065 8891
rect 3099 8888 3111 8891
rect 3234 8888 3240 8900
rect 3099 8860 3240 8888
rect 3099 8857 3111 8860
rect 3053 8851 3111 8857
rect 3234 8848 3240 8860
rect 3292 8848 3298 8900
rect 11164 8888 11192 9064
rect 13630 9052 13636 9064
rect 13688 9052 13694 9104
rect 14921 9027 14979 9033
rect 14921 8993 14933 9027
rect 14967 9024 14979 9027
rect 15470 9024 15476 9036
rect 14967 8996 15476 9024
rect 14967 8993 14979 8996
rect 14921 8987 14979 8993
rect 15470 8984 15476 8996
rect 15528 8984 15534 9036
rect 16942 8984 16948 9036
rect 17000 9024 17006 9036
rect 17405 9027 17463 9033
rect 17405 9024 17417 9027
rect 17000 8996 17417 9024
rect 17000 8984 17006 8996
rect 17405 8993 17417 8996
rect 17451 8993 17463 9027
rect 17405 8987 17463 8993
rect 19150 8984 19156 9036
rect 19208 9024 19214 9036
rect 19981 9027 20039 9033
rect 19981 9024 19993 9027
rect 19208 8996 19993 9024
rect 19208 8984 19214 8996
rect 19981 8993 19993 8996
rect 20027 8993 20039 9027
rect 19981 8987 20039 8993
rect 11790 8916 11796 8968
rect 11848 8916 11854 8968
rect 13170 8916 13176 8968
rect 13228 8956 13234 8968
rect 14645 8959 14703 8965
rect 14645 8956 14657 8959
rect 13228 8928 14657 8956
rect 13228 8916 13234 8928
rect 14645 8925 14657 8928
rect 14691 8925 14703 8959
rect 14645 8919 14703 8925
rect 16393 8959 16451 8965
rect 16393 8925 16405 8959
rect 16439 8956 16451 8959
rect 16850 8956 16856 8968
rect 16439 8928 16856 8956
rect 16439 8925 16451 8928
rect 16393 8919 16451 8925
rect 8220 8860 11192 8888
rect 14660 8888 14688 8919
rect 16850 8916 16856 8928
rect 16908 8916 16914 8968
rect 17037 8959 17095 8965
rect 17037 8925 17049 8959
rect 17083 8956 17095 8959
rect 17126 8956 17132 8968
rect 17083 8928 17132 8956
rect 17083 8925 17095 8928
rect 17037 8919 17095 8925
rect 17126 8916 17132 8928
rect 17184 8916 17190 8968
rect 14660 8860 16620 8888
rect 2041 8823 2099 8829
rect 2041 8789 2053 8823
rect 2087 8820 2099 8823
rect 2222 8820 2228 8832
rect 2087 8792 2228 8820
rect 2087 8789 2099 8792
rect 2041 8783 2099 8789
rect 2222 8780 2228 8792
rect 2280 8780 2286 8832
rect 3145 8823 3203 8829
rect 3145 8789 3157 8823
rect 3191 8820 3203 8823
rect 4617 8823 4675 8829
rect 4617 8820 4629 8823
rect 3191 8792 4629 8820
rect 3191 8789 3203 8792
rect 3145 8783 3203 8789
rect 4617 8789 4629 8792
rect 4663 8789 4675 8823
rect 4617 8783 4675 8789
rect 6822 8780 6828 8832
rect 6880 8820 6886 8832
rect 8220 8829 8248 8860
rect 6917 8823 6975 8829
rect 6917 8820 6929 8823
rect 6880 8792 6929 8820
rect 6880 8780 6886 8792
rect 6917 8789 6929 8792
rect 6963 8789 6975 8823
rect 6917 8783 6975 8789
rect 8205 8823 8263 8829
rect 8205 8789 8217 8823
rect 8251 8789 8263 8823
rect 8205 8783 8263 8789
rect 8938 8780 8944 8832
rect 8996 8820 9002 8832
rect 11164 8829 11192 8860
rect 9125 8823 9183 8829
rect 9125 8820 9137 8823
rect 8996 8792 9137 8820
rect 8996 8780 9002 8792
rect 9125 8789 9137 8792
rect 9171 8789 9183 8823
rect 9125 8783 9183 8789
rect 11149 8823 11207 8829
rect 11149 8789 11161 8823
rect 11195 8789 11207 8823
rect 11149 8783 11207 8789
rect 14734 8780 14740 8832
rect 14792 8780 14798 8832
rect 16206 8780 16212 8832
rect 16264 8780 16270 8832
rect 16592 8820 16620 8860
rect 17770 8848 17776 8900
rect 17828 8848 17834 8900
rect 19797 8891 19855 8897
rect 19797 8857 19809 8891
rect 19843 8888 19855 8891
rect 20714 8888 20720 8900
rect 19843 8860 20720 8888
rect 19843 8857 19855 8860
rect 19797 8851 19855 8857
rect 20714 8848 20720 8860
rect 20772 8848 20778 8900
rect 19889 8823 19947 8829
rect 19889 8820 19901 8823
rect 16592 8792 19901 8820
rect 19889 8789 19901 8792
rect 19935 8820 19947 8823
rect 20824 8820 20852 9132
rect 32950 9120 32956 9132
rect 33008 9120 33014 9172
rect 33045 9163 33103 9169
rect 33045 9129 33057 9163
rect 33091 9160 33103 9163
rect 33686 9160 33692 9172
rect 33091 9132 33692 9160
rect 33091 9129 33103 9132
rect 33045 9123 33103 9129
rect 33686 9120 33692 9132
rect 33744 9120 33750 9172
rect 34146 9120 34152 9172
rect 34204 9120 34210 9172
rect 35710 9160 35716 9172
rect 34440 9132 35716 9160
rect 20990 9052 20996 9104
rect 21048 9092 21054 9104
rect 21910 9092 21916 9104
rect 21048 9064 21916 9092
rect 21048 9052 21054 9064
rect 21910 9052 21916 9064
rect 21968 9092 21974 9104
rect 22005 9095 22063 9101
rect 22005 9092 22017 9095
rect 21968 9064 22017 9092
rect 21968 9052 21974 9064
rect 22005 9061 22017 9064
rect 22051 9061 22063 9095
rect 22005 9055 22063 9061
rect 27249 9095 27307 9101
rect 27249 9061 27261 9095
rect 27295 9092 27307 9095
rect 27522 9092 27528 9104
rect 27295 9064 27528 9092
rect 27295 9061 27307 9064
rect 27249 9055 27307 9061
rect 27522 9052 27528 9064
rect 27580 9052 27586 9104
rect 29089 9095 29147 9101
rect 29089 9061 29101 9095
rect 29135 9092 29147 9095
rect 29178 9092 29184 9104
rect 29135 9064 29184 9092
rect 29135 9061 29147 9064
rect 29089 9055 29147 9061
rect 29178 9052 29184 9064
rect 29236 9052 29242 9104
rect 29822 9052 29828 9104
rect 29880 9052 29886 9104
rect 32401 9095 32459 9101
rect 32401 9061 32413 9095
rect 32447 9092 32459 9095
rect 32674 9092 32680 9104
rect 32447 9064 32680 9092
rect 32447 9061 32459 9064
rect 32401 9055 32459 9061
rect 32674 9052 32680 9064
rect 32732 9092 32738 9104
rect 34440 9092 34468 9132
rect 35710 9120 35716 9132
rect 35768 9120 35774 9172
rect 36354 9120 36360 9172
rect 36412 9120 36418 9172
rect 32732 9064 34468 9092
rect 32732 9052 32738 9064
rect 25038 8984 25044 9036
rect 25096 8984 25102 9036
rect 25774 8984 25780 9036
rect 25832 9024 25838 9036
rect 25832 8996 26280 9024
rect 25832 8984 25838 8996
rect 21542 8916 21548 8968
rect 21600 8956 21606 8968
rect 22649 8959 22707 8965
rect 22649 8956 22661 8959
rect 21600 8928 22661 8956
rect 21600 8916 21606 8928
rect 22649 8925 22661 8928
rect 22695 8925 22707 8959
rect 22649 8919 22707 8925
rect 24578 8916 24584 8968
rect 24636 8956 24642 8968
rect 24765 8959 24823 8965
rect 24765 8956 24777 8959
rect 24636 8928 24777 8956
rect 24636 8916 24642 8928
rect 24765 8925 24777 8928
rect 24811 8925 24823 8959
rect 26252 8956 26280 8996
rect 26602 8984 26608 9036
rect 26660 9024 26666 9036
rect 27338 9024 27344 9036
rect 26660 8996 27344 9024
rect 26660 8984 26666 8996
rect 27338 8984 27344 8996
rect 27396 9024 27402 9036
rect 27801 9027 27859 9033
rect 27801 9024 27813 9027
rect 27396 8996 27813 9024
rect 27396 8984 27402 8996
rect 27801 8993 27813 8996
rect 27847 8993 27859 9027
rect 30469 9027 30527 9033
rect 27801 8987 27859 8993
rect 27908 8996 29132 9024
rect 27908 8956 27936 8996
rect 26252 8928 27936 8956
rect 24765 8919 24823 8925
rect 28994 8916 29000 8968
rect 29052 8916 29058 8968
rect 29104 8956 29132 8996
rect 30469 8993 30481 9027
rect 30515 9024 30527 9027
rect 30650 9024 30656 9036
rect 30515 8996 30656 9024
rect 30515 8993 30527 8996
rect 30469 8987 30527 8993
rect 30650 8984 30656 8996
rect 30708 8984 30714 9036
rect 34514 9024 34520 9036
rect 30760 8996 31156 9024
rect 30760 8956 30788 8996
rect 29104 8928 30788 8956
rect 31021 8959 31079 8965
rect 31021 8925 31033 8959
rect 31067 8925 31079 8959
rect 31021 8919 31079 8925
rect 21082 8848 21088 8900
rect 21140 8888 21146 8900
rect 21729 8891 21787 8897
rect 21729 8888 21741 8891
rect 21140 8860 21741 8888
rect 21140 8848 21146 8860
rect 21729 8857 21741 8860
rect 21775 8857 21787 8891
rect 21729 8851 21787 8857
rect 22738 8848 22744 8900
rect 22796 8888 22802 8900
rect 22894 8891 22952 8897
rect 22894 8888 22906 8891
rect 22796 8860 22906 8888
rect 22796 8848 22802 8860
rect 22894 8857 22906 8860
rect 22940 8857 22952 8891
rect 22894 8851 22952 8857
rect 25682 8848 25688 8900
rect 25740 8848 25746 8900
rect 27706 8848 27712 8900
rect 27764 8848 27770 8900
rect 28902 8848 28908 8900
rect 28960 8888 28966 8900
rect 31036 8888 31064 8919
rect 28960 8860 31064 8888
rect 28960 8848 28966 8860
rect 19935 8792 20852 8820
rect 22189 8823 22247 8829
rect 19935 8789 19947 8792
rect 19889 8783 19947 8789
rect 22189 8789 22201 8823
rect 22235 8820 22247 8823
rect 22646 8820 22652 8832
rect 22235 8792 22652 8820
rect 22235 8789 22247 8792
rect 22189 8783 22247 8789
rect 22646 8780 22652 8792
rect 22704 8780 22710 8832
rect 24026 8780 24032 8832
rect 24084 8780 24090 8832
rect 25958 8780 25964 8832
rect 26016 8820 26022 8832
rect 26513 8823 26571 8829
rect 26513 8820 26525 8823
rect 26016 8792 26525 8820
rect 26016 8780 26022 8792
rect 26513 8789 26525 8792
rect 26559 8789 26571 8823
rect 26513 8783 26571 8789
rect 27614 8780 27620 8832
rect 27672 8780 27678 8832
rect 30190 8780 30196 8832
rect 30248 8780 30254 8832
rect 30282 8780 30288 8832
rect 30340 8780 30346 8832
rect 31128 8820 31156 8996
rect 32876 8996 34520 9024
rect 31570 8916 31576 8968
rect 31628 8956 31634 8968
rect 32876 8956 32904 8996
rect 34514 8984 34520 8996
rect 34572 8984 34578 9036
rect 31628 8928 32904 8956
rect 31628 8916 31634 8928
rect 32950 8916 32956 8968
rect 33008 8916 33014 8968
rect 34330 8916 34336 8968
rect 34388 8916 34394 8968
rect 34606 8916 34612 8968
rect 34664 8956 34670 8968
rect 34977 8959 35035 8965
rect 34977 8956 34989 8959
rect 34664 8928 34989 8956
rect 34664 8916 34670 8928
rect 34977 8925 34989 8928
rect 35023 8956 35035 8959
rect 37458 8956 37464 8968
rect 35023 8928 37464 8956
rect 35023 8925 35035 8928
rect 34977 8919 35035 8925
rect 37458 8916 37464 8928
rect 37516 8916 37522 8968
rect 37550 8916 37556 8968
rect 37608 8956 37614 8968
rect 37717 8959 37775 8965
rect 37717 8956 37729 8959
rect 37608 8928 37729 8956
rect 37608 8916 37614 8928
rect 37717 8925 37729 8928
rect 37763 8925 37775 8959
rect 37717 8919 37775 8925
rect 44358 8916 44364 8968
rect 44416 8916 44422 8968
rect 31288 8891 31346 8897
rect 31288 8857 31300 8891
rect 31334 8888 31346 8891
rect 31478 8888 31484 8900
rect 31334 8860 31484 8888
rect 31334 8857 31346 8860
rect 31288 8851 31346 8857
rect 31478 8848 31484 8860
rect 31536 8848 31542 8900
rect 34146 8848 34152 8900
rect 34204 8888 34210 8900
rect 35222 8891 35280 8897
rect 35222 8888 35234 8891
rect 34204 8860 35234 8888
rect 34204 8848 34210 8860
rect 35222 8857 35234 8860
rect 35268 8857 35280 8891
rect 38930 8888 38936 8900
rect 35222 8851 35280 8857
rect 37844 8860 38936 8888
rect 31938 8820 31944 8832
rect 31128 8792 31944 8820
rect 31938 8780 31944 8792
rect 31996 8820 32002 8832
rect 34974 8820 34980 8832
rect 31996 8792 34980 8820
rect 31996 8780 32002 8792
rect 34974 8780 34980 8792
rect 35032 8820 35038 8832
rect 37844 8820 37872 8860
rect 38930 8848 38936 8860
rect 38988 8848 38994 8900
rect 35032 8792 37872 8820
rect 35032 8780 35038 8792
rect 37918 8780 37924 8832
rect 37976 8820 37982 8832
rect 38841 8823 38899 8829
rect 38841 8820 38853 8823
rect 37976 8792 38853 8820
rect 37976 8780 37982 8792
rect 38841 8789 38853 8792
rect 38887 8789 38899 8823
rect 38841 8783 38899 8789
rect 44174 8780 44180 8832
rect 44232 8780 44238 8832
rect 1104 8730 45051 8752
rect 1104 8678 11896 8730
rect 11948 8678 11960 8730
rect 12012 8678 12024 8730
rect 12076 8678 12088 8730
rect 12140 8678 12152 8730
rect 12204 8678 22843 8730
rect 22895 8678 22907 8730
rect 22959 8678 22971 8730
rect 23023 8678 23035 8730
rect 23087 8678 23099 8730
rect 23151 8678 33790 8730
rect 33842 8678 33854 8730
rect 33906 8678 33918 8730
rect 33970 8678 33982 8730
rect 34034 8678 34046 8730
rect 34098 8678 44737 8730
rect 44789 8678 44801 8730
rect 44853 8678 44865 8730
rect 44917 8678 44929 8730
rect 44981 8678 44993 8730
rect 45045 8678 45051 8730
rect 1104 8656 45051 8678
rect 2038 8576 2044 8628
rect 2096 8616 2102 8628
rect 2096 8588 3556 8616
rect 2096 8576 2102 8588
rect 3528 8548 3556 8588
rect 4338 8576 4344 8628
rect 4396 8616 4402 8628
rect 5353 8619 5411 8625
rect 5353 8616 5365 8619
rect 4396 8588 5365 8616
rect 4396 8576 4402 8588
rect 5353 8585 5365 8588
rect 5399 8585 5411 8619
rect 5353 8579 5411 8585
rect 4218 8551 4276 8557
rect 4218 8548 4230 8551
rect 2148 8520 2774 8548
rect 3528 8520 4230 8548
rect 2148 8489 2176 8520
rect 2133 8483 2191 8489
rect 2133 8449 2145 8483
rect 2179 8449 2191 8483
rect 2133 8443 2191 8449
rect 2222 8440 2228 8492
rect 2280 8480 2286 8492
rect 2389 8483 2447 8489
rect 2389 8480 2401 8483
rect 2280 8452 2401 8480
rect 2280 8440 2286 8452
rect 2389 8449 2401 8452
rect 2435 8449 2447 8483
rect 2746 8480 2774 8520
rect 4218 8517 4230 8520
rect 4264 8517 4276 8551
rect 5368 8548 5396 8579
rect 8202 8576 8208 8628
rect 8260 8576 8266 8628
rect 9674 8616 9680 8628
rect 8312 8588 9680 8616
rect 8312 8548 8340 8588
rect 9674 8576 9680 8588
rect 9732 8576 9738 8628
rect 10042 8576 10048 8628
rect 10100 8576 10106 8628
rect 15654 8576 15660 8628
rect 15712 8616 15718 8628
rect 15712 8588 24808 8616
rect 15712 8576 15718 8588
rect 8938 8557 8944 8560
rect 8932 8548 8944 8557
rect 5368 8520 8340 8548
rect 8899 8520 8944 8548
rect 4218 8511 4276 8517
rect 8932 8511 8944 8520
rect 8938 8508 8944 8511
rect 8996 8508 9002 8560
rect 17126 8548 17132 8560
rect 16868 8520 17132 8548
rect 3970 8480 3976 8492
rect 2746 8452 3976 8480
rect 2389 8443 2447 8449
rect 3970 8440 3976 8452
rect 4028 8440 4034 8492
rect 7101 8483 7159 8489
rect 7101 8449 7113 8483
rect 7147 8480 7159 8483
rect 9490 8480 9496 8492
rect 7147 8452 9496 8480
rect 7147 8449 7159 8452
rect 7101 8443 7159 8449
rect 9490 8440 9496 8452
rect 9548 8440 9554 8492
rect 14185 8483 14243 8489
rect 14185 8449 14197 8483
rect 14231 8449 14243 8483
rect 14185 8443 14243 8449
rect 7653 8415 7711 8421
rect 7653 8381 7665 8415
rect 7699 8412 7711 8415
rect 8294 8412 8300 8424
rect 7699 8384 8300 8412
rect 7699 8381 7711 8384
rect 7653 8375 7711 8381
rect 8294 8372 8300 8384
rect 8352 8372 8358 8424
rect 8662 8372 8668 8424
rect 8720 8372 8726 8424
rect 14200 8412 14228 8443
rect 14366 8440 14372 8492
rect 14424 8440 14430 8492
rect 16114 8440 16120 8492
rect 16172 8440 16178 8492
rect 16868 8489 16896 8520
rect 17126 8508 17132 8520
rect 17184 8508 17190 8560
rect 17218 8508 17224 8560
rect 17276 8548 17282 8560
rect 19981 8551 20039 8557
rect 17276 8520 17618 8548
rect 17276 8508 17282 8520
rect 19981 8517 19993 8551
rect 20027 8548 20039 8551
rect 20254 8548 20260 8560
rect 20027 8520 20260 8548
rect 20027 8517 20039 8520
rect 19981 8511 20039 8517
rect 20254 8508 20260 8520
rect 20312 8548 20318 8560
rect 20809 8551 20867 8557
rect 20809 8548 20821 8551
rect 20312 8520 20821 8548
rect 20312 8508 20318 8520
rect 20809 8517 20821 8520
rect 20855 8517 20867 8551
rect 20809 8511 20867 8517
rect 21082 8508 21088 8560
rect 21140 8548 21146 8560
rect 22189 8551 22247 8557
rect 22189 8548 22201 8551
rect 21140 8520 22201 8548
rect 21140 8508 21146 8520
rect 22189 8517 22201 8520
rect 22235 8548 22247 8551
rect 24026 8548 24032 8560
rect 22235 8520 24032 8548
rect 22235 8517 22247 8520
rect 22189 8511 22247 8517
rect 24026 8508 24032 8520
rect 24084 8508 24090 8560
rect 24780 8557 24808 8588
rect 25590 8576 25596 8628
rect 25648 8576 25654 8628
rect 25958 8576 25964 8628
rect 26016 8576 26022 8628
rect 30190 8576 30196 8628
rect 30248 8616 30254 8628
rect 31021 8619 31079 8625
rect 31021 8616 31033 8619
rect 30248 8588 31033 8616
rect 30248 8576 30254 8588
rect 31021 8585 31033 8588
rect 31067 8585 31079 8619
rect 31021 8579 31079 8585
rect 31478 8576 31484 8628
rect 31536 8576 31542 8628
rect 33965 8619 34023 8625
rect 33965 8585 33977 8619
rect 34011 8585 34023 8619
rect 33965 8579 34023 8585
rect 24765 8551 24823 8557
rect 24765 8517 24777 8551
rect 24811 8548 24823 8551
rect 28718 8548 28724 8560
rect 24811 8520 28724 8548
rect 24811 8517 24823 8520
rect 24765 8511 24823 8517
rect 28718 8508 28724 8520
rect 28776 8508 28782 8560
rect 32490 8548 32496 8560
rect 28828 8520 32496 8548
rect 16853 8483 16911 8489
rect 16853 8449 16865 8483
rect 16899 8449 16911 8483
rect 16853 8443 16911 8449
rect 19058 8440 19064 8492
rect 19116 8440 19122 8492
rect 19153 8483 19211 8489
rect 19153 8449 19165 8483
rect 19199 8480 19211 8483
rect 19705 8483 19763 8489
rect 19705 8480 19717 8483
rect 19199 8452 19717 8480
rect 19199 8449 19211 8452
rect 19153 8443 19211 8449
rect 19705 8449 19717 8452
rect 19751 8480 19763 8483
rect 19794 8480 19800 8492
rect 19751 8452 19800 8480
rect 19751 8449 19763 8452
rect 19705 8443 19763 8449
rect 19794 8440 19800 8452
rect 19852 8440 19858 8492
rect 19886 8440 19892 8492
rect 19944 8440 19950 8492
rect 20073 8483 20131 8489
rect 20073 8449 20085 8483
rect 20119 8480 20131 8483
rect 20346 8480 20352 8492
rect 20119 8452 20352 8480
rect 20119 8449 20131 8452
rect 20073 8443 20131 8449
rect 20346 8440 20352 8452
rect 20404 8440 20410 8492
rect 20714 8440 20720 8492
rect 20772 8440 20778 8492
rect 22002 8440 22008 8492
rect 22060 8440 22066 8492
rect 23109 8483 23167 8489
rect 23109 8449 23121 8483
rect 23155 8480 23167 8483
rect 23382 8480 23388 8492
rect 23155 8452 23388 8480
rect 23155 8449 23167 8452
rect 23109 8443 23167 8449
rect 23382 8440 23388 8452
rect 23440 8440 23446 8492
rect 26053 8483 26111 8489
rect 26053 8449 26065 8483
rect 26099 8480 26111 8483
rect 27614 8480 27620 8492
rect 26099 8452 27620 8480
rect 26099 8449 26111 8452
rect 26053 8443 26111 8449
rect 27614 8440 27620 8452
rect 27672 8480 27678 8492
rect 28068 8483 28126 8489
rect 28068 8480 28080 8483
rect 27672 8452 28080 8480
rect 27672 8440 27678 8452
rect 28068 8449 28080 8452
rect 28114 8480 28126 8483
rect 28828 8480 28856 8520
rect 32490 8508 32496 8520
rect 32548 8508 32554 8560
rect 33980 8548 34008 8579
rect 34514 8576 34520 8628
rect 34572 8616 34578 8628
rect 37461 8619 37519 8625
rect 34572 8588 37412 8616
rect 34572 8576 34578 8588
rect 34854 8551 34912 8557
rect 34854 8548 34866 8551
rect 33980 8520 34866 8548
rect 34854 8517 34866 8520
rect 34900 8517 34912 8551
rect 37384 8548 37412 8588
rect 37461 8585 37473 8619
rect 37507 8616 37519 8619
rect 37734 8616 37740 8628
rect 37507 8588 37740 8616
rect 37507 8585 37519 8588
rect 37461 8579 37519 8585
rect 37734 8576 37740 8588
rect 37792 8576 37798 8628
rect 37826 8576 37832 8628
rect 37884 8616 37890 8628
rect 37921 8619 37979 8625
rect 37921 8616 37933 8619
rect 37884 8588 37933 8616
rect 37884 8576 37890 8588
rect 37921 8585 37933 8588
rect 37967 8585 37979 8619
rect 37921 8579 37979 8585
rect 37384 8520 40540 8548
rect 34854 8511 34912 8517
rect 28114 8452 28856 8480
rect 28114 8449 28126 8452
rect 28068 8443 28126 8449
rect 29730 8440 29736 8492
rect 29788 8480 29794 8492
rect 29897 8483 29955 8489
rect 29897 8480 29909 8483
rect 29788 8452 29909 8480
rect 29788 8440 29794 8452
rect 29897 8449 29909 8452
rect 29943 8449 29955 8483
rect 29897 8443 29955 8449
rect 30190 8440 30196 8492
rect 30248 8480 30254 8492
rect 31570 8480 31576 8492
rect 30248 8452 31576 8480
rect 30248 8440 30254 8452
rect 31570 8440 31576 8452
rect 31628 8440 31634 8492
rect 31662 8440 31668 8492
rect 31720 8440 31726 8492
rect 34149 8483 34207 8489
rect 34149 8449 34161 8483
rect 34195 8480 34207 8483
rect 34514 8480 34520 8492
rect 34195 8452 34520 8480
rect 34195 8449 34207 8452
rect 34149 8443 34207 8449
rect 34514 8440 34520 8452
rect 34572 8440 34578 8492
rect 34606 8440 34612 8492
rect 34664 8440 34670 8492
rect 37829 8483 37887 8489
rect 37829 8449 37841 8483
rect 37875 8480 37887 8483
rect 37918 8480 37924 8492
rect 37875 8452 37924 8480
rect 37875 8449 37887 8452
rect 37829 8443 37887 8449
rect 37918 8440 37924 8452
rect 37976 8440 37982 8492
rect 40512 8489 40540 8520
rect 40497 8483 40555 8489
rect 40497 8449 40509 8483
rect 40543 8480 40555 8483
rect 42610 8480 42616 8492
rect 40543 8452 42616 8480
rect 40543 8449 40555 8452
rect 40497 8443 40555 8449
rect 42610 8440 42616 8452
rect 42668 8440 42674 8492
rect 14918 8412 14924 8424
rect 14200 8384 14924 8412
rect 14918 8372 14924 8384
rect 14976 8372 14982 8424
rect 16206 8372 16212 8424
rect 16264 8412 16270 8424
rect 17129 8415 17187 8421
rect 17129 8412 17141 8415
rect 16264 8384 17141 8412
rect 16264 8372 16270 8384
rect 17129 8381 17141 8384
rect 17175 8381 17187 8415
rect 17129 8375 17187 8381
rect 26142 8372 26148 8424
rect 26200 8372 26206 8424
rect 27801 8415 27859 8421
rect 27801 8381 27813 8415
rect 27847 8381 27859 8415
rect 28902 8412 28908 8424
rect 27801 8375 27859 8381
rect 28828 8384 28908 8412
rect 3234 8304 3240 8356
rect 3292 8344 3298 8356
rect 3513 8347 3571 8353
rect 3513 8344 3525 8347
rect 3292 8316 3525 8344
rect 3292 8304 3298 8316
rect 3513 8313 3525 8316
rect 3559 8313 3571 8347
rect 3513 8307 3571 8313
rect 6914 8304 6920 8356
rect 6972 8304 6978 8356
rect 16224 8316 16988 8344
rect 14277 8279 14335 8285
rect 14277 8245 14289 8279
rect 14323 8276 14335 8279
rect 14642 8276 14648 8288
rect 14323 8248 14648 8276
rect 14323 8245 14335 8248
rect 14277 8239 14335 8245
rect 14642 8236 14648 8248
rect 14700 8236 14706 8288
rect 16224 8285 16252 8316
rect 16209 8279 16267 8285
rect 16209 8245 16221 8279
rect 16255 8245 16267 8279
rect 16960 8276 16988 8316
rect 18598 8304 18604 8356
rect 18656 8304 18662 8356
rect 17218 8276 17224 8288
rect 16960 8248 17224 8276
rect 16209 8239 16267 8245
rect 17218 8236 17224 8248
rect 17276 8236 17282 8288
rect 20070 8236 20076 8288
rect 20128 8276 20134 8288
rect 20257 8279 20315 8285
rect 20257 8276 20269 8279
rect 20128 8248 20269 8276
rect 20128 8236 20134 8248
rect 20257 8245 20269 8248
rect 20303 8245 20315 8279
rect 20257 8239 20315 8245
rect 22186 8236 22192 8288
rect 22244 8276 22250 8288
rect 22373 8279 22431 8285
rect 22373 8276 22385 8279
rect 22244 8248 22385 8276
rect 22244 8236 22250 8248
rect 22373 8245 22385 8248
rect 22419 8245 22431 8279
rect 27816 8276 27844 8375
rect 28166 8276 28172 8288
rect 27816 8248 28172 8276
rect 22373 8239 22431 8245
rect 28166 8236 28172 8248
rect 28224 8276 28230 8288
rect 28828 8276 28856 8384
rect 28902 8372 28908 8384
rect 28960 8412 28966 8424
rect 29641 8415 29699 8421
rect 29641 8412 29653 8415
rect 28960 8384 29653 8412
rect 28960 8372 28966 8384
rect 29641 8381 29653 8384
rect 29687 8381 29699 8415
rect 29641 8375 29699 8381
rect 35710 8372 35716 8424
rect 35768 8412 35774 8424
rect 38013 8415 38071 8421
rect 38013 8412 38025 8415
rect 35768 8384 38025 8412
rect 35768 8372 35774 8384
rect 38013 8381 38025 8384
rect 38059 8381 38071 8415
rect 38013 8375 38071 8381
rect 35618 8304 35624 8356
rect 35676 8344 35682 8356
rect 35989 8347 36047 8353
rect 35989 8344 36001 8347
rect 35676 8316 36001 8344
rect 35676 8304 35682 8316
rect 35989 8313 36001 8316
rect 36035 8313 36047 8347
rect 35989 8307 36047 8313
rect 40589 8347 40647 8353
rect 40589 8313 40601 8347
rect 40635 8344 40647 8347
rect 41414 8344 41420 8356
rect 40635 8316 41420 8344
rect 40635 8313 40647 8316
rect 40589 8307 40647 8313
rect 41414 8304 41420 8316
rect 41472 8304 41478 8356
rect 28224 8248 28856 8276
rect 28224 8236 28230 8248
rect 29178 8236 29184 8288
rect 29236 8236 29242 8288
rect 1104 8186 44896 8208
rect 1104 8134 6423 8186
rect 6475 8134 6487 8186
rect 6539 8134 6551 8186
rect 6603 8134 6615 8186
rect 6667 8134 6679 8186
rect 6731 8134 17370 8186
rect 17422 8134 17434 8186
rect 17486 8134 17498 8186
rect 17550 8134 17562 8186
rect 17614 8134 17626 8186
rect 17678 8134 28317 8186
rect 28369 8134 28381 8186
rect 28433 8134 28445 8186
rect 28497 8134 28509 8186
rect 28561 8134 28573 8186
rect 28625 8134 39264 8186
rect 39316 8134 39328 8186
rect 39380 8134 39392 8186
rect 39444 8134 39456 8186
rect 39508 8134 39520 8186
rect 39572 8134 44896 8186
rect 1104 8112 44896 8134
rect 5350 8032 5356 8084
rect 5408 8032 5414 8084
rect 6270 8032 6276 8084
rect 6328 8072 6334 8084
rect 6457 8075 6515 8081
rect 6457 8072 6469 8075
rect 6328 8044 6469 8072
rect 6328 8032 6334 8044
rect 6457 8041 6469 8044
rect 6503 8041 6515 8075
rect 6457 8035 6515 8041
rect 8389 8075 8447 8081
rect 8389 8041 8401 8075
rect 8435 8072 8447 8075
rect 8570 8072 8576 8084
rect 8435 8044 8576 8072
rect 8435 8041 8447 8044
rect 8389 8035 8447 8041
rect 8570 8032 8576 8044
rect 8628 8032 8634 8084
rect 11790 8032 11796 8084
rect 11848 8072 11854 8084
rect 12437 8075 12495 8081
rect 12437 8072 12449 8075
rect 11848 8044 12449 8072
rect 11848 8032 11854 8044
rect 12437 8041 12449 8044
rect 12483 8041 12495 8075
rect 12437 8035 12495 8041
rect 14918 8032 14924 8084
rect 14976 8072 14982 8084
rect 25041 8075 25099 8081
rect 25041 8072 25053 8075
rect 14976 8044 18460 8072
rect 14976 8032 14982 8044
rect 3326 7896 3332 7948
rect 3384 7936 3390 7948
rect 3878 7936 3884 7948
rect 3384 7908 3884 7936
rect 3384 7896 3390 7908
rect 3878 7896 3884 7908
rect 3936 7936 3942 7948
rect 3973 7939 4031 7945
rect 3973 7936 3985 7939
rect 3936 7908 3985 7936
rect 3936 7896 3942 7908
rect 3973 7905 3985 7908
rect 4019 7905 4031 7939
rect 3973 7899 4031 7905
rect 5902 7896 5908 7948
rect 5960 7896 5966 7948
rect 9122 7896 9128 7948
rect 9180 7896 9186 7948
rect 14090 7936 14096 7948
rect 12084 7908 14096 7936
rect 2041 7871 2099 7877
rect 2041 7837 2053 7871
rect 2087 7868 2099 7871
rect 3344 7868 3372 7896
rect 4240 7871 4298 7877
rect 4240 7868 4252 7871
rect 2087 7840 3372 7868
rect 4172 7840 4252 7868
rect 2087 7837 2099 7840
rect 2041 7831 2099 7837
rect 2314 7809 2320 7812
rect 2308 7763 2320 7809
rect 2314 7760 2320 7763
rect 2372 7760 2378 7812
rect 3421 7735 3479 7741
rect 3421 7701 3433 7735
rect 3467 7732 3479 7735
rect 4172 7732 4200 7840
rect 4240 7837 4252 7840
rect 4286 7868 4298 7871
rect 6917 7871 6975 7877
rect 6917 7868 6929 7871
rect 4286 7840 6929 7868
rect 4286 7837 4298 7840
rect 4240 7831 4298 7837
rect 6917 7837 6929 7840
rect 6963 7837 6975 7871
rect 6917 7831 6975 7837
rect 8018 7828 8024 7880
rect 8076 7828 8082 7880
rect 8205 7871 8263 7877
rect 8205 7837 8217 7871
rect 8251 7868 8263 7871
rect 8570 7868 8576 7880
rect 8251 7840 8576 7868
rect 8251 7837 8263 7840
rect 8205 7831 8263 7837
rect 8570 7828 8576 7840
rect 8628 7828 8634 7880
rect 10502 7828 10508 7880
rect 10560 7868 10566 7880
rect 12084 7877 12112 7908
rect 14090 7896 14096 7908
rect 14148 7896 14154 7948
rect 18138 7936 18144 7948
rect 16040 7908 18144 7936
rect 10965 7871 11023 7877
rect 10965 7868 10977 7871
rect 10560 7840 10977 7868
rect 10560 7828 10566 7840
rect 10965 7837 10977 7840
rect 11011 7837 11023 7871
rect 12069 7871 12127 7877
rect 12069 7868 12081 7871
rect 10965 7831 11023 7837
rect 11072 7840 12081 7868
rect 4430 7760 4436 7812
rect 4488 7800 4494 7812
rect 7926 7800 7932 7812
rect 4488 7772 7932 7800
rect 4488 7760 4494 7772
rect 7926 7760 7932 7772
rect 7984 7760 7990 7812
rect 8294 7760 8300 7812
rect 8352 7800 8358 7812
rect 9370 7803 9428 7809
rect 9370 7800 9382 7803
rect 8352 7772 9382 7800
rect 8352 7760 8358 7772
rect 9370 7769 9382 7772
rect 9416 7769 9428 7803
rect 9370 7763 9428 7769
rect 9766 7760 9772 7812
rect 9824 7800 9830 7812
rect 11072 7800 11100 7840
rect 12069 7837 12081 7840
rect 12115 7837 12127 7871
rect 12069 7831 12127 7837
rect 12253 7871 12311 7877
rect 12253 7837 12265 7871
rect 12299 7837 12311 7871
rect 12253 7831 12311 7837
rect 13265 7871 13323 7877
rect 13265 7837 13277 7871
rect 13311 7837 13323 7871
rect 13265 7831 13323 7837
rect 9824 7772 11100 7800
rect 9824 7760 9830 7772
rect 11146 7760 11152 7812
rect 11204 7800 11210 7812
rect 12268 7800 12296 7831
rect 11204 7772 12296 7800
rect 13280 7800 13308 7831
rect 13354 7828 13360 7880
rect 13412 7828 13418 7880
rect 14458 7828 14464 7880
rect 14516 7868 14522 7880
rect 14553 7871 14611 7877
rect 14553 7868 14565 7871
rect 14516 7840 14565 7868
rect 14516 7828 14522 7840
rect 14553 7837 14565 7840
rect 14599 7837 14611 7871
rect 14553 7831 14611 7837
rect 15286 7828 15292 7880
rect 15344 7868 15350 7880
rect 16040 7877 16068 7908
rect 18138 7896 18144 7908
rect 18196 7896 18202 7948
rect 18432 7936 18460 8044
rect 19720 8044 25053 8072
rect 18432 7908 18644 7936
rect 15381 7871 15439 7877
rect 15381 7868 15393 7871
rect 15344 7840 15393 7868
rect 15344 7828 15350 7840
rect 15381 7837 15393 7840
rect 15427 7837 15439 7871
rect 15381 7831 15439 7837
rect 16025 7871 16083 7877
rect 16025 7837 16037 7871
rect 16071 7837 16083 7871
rect 16025 7831 16083 7837
rect 16114 7828 16120 7880
rect 16172 7868 16178 7880
rect 16485 7871 16543 7877
rect 16485 7868 16497 7871
rect 16172 7840 16497 7868
rect 16172 7828 16178 7840
rect 16485 7837 16497 7840
rect 16531 7837 16543 7871
rect 16485 7831 16543 7837
rect 17126 7828 17132 7880
rect 17184 7828 17190 7880
rect 18616 7868 18644 7908
rect 19720 7877 19748 8044
rect 25041 8041 25053 8044
rect 25087 8041 25099 8075
rect 25041 8035 25099 8041
rect 25682 8032 25688 8084
rect 25740 8032 25746 8084
rect 29730 8032 29736 8084
rect 29788 8032 29794 8084
rect 34514 8032 34520 8084
rect 34572 8072 34578 8084
rect 34885 8075 34943 8081
rect 34885 8072 34897 8075
rect 34572 8044 34897 8072
rect 34572 8032 34578 8044
rect 34885 8041 34897 8044
rect 34931 8041 34943 8075
rect 40494 8072 40500 8084
rect 34885 8035 34943 8041
rect 39500 8044 40500 8072
rect 23934 7964 23940 8016
rect 23992 8004 23998 8016
rect 28994 8004 29000 8016
rect 23992 7976 29000 8004
rect 23992 7964 23998 7976
rect 28994 7964 29000 7976
rect 29052 8004 29058 8016
rect 30190 8004 30196 8016
rect 29052 7976 30196 8004
rect 29052 7964 29058 7976
rect 30190 7964 30196 7976
rect 30248 7964 30254 8016
rect 19794 7896 19800 7948
rect 19852 7936 19858 7948
rect 19981 7939 20039 7945
rect 19981 7936 19993 7939
rect 19852 7908 19993 7936
rect 19852 7896 19858 7908
rect 19981 7905 19993 7908
rect 20027 7905 20039 7939
rect 19981 7899 20039 7905
rect 20073 7939 20131 7945
rect 20073 7905 20085 7939
rect 20119 7936 20131 7939
rect 20346 7936 20352 7948
rect 20119 7908 20352 7936
rect 20119 7905 20131 7908
rect 20073 7899 20131 7905
rect 20346 7896 20352 7908
rect 20404 7936 20410 7948
rect 20404 7908 20944 7936
rect 20404 7896 20410 7908
rect 19705 7871 19763 7877
rect 18616 7840 18736 7868
rect 13722 7800 13728 7812
rect 13280 7772 13728 7800
rect 11204 7760 11210 7772
rect 13722 7760 13728 7772
rect 13780 7800 13786 7812
rect 15010 7800 15016 7812
rect 13780 7772 15016 7800
rect 13780 7760 13786 7772
rect 15010 7760 15016 7772
rect 15068 7760 15074 7812
rect 17405 7803 17463 7809
rect 17405 7800 17417 7803
rect 15856 7772 17417 7800
rect 3467 7704 4200 7732
rect 3467 7701 3479 7704
rect 3421 7695 3479 7701
rect 5626 7692 5632 7744
rect 5684 7732 5690 7744
rect 7561 7735 7619 7741
rect 7561 7732 7573 7735
rect 5684 7704 7573 7732
rect 5684 7692 5690 7704
rect 7561 7701 7573 7704
rect 7607 7701 7619 7735
rect 7561 7695 7619 7701
rect 10502 7692 10508 7744
rect 10560 7692 10566 7744
rect 11606 7692 11612 7744
rect 11664 7692 11670 7744
rect 12986 7692 12992 7744
rect 13044 7732 13050 7744
rect 13541 7735 13599 7741
rect 13541 7732 13553 7735
rect 13044 7704 13553 7732
rect 13044 7692 13050 7704
rect 13541 7701 13553 7704
rect 13587 7701 13599 7735
rect 13541 7695 13599 7701
rect 14366 7692 14372 7744
rect 14424 7732 14430 7744
rect 14645 7735 14703 7741
rect 14645 7732 14657 7735
rect 14424 7704 14657 7732
rect 14424 7692 14430 7704
rect 14645 7701 14657 7704
rect 14691 7732 14703 7735
rect 15102 7732 15108 7744
rect 14691 7704 15108 7732
rect 14691 7701 14703 7704
rect 14645 7695 14703 7701
rect 15102 7692 15108 7704
rect 15160 7692 15166 7744
rect 15194 7692 15200 7744
rect 15252 7692 15258 7744
rect 15856 7741 15884 7772
rect 17405 7769 17417 7772
rect 17451 7769 17463 7803
rect 18708 7800 18736 7840
rect 19705 7837 19717 7871
rect 19751 7837 19763 7871
rect 19705 7831 19763 7837
rect 19886 7828 19892 7880
rect 19944 7828 19950 7880
rect 20254 7828 20260 7880
rect 20312 7828 20318 7880
rect 20916 7877 20944 7908
rect 21542 7896 21548 7948
rect 21600 7896 21606 7948
rect 24026 7896 24032 7948
rect 24084 7936 24090 7948
rect 24673 7939 24731 7945
rect 24673 7936 24685 7939
rect 24084 7908 24685 7936
rect 24084 7896 24090 7908
rect 24673 7905 24685 7908
rect 24719 7905 24731 7939
rect 25958 7936 25964 7948
rect 24673 7899 24731 7905
rect 24780 7908 25964 7936
rect 20901 7871 20959 7877
rect 20901 7837 20913 7871
rect 20947 7837 20959 7871
rect 20901 7831 20959 7837
rect 20916 7800 20944 7831
rect 21082 7828 21088 7880
rect 21140 7828 21146 7880
rect 22370 7828 22376 7880
rect 22428 7868 22434 7880
rect 24780 7877 24808 7908
rect 25958 7896 25964 7908
rect 26016 7896 26022 7948
rect 27614 7896 27620 7948
rect 27672 7936 27678 7948
rect 28721 7939 28779 7945
rect 28721 7936 28733 7939
rect 27672 7908 28733 7936
rect 27672 7896 27678 7908
rect 28721 7905 28733 7908
rect 28767 7905 28779 7939
rect 28721 7899 28779 7905
rect 31389 7939 31447 7945
rect 31389 7905 31401 7939
rect 31435 7936 31447 7939
rect 32950 7936 32956 7948
rect 31435 7908 32956 7936
rect 31435 7905 31447 7908
rect 31389 7899 31447 7905
rect 32950 7896 32956 7908
rect 33008 7896 33014 7948
rect 34698 7896 34704 7948
rect 34756 7936 34762 7948
rect 35345 7939 35403 7945
rect 35345 7936 35357 7939
rect 34756 7908 35357 7936
rect 34756 7896 34762 7908
rect 35345 7905 35357 7908
rect 35391 7905 35403 7939
rect 35345 7899 35403 7905
rect 35529 7939 35587 7945
rect 35529 7905 35541 7939
rect 35575 7936 35587 7939
rect 35710 7936 35716 7948
rect 35575 7908 35716 7936
rect 35575 7905 35587 7908
rect 35529 7899 35587 7905
rect 35710 7896 35716 7908
rect 35768 7896 35774 7948
rect 37918 7896 37924 7948
rect 37976 7936 37982 7948
rect 39500 7945 39528 8044
rect 40494 8032 40500 8044
rect 40552 8032 40558 8084
rect 38197 7939 38255 7945
rect 38197 7936 38209 7939
rect 37976 7908 38209 7936
rect 37976 7896 37982 7908
rect 38197 7905 38209 7908
rect 38243 7905 38255 7939
rect 38197 7899 38255 7905
rect 39485 7939 39543 7945
rect 39485 7905 39497 7939
rect 39531 7905 39543 7939
rect 42245 7939 42303 7945
rect 42245 7936 42257 7939
rect 39485 7899 39543 7905
rect 40052 7908 42257 7936
rect 40052 7880 40080 7908
rect 42245 7905 42257 7908
rect 42291 7905 42303 7939
rect 42245 7899 42303 7905
rect 23569 7871 23627 7877
rect 23569 7868 23581 7871
rect 22428 7840 23581 7868
rect 22428 7828 22434 7840
rect 23569 7837 23581 7840
rect 23615 7837 23627 7871
rect 23569 7831 23627 7837
rect 24765 7871 24823 7877
rect 24765 7837 24777 7871
rect 24811 7837 24823 7871
rect 24765 7831 24823 7837
rect 25498 7828 25504 7880
rect 25556 7868 25562 7880
rect 25593 7871 25651 7877
rect 25593 7868 25605 7871
rect 25556 7840 25605 7868
rect 25556 7828 25562 7840
rect 25593 7837 25605 7840
rect 25639 7837 25651 7871
rect 25593 7831 25651 7837
rect 28905 7871 28963 7877
rect 28905 7837 28917 7871
rect 28951 7868 28963 7871
rect 29178 7868 29184 7880
rect 28951 7840 29184 7868
rect 28951 7837 28963 7840
rect 28905 7831 28963 7837
rect 29178 7828 29184 7840
rect 29236 7828 29242 7880
rect 29917 7871 29975 7877
rect 29917 7837 29929 7871
rect 29963 7837 29975 7871
rect 29917 7831 29975 7837
rect 21812 7803 21870 7809
rect 17405 7763 17463 7769
rect 17512 7772 17894 7800
rect 18708 7772 20852 7800
rect 20916 7772 21128 7800
rect 15841 7735 15899 7741
rect 15841 7701 15853 7735
rect 15887 7701 15899 7735
rect 15841 7695 15899 7701
rect 16577 7735 16635 7741
rect 16577 7701 16589 7735
rect 16623 7732 16635 7735
rect 17512 7732 17540 7772
rect 16623 7704 17540 7732
rect 18877 7735 18935 7741
rect 16623 7701 16635 7704
rect 16577 7695 16635 7701
rect 18877 7701 18889 7735
rect 18923 7732 18935 7735
rect 19334 7732 19340 7744
rect 18923 7704 19340 7732
rect 18923 7701 18935 7704
rect 18877 7695 18935 7701
rect 19334 7692 19340 7704
rect 19392 7732 19398 7744
rect 19978 7732 19984 7744
rect 19392 7704 19984 7732
rect 19392 7692 19398 7704
rect 19978 7692 19984 7704
rect 20036 7692 20042 7744
rect 20441 7735 20499 7741
rect 20441 7701 20453 7735
rect 20487 7732 20499 7735
rect 20714 7732 20720 7744
rect 20487 7704 20720 7732
rect 20487 7701 20499 7704
rect 20441 7695 20499 7701
rect 20714 7692 20720 7704
rect 20772 7692 20778 7744
rect 20824 7732 20852 7772
rect 20990 7732 20996 7744
rect 20824 7704 20996 7732
rect 20990 7692 20996 7704
rect 21048 7692 21054 7744
rect 21100 7732 21128 7772
rect 21812 7769 21824 7803
rect 21858 7800 21870 7803
rect 29089 7803 29147 7809
rect 21858 7772 23428 7800
rect 21858 7769 21870 7772
rect 21812 7763 21870 7769
rect 22002 7732 22008 7744
rect 21100 7704 22008 7732
rect 22002 7692 22008 7704
rect 22060 7732 22066 7744
rect 23400 7741 23428 7772
rect 29089 7769 29101 7803
rect 29135 7800 29147 7803
rect 29932 7800 29960 7831
rect 31018 7828 31024 7880
rect 31076 7868 31082 7880
rect 31113 7871 31171 7877
rect 31113 7868 31125 7871
rect 31076 7840 31125 7868
rect 31076 7828 31082 7840
rect 31113 7837 31125 7840
rect 31159 7837 31171 7871
rect 31113 7831 31171 7837
rect 32582 7828 32588 7880
rect 32640 7828 32646 7880
rect 35253 7871 35311 7877
rect 35253 7837 35265 7871
rect 35299 7868 35311 7871
rect 35618 7868 35624 7880
rect 35299 7840 35624 7868
rect 35299 7837 35311 7840
rect 35253 7831 35311 7837
rect 35618 7828 35624 7840
rect 35676 7828 35682 7880
rect 38289 7871 38347 7877
rect 38289 7837 38301 7871
rect 38335 7868 38347 7871
rect 39114 7868 39120 7880
rect 38335 7840 39120 7868
rect 38335 7837 38347 7840
rect 38289 7831 38347 7837
rect 39114 7828 39120 7840
rect 39172 7828 39178 7880
rect 39209 7871 39267 7877
rect 39209 7837 39221 7871
rect 39255 7837 39267 7871
rect 39209 7831 39267 7837
rect 29135 7772 29960 7800
rect 29135 7769 29147 7772
rect 29089 7763 29147 7769
rect 38930 7760 38936 7812
rect 38988 7800 38994 7812
rect 39224 7800 39252 7831
rect 39298 7828 39304 7880
rect 39356 7828 39362 7880
rect 40034 7828 40040 7880
rect 40092 7828 40098 7880
rect 41414 7828 41420 7880
rect 41472 7828 41478 7880
rect 39850 7800 39856 7812
rect 38988 7772 39856 7800
rect 38988 7760 38994 7772
rect 39850 7760 39856 7772
rect 39908 7760 39914 7812
rect 40310 7760 40316 7812
rect 40368 7760 40374 7812
rect 42518 7760 42524 7812
rect 42576 7760 42582 7812
rect 42978 7760 42984 7812
rect 43036 7760 43042 7812
rect 22925 7735 22983 7741
rect 22925 7732 22937 7735
rect 22060 7704 22937 7732
rect 22060 7692 22066 7704
rect 22925 7701 22937 7704
rect 22971 7701 22983 7735
rect 22925 7695 22983 7701
rect 23385 7735 23443 7741
rect 23385 7701 23397 7735
rect 23431 7701 23443 7735
rect 23385 7695 23443 7701
rect 32398 7692 32404 7744
rect 32456 7692 32462 7744
rect 35526 7692 35532 7744
rect 35584 7732 35590 7744
rect 38657 7735 38715 7741
rect 38657 7732 38669 7735
rect 35584 7704 38669 7732
rect 35584 7692 35590 7704
rect 38657 7701 38669 7704
rect 38703 7701 38715 7735
rect 38657 7695 38715 7701
rect 38746 7692 38752 7744
rect 38804 7732 38810 7744
rect 39485 7735 39543 7741
rect 39485 7732 39497 7735
rect 38804 7704 39497 7732
rect 38804 7692 38810 7704
rect 39485 7701 39497 7704
rect 39531 7701 39543 7735
rect 39485 7695 39543 7701
rect 40218 7692 40224 7744
rect 40276 7732 40282 7744
rect 40402 7732 40408 7744
rect 40276 7704 40408 7732
rect 40276 7692 40282 7704
rect 40402 7692 40408 7704
rect 40460 7732 40466 7744
rect 41785 7735 41843 7741
rect 41785 7732 41797 7735
rect 40460 7704 41797 7732
rect 40460 7692 40466 7704
rect 41785 7701 41797 7704
rect 41831 7701 41843 7735
rect 41785 7695 41843 7701
rect 43990 7692 43996 7744
rect 44048 7692 44054 7744
rect 1104 7642 45051 7664
rect 1104 7590 11896 7642
rect 11948 7590 11960 7642
rect 12012 7590 12024 7642
rect 12076 7590 12088 7642
rect 12140 7590 12152 7642
rect 12204 7590 22843 7642
rect 22895 7590 22907 7642
rect 22959 7590 22971 7642
rect 23023 7590 23035 7642
rect 23087 7590 23099 7642
rect 23151 7590 33790 7642
rect 33842 7590 33854 7642
rect 33906 7590 33918 7642
rect 33970 7590 33982 7642
rect 34034 7590 34046 7642
rect 34098 7590 44737 7642
rect 44789 7590 44801 7642
rect 44853 7590 44865 7642
rect 44917 7590 44929 7642
rect 44981 7590 44993 7642
rect 45045 7590 45051 7642
rect 1104 7568 45051 7590
rect 3878 7488 3884 7540
rect 3936 7488 3942 7540
rect 5626 7488 5632 7540
rect 5684 7488 5690 7540
rect 5718 7488 5724 7540
rect 5776 7528 5782 7540
rect 6917 7531 6975 7537
rect 6917 7528 6929 7531
rect 5776 7500 6929 7528
rect 5776 7488 5782 7500
rect 6917 7497 6929 7500
rect 6963 7497 6975 7531
rect 6917 7491 6975 7497
rect 9122 7488 9128 7540
rect 9180 7488 9186 7540
rect 9490 7488 9496 7540
rect 9548 7528 9554 7540
rect 10045 7531 10103 7537
rect 10045 7528 10057 7531
rect 9548 7500 10057 7528
rect 9548 7488 9554 7500
rect 10045 7497 10057 7500
rect 10091 7497 10103 7531
rect 10045 7491 10103 7497
rect 10505 7531 10563 7537
rect 10505 7497 10517 7531
rect 10551 7528 10563 7531
rect 11606 7528 11612 7540
rect 10551 7500 11612 7528
rect 10551 7497 10563 7500
rect 10505 7491 10563 7497
rect 11606 7488 11612 7500
rect 11664 7488 11670 7540
rect 14458 7488 14464 7540
rect 14516 7488 14522 7540
rect 16850 7488 16856 7540
rect 16908 7488 16914 7540
rect 17313 7531 17371 7537
rect 17313 7497 17325 7531
rect 17359 7528 17371 7531
rect 17862 7528 17868 7540
rect 17359 7500 17868 7528
rect 17359 7497 17371 7500
rect 17313 7491 17371 7497
rect 17862 7488 17868 7500
rect 17920 7488 17926 7540
rect 18138 7488 18144 7540
rect 18196 7488 18202 7540
rect 18509 7531 18567 7537
rect 18509 7497 18521 7531
rect 18555 7528 18567 7531
rect 19334 7528 19340 7540
rect 18555 7500 19340 7528
rect 18555 7497 18567 7500
rect 18509 7491 18567 7497
rect 19334 7488 19340 7500
rect 19392 7488 19398 7540
rect 20162 7488 20168 7540
rect 20220 7528 20226 7540
rect 20257 7531 20315 7537
rect 20257 7528 20269 7531
rect 20220 7500 20269 7528
rect 20220 7488 20226 7500
rect 20257 7497 20269 7500
rect 20303 7497 20315 7531
rect 20257 7491 20315 7497
rect 20990 7488 20996 7540
rect 21048 7528 21054 7540
rect 22205 7531 22263 7537
rect 22205 7528 22217 7531
rect 21048 7500 22217 7528
rect 21048 7488 21054 7500
rect 22205 7497 22217 7500
rect 22251 7497 22263 7531
rect 22205 7491 22263 7497
rect 22370 7488 22376 7540
rect 22428 7488 22434 7540
rect 22738 7488 22744 7540
rect 22796 7528 22802 7540
rect 22833 7531 22891 7537
rect 22833 7528 22845 7531
rect 22796 7500 22845 7528
rect 22796 7488 22802 7500
rect 22833 7497 22845 7500
rect 22879 7497 22891 7531
rect 22833 7491 22891 7497
rect 29917 7531 29975 7537
rect 29917 7497 29929 7531
rect 29963 7528 29975 7531
rect 30742 7528 30748 7540
rect 29963 7500 30748 7528
rect 29963 7497 29975 7500
rect 29917 7491 29975 7497
rect 30742 7488 30748 7500
rect 30800 7488 30806 7540
rect 39298 7528 39304 7540
rect 34348 7500 39304 7528
rect 2593 7463 2651 7469
rect 2593 7429 2605 7463
rect 2639 7460 2651 7463
rect 6822 7460 6828 7472
rect 2639 7432 6828 7460
rect 2639 7429 2651 7432
rect 2593 7423 2651 7429
rect 6822 7420 6828 7432
rect 6880 7460 6886 7472
rect 7837 7463 7895 7469
rect 7837 7460 7849 7463
rect 6880 7432 7849 7460
rect 6880 7420 6886 7432
rect 7837 7429 7849 7432
rect 7883 7429 7895 7463
rect 7837 7423 7895 7429
rect 7926 7420 7932 7472
rect 7984 7460 7990 7472
rect 13348 7463 13406 7469
rect 7984 7432 13308 7460
rect 7984 7420 7990 7432
rect 934 7352 940 7404
rect 992 7392 998 7404
rect 1765 7395 1823 7401
rect 1765 7392 1777 7395
rect 992 7364 1777 7392
rect 992 7352 998 7364
rect 1765 7361 1777 7364
rect 1811 7361 1823 7395
rect 1765 7355 1823 7361
rect 5534 7352 5540 7404
rect 5592 7352 5598 7404
rect 6733 7395 6791 7401
rect 6733 7392 6745 7395
rect 5644 7364 6745 7392
rect 5350 7284 5356 7336
rect 5408 7324 5414 7336
rect 5644 7324 5672 7364
rect 6733 7361 6745 7364
rect 6779 7361 6791 7395
rect 6733 7355 6791 7361
rect 9306 7352 9312 7404
rect 9364 7392 9370 7404
rect 10413 7395 10471 7401
rect 10413 7392 10425 7395
rect 9364 7364 10425 7392
rect 9364 7352 9370 7364
rect 10413 7361 10425 7364
rect 10459 7361 10471 7395
rect 10413 7355 10471 7361
rect 12618 7352 12624 7404
rect 12676 7352 12682 7404
rect 13280 7392 13308 7432
rect 13348 7429 13360 7463
rect 13394 7460 13406 7463
rect 15194 7460 15200 7472
rect 13394 7432 15200 7460
rect 13394 7429 13406 7432
rect 13348 7423 13406 7429
rect 15194 7420 15200 7432
rect 15252 7420 15258 7472
rect 17218 7420 17224 7472
rect 17276 7460 17282 7472
rect 18598 7460 18604 7472
rect 17276 7432 18604 7460
rect 17276 7420 17282 7432
rect 18598 7420 18604 7432
rect 18656 7420 18662 7472
rect 18800 7432 20852 7460
rect 13280 7364 14872 7392
rect 5408 7296 5672 7324
rect 5408 7284 5414 7296
rect 5810 7284 5816 7336
rect 5868 7284 5874 7336
rect 6549 7327 6607 7333
rect 6549 7293 6561 7327
rect 6595 7324 6607 7327
rect 8018 7324 8024 7336
rect 6595 7296 8024 7324
rect 6595 7293 6607 7296
rect 6549 7287 6607 7293
rect 8018 7284 8024 7296
rect 8076 7324 8082 7336
rect 9766 7324 9772 7336
rect 8076 7296 9772 7324
rect 8076 7284 8082 7296
rect 9766 7284 9772 7296
rect 9824 7284 9830 7336
rect 10594 7284 10600 7336
rect 10652 7284 10658 7336
rect 12250 7284 12256 7336
rect 12308 7324 12314 7336
rect 13081 7327 13139 7333
rect 13081 7324 13093 7327
rect 12308 7296 13093 7324
rect 12308 7284 12314 7296
rect 13081 7293 13093 7296
rect 13127 7293 13139 7327
rect 13081 7287 13139 7293
rect 1581 7259 1639 7265
rect 1581 7225 1593 7259
rect 1627 7256 1639 7259
rect 14844 7256 14872 7364
rect 14918 7352 14924 7404
rect 14976 7352 14982 7404
rect 15102 7352 15108 7404
rect 15160 7352 15166 7404
rect 18800 7392 18828 7432
rect 18616 7364 18828 7392
rect 17497 7327 17555 7333
rect 17497 7293 17509 7327
rect 17543 7324 17555 7327
rect 18322 7324 18328 7336
rect 17543 7296 18328 7324
rect 17543 7293 17555 7296
rect 17497 7287 17555 7293
rect 18322 7284 18328 7296
rect 18380 7284 18386 7336
rect 18616 7333 18644 7364
rect 18874 7352 18880 7404
rect 18932 7392 18938 7404
rect 19613 7395 19671 7401
rect 19613 7392 19625 7395
rect 18932 7364 19625 7392
rect 18932 7352 18938 7364
rect 19613 7361 19625 7364
rect 19659 7361 19671 7395
rect 19613 7355 19671 7361
rect 20070 7352 20076 7404
rect 20128 7352 20134 7404
rect 20714 7352 20720 7404
rect 20772 7352 20778 7404
rect 20824 7392 20852 7432
rect 21910 7420 21916 7472
rect 21968 7460 21974 7472
rect 22005 7463 22063 7469
rect 22005 7460 22017 7463
rect 21968 7432 22017 7460
rect 21968 7420 21974 7432
rect 22005 7429 22017 7432
rect 22051 7429 22063 7463
rect 30837 7463 30895 7469
rect 30837 7460 30849 7463
rect 22005 7423 22063 7429
rect 22572 7432 30849 7460
rect 22572 7392 22600 7432
rect 30837 7429 30849 7432
rect 30883 7429 30895 7463
rect 30837 7423 30895 7429
rect 32398 7420 32404 7472
rect 32456 7460 32462 7472
rect 32554 7463 32612 7469
rect 32554 7460 32566 7463
rect 32456 7432 32566 7460
rect 32456 7420 32462 7432
rect 32554 7429 32566 7432
rect 32600 7429 32612 7463
rect 32554 7423 32612 7429
rect 32674 7420 32680 7472
rect 32732 7420 32738 7472
rect 20824 7364 22600 7392
rect 22646 7352 22652 7404
rect 22704 7392 22710 7404
rect 23017 7395 23075 7401
rect 23017 7392 23029 7395
rect 22704 7364 23029 7392
rect 22704 7352 22710 7364
rect 23017 7361 23029 7364
rect 23063 7361 23075 7395
rect 23017 7355 23075 7361
rect 23750 7352 23756 7404
rect 23808 7392 23814 7404
rect 24673 7395 24731 7401
rect 24673 7392 24685 7395
rect 23808 7364 24685 7392
rect 23808 7352 23814 7364
rect 24673 7361 24685 7364
rect 24719 7361 24731 7395
rect 24673 7355 24731 7361
rect 24949 7395 25007 7401
rect 24949 7361 24961 7395
rect 24995 7392 25007 7395
rect 25498 7392 25504 7404
rect 24995 7364 25504 7392
rect 24995 7361 25007 7364
rect 24949 7355 25007 7361
rect 25498 7352 25504 7364
rect 25556 7392 25562 7404
rect 28810 7401 28816 7404
rect 25593 7395 25651 7401
rect 25593 7392 25605 7395
rect 25556 7364 25605 7392
rect 25556 7352 25562 7364
rect 25593 7361 25605 7364
rect 25639 7361 25651 7395
rect 25593 7355 25651 7361
rect 28804 7355 28816 7401
rect 28810 7352 28816 7355
rect 28868 7352 28874 7404
rect 32692 7392 32720 7420
rect 34348 7401 34376 7500
rect 37553 7463 37611 7469
rect 37553 7460 37565 7463
rect 36096 7432 37565 7460
rect 36096 7404 36124 7432
rect 37553 7429 37565 7432
rect 37599 7429 37611 7463
rect 37553 7423 37611 7429
rect 38746 7420 38752 7472
rect 38804 7420 38810 7472
rect 38930 7420 38936 7472
rect 38988 7420 38994 7472
rect 30944 7364 32720 7392
rect 34333 7395 34391 7401
rect 18601 7327 18659 7333
rect 18601 7293 18613 7327
rect 18647 7293 18659 7327
rect 18601 7287 18659 7293
rect 18785 7327 18843 7333
rect 18785 7293 18797 7327
rect 18831 7324 18843 7327
rect 19150 7324 19156 7336
rect 18831 7296 19156 7324
rect 18831 7293 18843 7296
rect 18785 7287 18843 7293
rect 18616 7256 18644 7287
rect 19150 7284 19156 7296
rect 19208 7284 19214 7336
rect 19981 7327 20039 7333
rect 19981 7293 19993 7327
rect 20027 7293 20039 7327
rect 19981 7287 20039 7293
rect 1627 7228 13124 7256
rect 14844 7228 18644 7256
rect 19996 7256 20024 7287
rect 20990 7284 20996 7336
rect 21048 7284 21054 7336
rect 23934 7284 23940 7336
rect 23992 7284 23998 7336
rect 28166 7284 28172 7336
rect 28224 7324 28230 7336
rect 28537 7327 28595 7333
rect 28537 7324 28549 7327
rect 28224 7296 28549 7324
rect 28224 7284 28230 7296
rect 28537 7293 28549 7296
rect 28583 7293 28595 7327
rect 28537 7287 28595 7293
rect 30466 7284 30472 7336
rect 30524 7324 30530 7336
rect 30944 7333 30972 7364
rect 34333 7361 34345 7395
rect 34379 7361 34391 7395
rect 34333 7355 34391 7361
rect 35526 7352 35532 7404
rect 35584 7352 35590 7404
rect 35618 7352 35624 7404
rect 35676 7392 35682 7404
rect 35713 7395 35771 7401
rect 35713 7392 35725 7395
rect 35676 7364 35725 7392
rect 35676 7352 35682 7364
rect 35713 7361 35725 7364
rect 35759 7361 35771 7395
rect 35713 7355 35771 7361
rect 36078 7352 36084 7404
rect 36136 7352 36142 7404
rect 39040 7401 39068 7500
rect 39298 7488 39304 7500
rect 39356 7488 39362 7540
rect 39485 7531 39543 7537
rect 39485 7497 39497 7531
rect 39531 7528 39543 7531
rect 40605 7531 40663 7537
rect 40605 7528 40617 7531
rect 39531 7500 40617 7528
rect 39531 7497 39543 7500
rect 39485 7491 39543 7497
rect 40605 7497 40617 7500
rect 40651 7497 40663 7531
rect 40605 7491 40663 7497
rect 41233 7531 41291 7537
rect 41233 7497 41245 7531
rect 41279 7528 41291 7531
rect 42518 7528 42524 7540
rect 41279 7500 42524 7528
rect 41279 7497 41291 7500
rect 41233 7491 41291 7497
rect 42518 7488 42524 7500
rect 42576 7488 42582 7540
rect 42705 7531 42763 7537
rect 42705 7497 42717 7531
rect 42751 7528 42763 7531
rect 42978 7528 42984 7540
rect 42751 7500 42984 7528
rect 42751 7497 42763 7500
rect 42705 7491 42763 7497
rect 42978 7488 42984 7500
rect 43036 7488 43042 7540
rect 44177 7531 44235 7537
rect 44177 7497 44189 7531
rect 44223 7528 44235 7531
rect 44266 7528 44272 7540
rect 44223 7500 44272 7528
rect 44223 7497 44235 7500
rect 44177 7491 44235 7497
rect 44266 7488 44272 7500
rect 44324 7488 44330 7540
rect 39316 7460 39344 7488
rect 40218 7460 40224 7472
rect 39316 7432 40224 7460
rect 37461 7395 37519 7401
rect 37461 7361 37473 7395
rect 37507 7361 37519 7395
rect 37461 7355 37519 7361
rect 39025 7395 39083 7401
rect 39025 7361 39037 7395
rect 39071 7361 39083 7395
rect 39025 7355 39083 7361
rect 39669 7395 39727 7401
rect 39669 7361 39681 7395
rect 39715 7361 39727 7395
rect 39669 7355 39727 7361
rect 30929 7327 30987 7333
rect 30929 7324 30941 7327
rect 30524 7296 30941 7324
rect 30524 7284 30530 7296
rect 30929 7293 30941 7296
rect 30975 7293 30987 7327
rect 30929 7287 30987 7293
rect 31202 7284 31208 7336
rect 31260 7324 31266 7336
rect 32309 7327 32367 7333
rect 32309 7324 32321 7327
rect 31260 7296 32321 7324
rect 31260 7284 31266 7296
rect 32309 7293 32321 7296
rect 32355 7293 32367 7327
rect 34241 7327 34299 7333
rect 34241 7324 34253 7327
rect 32309 7287 32367 7293
rect 33704 7296 34253 7324
rect 21269 7259 21327 7265
rect 21269 7256 21281 7259
rect 19996 7228 21281 7256
rect 1627 7225 1639 7228
rect 1581 7219 1639 7225
rect 5166 7148 5172 7200
rect 5224 7148 5230 7200
rect 12434 7148 12440 7200
rect 12492 7148 12498 7200
rect 13096 7188 13124 7228
rect 21269 7225 21281 7228
rect 21315 7225 21327 7259
rect 21269 7219 21327 7225
rect 14734 7188 14740 7200
rect 13096 7160 14740 7188
rect 14734 7148 14740 7160
rect 14792 7148 14798 7200
rect 14918 7148 14924 7200
rect 14976 7148 14982 7200
rect 15010 7148 15016 7200
rect 15068 7188 15074 7200
rect 19886 7188 19892 7200
rect 15068 7160 19892 7188
rect 15068 7148 15074 7160
rect 19886 7148 19892 7160
rect 19944 7148 19950 7200
rect 20073 7191 20131 7197
rect 20073 7157 20085 7191
rect 20119 7188 20131 7191
rect 20714 7188 20720 7200
rect 20119 7160 20720 7188
rect 20119 7157 20131 7160
rect 20073 7151 20131 7157
rect 20714 7148 20720 7160
rect 20772 7148 20778 7200
rect 20806 7148 20812 7200
rect 20864 7148 20870 7200
rect 22186 7148 22192 7200
rect 22244 7148 22250 7200
rect 25590 7148 25596 7200
rect 25648 7188 25654 7200
rect 25685 7191 25743 7197
rect 25685 7188 25697 7191
rect 25648 7160 25697 7188
rect 25648 7148 25654 7160
rect 25685 7157 25697 7160
rect 25731 7157 25743 7191
rect 25685 7151 25743 7157
rect 30006 7148 30012 7200
rect 30064 7188 30070 7200
rect 30377 7191 30435 7197
rect 30377 7188 30389 7191
rect 30064 7160 30389 7188
rect 30064 7148 30070 7160
rect 30377 7157 30389 7160
rect 30423 7157 30435 7191
rect 30377 7151 30435 7157
rect 33502 7148 33508 7200
rect 33560 7188 33566 7200
rect 33704 7197 33732 7296
rect 34241 7293 34253 7296
rect 34287 7293 34299 7327
rect 34241 7287 34299 7293
rect 35434 7284 35440 7336
rect 35492 7324 35498 7336
rect 35805 7327 35863 7333
rect 35805 7324 35817 7327
rect 35492 7296 35817 7324
rect 35492 7284 35498 7296
rect 35805 7293 35817 7296
rect 35851 7293 35863 7327
rect 35805 7287 35863 7293
rect 35894 7284 35900 7336
rect 35952 7324 35958 7336
rect 36354 7324 36360 7336
rect 35952 7296 36360 7324
rect 35952 7284 35958 7296
rect 36354 7284 36360 7296
rect 36412 7284 36418 7336
rect 37476 7324 37504 7355
rect 39684 7324 39712 7355
rect 39850 7352 39856 7404
rect 39908 7352 39914 7404
rect 39960 7401 39988 7432
rect 40218 7420 40224 7432
rect 40276 7420 40282 7472
rect 40405 7463 40463 7469
rect 40405 7429 40417 7463
rect 40451 7460 40463 7463
rect 40494 7460 40500 7472
rect 40451 7432 40500 7460
rect 40451 7429 40463 7432
rect 40405 7423 40463 7429
rect 40494 7420 40500 7432
rect 40552 7420 40558 7472
rect 39945 7395 40003 7401
rect 39945 7361 39957 7395
rect 39991 7361 40003 7395
rect 39945 7355 40003 7361
rect 41417 7395 41475 7401
rect 41417 7361 41429 7395
rect 41463 7361 41475 7395
rect 41417 7355 41475 7361
rect 40218 7324 40224 7336
rect 37476 7296 40224 7324
rect 40218 7284 40224 7296
rect 40276 7284 40282 7336
rect 38749 7259 38807 7265
rect 38749 7225 38761 7259
rect 38795 7256 38807 7259
rect 40310 7256 40316 7268
rect 38795 7228 40316 7256
rect 38795 7225 38807 7228
rect 38749 7219 38807 7225
rect 40310 7216 40316 7228
rect 40368 7216 40374 7268
rect 40773 7259 40831 7265
rect 40773 7225 40785 7259
rect 40819 7256 40831 7259
rect 41432 7256 41460 7355
rect 42610 7352 42616 7404
rect 42668 7352 42674 7404
rect 44358 7352 44364 7404
rect 44416 7352 44422 7404
rect 40819 7228 41460 7256
rect 40819 7225 40831 7228
rect 40773 7219 40831 7225
rect 33689 7191 33747 7197
rect 33689 7188 33701 7191
rect 33560 7160 33701 7188
rect 33560 7148 33566 7160
rect 33689 7157 33701 7160
rect 33735 7157 33747 7191
rect 33689 7151 33747 7157
rect 34701 7191 34759 7197
rect 34701 7157 34713 7191
rect 34747 7188 34759 7191
rect 35250 7188 35256 7200
rect 34747 7160 35256 7188
rect 34747 7157 34759 7160
rect 34701 7151 34759 7157
rect 35250 7148 35256 7160
rect 35308 7148 35314 7200
rect 36262 7148 36268 7200
rect 36320 7148 36326 7200
rect 39942 7148 39948 7200
rect 40000 7188 40006 7200
rect 40589 7191 40647 7197
rect 40589 7188 40601 7191
rect 40000 7160 40601 7188
rect 40000 7148 40006 7160
rect 40589 7157 40601 7160
rect 40635 7188 40647 7191
rect 41230 7188 41236 7200
rect 40635 7160 41236 7188
rect 40635 7157 40647 7160
rect 40589 7151 40647 7157
rect 41230 7148 41236 7160
rect 41288 7148 41294 7200
rect 1104 7098 44896 7120
rect 1104 7046 6423 7098
rect 6475 7046 6487 7098
rect 6539 7046 6551 7098
rect 6603 7046 6615 7098
rect 6667 7046 6679 7098
rect 6731 7046 17370 7098
rect 17422 7046 17434 7098
rect 17486 7046 17498 7098
rect 17550 7046 17562 7098
rect 17614 7046 17626 7098
rect 17678 7046 28317 7098
rect 28369 7046 28381 7098
rect 28433 7046 28445 7098
rect 28497 7046 28509 7098
rect 28561 7046 28573 7098
rect 28625 7046 39264 7098
rect 39316 7046 39328 7098
rect 39380 7046 39392 7098
rect 39444 7046 39456 7098
rect 39508 7046 39520 7098
rect 39572 7046 44896 7098
rect 1104 7024 44896 7046
rect 8570 6944 8576 6996
rect 8628 6944 8634 6996
rect 12526 6944 12532 6996
rect 12584 6984 12590 6996
rect 13722 6984 13728 6996
rect 12584 6956 13728 6984
rect 12584 6944 12590 6956
rect 13722 6944 13728 6956
rect 13780 6944 13786 6996
rect 14642 6944 14648 6996
rect 14700 6944 14706 6996
rect 17589 6987 17647 6993
rect 16960 6956 17448 6984
rect 11701 6919 11759 6925
rect 11701 6916 11713 6919
rect 11624 6888 11713 6916
rect 11624 6860 11652 6888
rect 11701 6885 11713 6888
rect 11747 6885 11759 6919
rect 11701 6879 11759 6885
rect 2685 6851 2743 6857
rect 2685 6817 2697 6851
rect 2731 6848 2743 6851
rect 3418 6848 3424 6860
rect 2731 6820 3424 6848
rect 2731 6817 2743 6820
rect 2685 6811 2743 6817
rect 3418 6808 3424 6820
rect 3476 6808 3482 6860
rect 3970 6808 3976 6860
rect 4028 6808 4034 6860
rect 11606 6808 11612 6860
rect 11664 6808 11670 6860
rect 11716 6820 12112 6848
rect 3988 6780 4016 6808
rect 7193 6783 7251 6789
rect 7193 6780 7205 6783
rect 3988 6752 7205 6780
rect 7193 6749 7205 6752
rect 7239 6780 7251 6783
rect 7926 6780 7932 6792
rect 7239 6752 7932 6780
rect 7239 6749 7251 6752
rect 7193 6743 7251 6749
rect 7926 6740 7932 6752
rect 7984 6780 7990 6792
rect 8662 6780 8668 6792
rect 7984 6752 8668 6780
rect 7984 6740 7990 6752
rect 8662 6740 8668 6752
rect 8720 6740 8726 6792
rect 9122 6740 9128 6792
rect 9180 6780 9186 6792
rect 9493 6783 9551 6789
rect 9493 6780 9505 6783
rect 9180 6752 9505 6780
rect 9180 6740 9186 6752
rect 9493 6749 9505 6752
rect 9539 6749 9551 6783
rect 9493 6743 9551 6749
rect 9766 6740 9772 6792
rect 9824 6740 9830 6792
rect 11716 6789 11744 6820
rect 11701 6783 11759 6789
rect 11701 6749 11713 6783
rect 11747 6749 11759 6783
rect 11701 6743 11759 6749
rect 11790 6740 11796 6792
rect 11848 6780 11854 6792
rect 11885 6783 11943 6789
rect 11885 6780 11897 6783
rect 11848 6752 11897 6780
rect 11848 6740 11854 6752
rect 11885 6749 11897 6752
rect 11931 6749 11943 6783
rect 11885 6743 11943 6749
rect 2501 6715 2559 6721
rect 2501 6681 2513 6715
rect 2547 6712 2559 6715
rect 2547 6684 3188 6712
rect 2547 6681 2559 6684
rect 2501 6675 2559 6681
rect 2130 6604 2136 6656
rect 2188 6604 2194 6656
rect 2593 6647 2651 6653
rect 2593 6613 2605 6647
rect 2639 6644 2651 6647
rect 2866 6644 2872 6656
rect 2639 6616 2872 6644
rect 2639 6613 2651 6616
rect 2593 6607 2651 6613
rect 2866 6604 2872 6616
rect 2924 6604 2930 6656
rect 3160 6644 3188 6684
rect 3234 6672 3240 6724
rect 3292 6712 3298 6724
rect 4218 6715 4276 6721
rect 4218 6712 4230 6715
rect 3292 6684 4230 6712
rect 3292 6672 3298 6684
rect 4218 6681 4230 6684
rect 4264 6681 4276 6715
rect 4218 6675 4276 6681
rect 7460 6715 7518 6721
rect 7460 6681 7472 6715
rect 7506 6712 7518 6715
rect 12084 6712 12112 6820
rect 14826 6808 14832 6860
rect 14884 6848 14890 6860
rect 15381 6851 15439 6857
rect 14884 6820 15332 6848
rect 14884 6808 14890 6820
rect 12250 6740 12256 6792
rect 12308 6780 12314 6792
rect 12345 6783 12403 6789
rect 12345 6780 12357 6783
rect 12308 6752 12357 6780
rect 12308 6740 12314 6752
rect 12345 6749 12357 6752
rect 12391 6749 12403 6783
rect 12345 6743 12403 6749
rect 12434 6740 12440 6792
rect 12492 6780 12498 6792
rect 12601 6783 12659 6789
rect 12601 6780 12613 6783
rect 12492 6752 12613 6780
rect 12492 6740 12498 6752
rect 12601 6749 12613 6752
rect 12647 6749 12659 6783
rect 12601 6743 12659 6749
rect 14274 6740 14280 6792
rect 14332 6780 14338 6792
rect 14918 6780 14924 6792
rect 14332 6752 14924 6780
rect 14332 6740 14338 6752
rect 14918 6740 14924 6752
rect 14976 6740 14982 6792
rect 15304 6789 15332 6820
rect 15381 6817 15393 6851
rect 15427 6848 15439 6851
rect 16960 6848 16988 6956
rect 17037 6919 17095 6925
rect 17037 6885 17049 6919
rect 17083 6885 17095 6919
rect 17037 6879 17095 6885
rect 15427 6820 16988 6848
rect 17052 6848 17080 6879
rect 17420 6848 17448 6956
rect 17589 6953 17601 6987
rect 17635 6984 17647 6987
rect 19334 6984 19340 6996
rect 17635 6956 19340 6984
rect 17635 6953 17647 6956
rect 17589 6947 17647 6953
rect 19334 6944 19340 6956
rect 19392 6944 19398 6996
rect 20901 6987 20959 6993
rect 20901 6953 20913 6987
rect 20947 6953 20959 6987
rect 20901 6947 20959 6953
rect 28629 6987 28687 6993
rect 28629 6953 28641 6987
rect 28675 6984 28687 6987
rect 28810 6984 28816 6996
rect 28675 6956 28816 6984
rect 28675 6953 28687 6956
rect 28629 6947 28687 6953
rect 18414 6876 18420 6928
rect 18472 6916 18478 6928
rect 20916 6916 20944 6947
rect 28810 6944 28816 6956
rect 28868 6944 28874 6996
rect 32401 6987 32459 6993
rect 32401 6953 32413 6987
rect 32447 6984 32459 6987
rect 32582 6984 32588 6996
rect 32447 6956 32588 6984
rect 32447 6953 32459 6956
rect 32401 6947 32459 6953
rect 32582 6944 32588 6956
rect 32640 6944 32646 6996
rect 39114 6944 39120 6996
rect 39172 6984 39178 6996
rect 39482 6984 39488 6996
rect 39172 6956 39488 6984
rect 39172 6944 39178 6956
rect 39482 6944 39488 6956
rect 39540 6944 39546 6996
rect 40034 6984 40040 6996
rect 39776 6956 40040 6984
rect 18472 6888 19012 6916
rect 20916 6888 21036 6916
rect 18472 6876 18478 6888
rect 17681 6851 17739 6857
rect 17681 6848 17693 6851
rect 17052 6820 17356 6848
rect 17420 6820 17693 6848
rect 15427 6817 15439 6820
rect 15381 6811 15439 6817
rect 15289 6783 15347 6789
rect 15289 6749 15301 6783
rect 15335 6749 15347 6783
rect 17218 6780 17224 6792
rect 17179 6752 17224 6780
rect 15289 6743 15347 6749
rect 17218 6740 17224 6752
rect 17276 6740 17282 6792
rect 17328 6780 17356 6820
rect 17681 6817 17693 6820
rect 17727 6848 17739 6851
rect 18782 6848 18788 6860
rect 17727 6820 18788 6848
rect 17727 6817 17739 6820
rect 17681 6811 17739 6817
rect 18782 6808 18788 6820
rect 18840 6808 18846 6860
rect 18874 6808 18880 6860
rect 18932 6808 18938 6860
rect 18984 6848 19012 6888
rect 19981 6851 20039 6857
rect 19981 6848 19993 6851
rect 18984 6820 19993 6848
rect 19981 6817 19993 6820
rect 20027 6817 20039 6851
rect 21008 6848 21036 6888
rect 19981 6811 20039 6817
rect 20088 6820 20944 6848
rect 21008 6820 21956 6848
rect 18141 6783 18199 6789
rect 18141 6780 18153 6783
rect 17328 6752 18153 6780
rect 18141 6749 18153 6752
rect 18187 6749 18199 6783
rect 18141 6743 18199 6749
rect 18325 6783 18383 6789
rect 18325 6749 18337 6783
rect 18371 6749 18383 6783
rect 18325 6743 18383 6749
rect 14458 6712 14464 6724
rect 7506 6684 10916 6712
rect 12084 6684 14464 6712
rect 7506 6681 7518 6684
rect 7460 6675 7518 6681
rect 5258 6644 5264 6656
rect 3160 6616 5264 6644
rect 5258 6604 5264 6616
rect 5316 6604 5322 6656
rect 5353 6647 5411 6653
rect 5353 6613 5365 6647
rect 5399 6644 5411 6647
rect 5534 6644 5540 6656
rect 5399 6616 5540 6644
rect 5399 6613 5411 6616
rect 5353 6607 5411 6613
rect 5534 6604 5540 6616
rect 5592 6644 5598 6656
rect 5994 6644 6000 6656
rect 5592 6616 6000 6644
rect 5592 6604 5598 6616
rect 5994 6604 6000 6616
rect 6052 6604 6058 6656
rect 9207 6647 9265 6653
rect 9207 6613 9219 6647
rect 9253 6644 9265 6647
rect 9398 6644 9404 6656
rect 9253 6616 9404 6644
rect 9253 6613 9265 6616
rect 9207 6607 9265 6613
rect 9398 6604 9404 6616
rect 9456 6604 9462 6656
rect 9674 6604 9680 6656
rect 9732 6604 9738 6656
rect 10888 6644 10916 6684
rect 14458 6672 14464 6684
rect 14516 6672 14522 6724
rect 15102 6672 15108 6724
rect 15160 6712 15166 6724
rect 18340 6712 18368 6743
rect 18414 6740 18420 6792
rect 18472 6740 18478 6792
rect 18506 6740 18512 6792
rect 18564 6740 18570 6792
rect 18598 6740 18604 6792
rect 18656 6780 18662 6792
rect 18693 6783 18751 6789
rect 18693 6780 18705 6783
rect 18656 6752 18705 6780
rect 18656 6740 18662 6752
rect 18693 6749 18705 6752
rect 18739 6749 18751 6783
rect 18693 6743 18751 6749
rect 19610 6740 19616 6792
rect 19668 6740 19674 6792
rect 19705 6783 19763 6789
rect 19705 6749 19717 6783
rect 19751 6780 19763 6783
rect 19886 6780 19892 6792
rect 19751 6752 19892 6780
rect 19751 6749 19763 6752
rect 19705 6743 19763 6749
rect 19886 6740 19892 6752
rect 19944 6740 19950 6792
rect 20088 6789 20116 6820
rect 20073 6783 20131 6789
rect 20073 6749 20085 6783
rect 20119 6749 20131 6783
rect 20073 6743 20131 6749
rect 20809 6783 20867 6789
rect 20809 6749 20821 6783
rect 20855 6749 20867 6783
rect 20916 6780 20944 6820
rect 20993 6783 21051 6789
rect 20993 6780 21005 6783
rect 20916 6752 21005 6780
rect 20809 6743 20867 6749
rect 20993 6749 21005 6752
rect 21039 6780 21051 6783
rect 21729 6783 21787 6789
rect 21729 6780 21741 6783
rect 21039 6752 21741 6780
rect 21039 6749 21051 6752
rect 20993 6743 21051 6749
rect 21729 6749 21741 6752
rect 21775 6749 21787 6783
rect 21729 6743 21787 6749
rect 20088 6712 20116 6743
rect 15160 6684 17264 6712
rect 18340 6684 20116 6712
rect 15160 6672 15166 6684
rect 12802 6644 12808 6656
rect 10888 6616 12808 6644
rect 12802 6604 12808 6616
rect 12860 6644 12866 6656
rect 13630 6644 13636 6656
rect 12860 6616 13636 6644
rect 12860 6604 12866 6616
rect 13630 6604 13636 6616
rect 13688 6604 13694 6656
rect 14642 6604 14648 6656
rect 14700 6604 14706 6656
rect 14829 6647 14887 6653
rect 14829 6613 14841 6647
rect 14875 6644 14887 6647
rect 15286 6644 15292 6656
rect 14875 6616 15292 6644
rect 14875 6613 14887 6616
rect 14829 6607 14887 6613
rect 15286 6604 15292 6616
rect 15344 6604 15350 6656
rect 17236 6653 17264 6684
rect 20714 6672 20720 6724
rect 20772 6712 20778 6724
rect 20824 6712 20852 6743
rect 21634 6712 21640 6724
rect 20772 6684 21640 6712
rect 20772 6672 20778 6684
rect 21634 6672 21640 6684
rect 21692 6672 21698 6724
rect 17221 6647 17279 6653
rect 17221 6613 17233 6647
rect 17267 6644 17279 6647
rect 18506 6644 18512 6656
rect 17267 6616 18512 6644
rect 17267 6613 17279 6616
rect 17221 6607 17279 6613
rect 18506 6604 18512 6616
rect 18564 6604 18570 6656
rect 19429 6647 19487 6653
rect 19429 6613 19441 6647
rect 19475 6644 19487 6647
rect 20990 6644 20996 6656
rect 19475 6616 20996 6644
rect 19475 6613 19487 6616
rect 19429 6607 19487 6613
rect 20990 6604 20996 6616
rect 21048 6604 21054 6656
rect 21450 6604 21456 6656
rect 21508 6604 21514 6656
rect 21744 6644 21772 6743
rect 21818 6740 21824 6792
rect 21876 6740 21882 6792
rect 21928 6789 21956 6820
rect 32674 6808 32680 6860
rect 32732 6848 32738 6860
rect 32953 6851 33011 6857
rect 32953 6848 32965 6851
rect 32732 6820 32965 6848
rect 32732 6808 32738 6820
rect 32953 6817 32965 6820
rect 32999 6817 33011 6851
rect 32953 6811 33011 6817
rect 33042 6808 33048 6860
rect 33100 6848 33106 6860
rect 34422 6848 34428 6860
rect 33100 6820 34428 6848
rect 33100 6808 33106 6820
rect 21913 6783 21971 6789
rect 21913 6749 21925 6783
rect 21959 6749 21971 6783
rect 21913 6743 21971 6749
rect 22002 6740 22008 6792
rect 22060 6780 22066 6792
rect 22097 6783 22155 6789
rect 22097 6780 22109 6783
rect 22060 6752 22109 6780
rect 22060 6740 22066 6752
rect 22097 6749 22109 6752
rect 22143 6749 22155 6783
rect 22097 6743 22155 6749
rect 22646 6740 22652 6792
rect 22704 6740 22710 6792
rect 24026 6740 24032 6792
rect 24084 6740 24090 6792
rect 24578 6740 24584 6792
rect 24636 6740 24642 6792
rect 28169 6783 28227 6789
rect 28169 6749 28181 6783
rect 28215 6749 28227 6783
rect 28169 6743 28227 6749
rect 28813 6783 28871 6789
rect 28813 6749 28825 6783
rect 28859 6780 28871 6783
rect 30006 6780 30012 6792
rect 28859 6752 30012 6780
rect 28859 6749 28871 6752
rect 28813 6743 28871 6749
rect 24857 6715 24915 6721
rect 24857 6681 24869 6715
rect 24903 6681 24915 6715
rect 24857 6675 24915 6681
rect 22741 6647 22799 6653
rect 22741 6644 22753 6647
rect 21744 6616 22753 6644
rect 22741 6613 22753 6616
rect 22787 6613 22799 6647
rect 22741 6607 22799 6613
rect 23845 6647 23903 6653
rect 23845 6613 23857 6647
rect 23891 6644 23903 6647
rect 24872 6644 24900 6675
rect 25590 6672 25596 6724
rect 25648 6672 25654 6724
rect 28184 6712 28212 6743
rect 30006 6740 30012 6752
rect 30064 6740 30070 6792
rect 30742 6740 30748 6792
rect 30800 6780 30806 6792
rect 31205 6783 31263 6789
rect 31205 6780 31217 6783
rect 30800 6752 31217 6780
rect 30800 6740 30806 6752
rect 31205 6749 31217 6752
rect 31251 6749 31263 6783
rect 31205 6743 31263 6749
rect 32769 6783 32827 6789
rect 32769 6749 32781 6783
rect 32815 6780 32827 6783
rect 33502 6780 33508 6792
rect 32815 6752 33508 6780
rect 32815 6749 32827 6752
rect 32769 6743 32827 6749
rect 33502 6740 33508 6752
rect 33560 6740 33566 6792
rect 33612 6789 33640 6820
rect 34422 6808 34428 6820
rect 34480 6808 34486 6860
rect 35618 6848 35624 6860
rect 35544 6820 35624 6848
rect 33597 6783 33655 6789
rect 33597 6749 33609 6783
rect 33643 6749 33655 6783
rect 33597 6743 33655 6749
rect 33686 6740 33692 6792
rect 33744 6780 33750 6792
rect 33965 6783 34023 6789
rect 33965 6780 33977 6783
rect 33744 6752 33977 6780
rect 33744 6740 33750 6752
rect 33965 6749 33977 6752
rect 34011 6749 34023 6783
rect 33965 6743 34023 6749
rect 35250 6740 35256 6792
rect 35308 6740 35314 6792
rect 35434 6789 35440 6792
rect 35401 6783 35440 6789
rect 35401 6749 35413 6783
rect 35401 6743 35440 6749
rect 35434 6740 35440 6743
rect 35492 6740 35498 6792
rect 35544 6789 35572 6820
rect 35618 6808 35624 6820
rect 35676 6808 35682 6860
rect 37458 6808 37464 6860
rect 37516 6848 37522 6860
rect 39776 6848 39804 6956
rect 40034 6944 40040 6956
rect 40092 6944 40098 6996
rect 40218 6944 40224 6996
rect 40276 6984 40282 6996
rect 43990 6984 43996 6996
rect 40276 6956 43996 6984
rect 40276 6944 40282 6956
rect 43990 6944 43996 6956
rect 44048 6944 44054 6996
rect 39850 6876 39856 6928
rect 39908 6916 39914 6928
rect 39908 6888 39988 6916
rect 39908 6876 39914 6888
rect 37516 6820 39804 6848
rect 39960 6848 39988 6888
rect 40494 6876 40500 6928
rect 40552 6916 40558 6928
rect 40552 6888 41184 6916
rect 40552 6876 40558 6888
rect 39960 6820 40080 6848
rect 37516 6808 37522 6820
rect 35529 6783 35587 6789
rect 35529 6749 35541 6783
rect 35575 6749 35587 6783
rect 35529 6743 35587 6749
rect 35759 6783 35817 6789
rect 35759 6749 35771 6783
rect 35805 6780 35817 6783
rect 35894 6780 35900 6792
rect 35805 6752 35900 6780
rect 35805 6749 35817 6752
rect 35759 6743 35817 6749
rect 35894 6740 35900 6752
rect 35952 6740 35958 6792
rect 38289 6783 38347 6789
rect 38289 6749 38301 6783
rect 38335 6749 38347 6783
rect 38289 6743 38347 6749
rect 29730 6712 29736 6724
rect 28184 6684 29736 6712
rect 29730 6672 29736 6684
rect 29788 6672 29794 6724
rect 32582 6672 32588 6724
rect 32640 6712 32646 6724
rect 32861 6715 32919 6721
rect 32861 6712 32873 6715
rect 32640 6684 32873 6712
rect 32640 6672 32646 6684
rect 32861 6681 32873 6684
rect 32907 6681 32919 6715
rect 32861 6675 32919 6681
rect 33134 6672 33140 6724
rect 33192 6712 33198 6724
rect 33781 6715 33839 6721
rect 33781 6712 33793 6715
rect 33192 6684 33793 6712
rect 33192 6672 33198 6684
rect 33781 6681 33793 6684
rect 33827 6681 33839 6715
rect 33781 6675 33839 6681
rect 33873 6715 33931 6721
rect 33873 6681 33885 6715
rect 33919 6681 33931 6715
rect 33873 6675 33931 6681
rect 35621 6715 35679 6721
rect 35621 6681 35633 6715
rect 35667 6712 35679 6715
rect 36078 6712 36084 6724
rect 35667 6684 36084 6712
rect 35667 6681 35679 6684
rect 35621 6675 35679 6681
rect 23891 6616 24900 6644
rect 23891 6613 23903 6616
rect 23845 6607 23903 6613
rect 25222 6604 25228 6656
rect 25280 6644 25286 6656
rect 26329 6647 26387 6653
rect 26329 6644 26341 6647
rect 25280 6616 26341 6644
rect 25280 6604 25286 6616
rect 26329 6613 26341 6616
rect 26375 6613 26387 6647
rect 26329 6607 26387 6613
rect 27982 6604 27988 6656
rect 28040 6604 28046 6656
rect 31297 6647 31355 6653
rect 31297 6613 31309 6647
rect 31343 6644 31355 6647
rect 32766 6644 32772 6656
rect 31343 6616 32772 6644
rect 31343 6613 31355 6616
rect 31297 6607 31355 6613
rect 32766 6604 32772 6616
rect 32824 6604 32830 6656
rect 33686 6604 33692 6656
rect 33744 6644 33750 6656
rect 33888 6644 33916 6675
rect 36078 6672 36084 6684
rect 36136 6672 36142 6724
rect 38304 6712 38332 6743
rect 38470 6740 38476 6792
rect 38528 6740 38534 6792
rect 39942 6780 39948 6792
rect 38856 6752 39948 6780
rect 38856 6712 38884 6752
rect 39942 6740 39948 6752
rect 40000 6740 40006 6792
rect 38304 6684 38884 6712
rect 38930 6672 38936 6724
rect 38988 6672 38994 6724
rect 40052 6721 40080 6820
rect 40126 6808 40132 6860
rect 40184 6848 40190 6860
rect 40770 6848 40776 6860
rect 40184 6820 40776 6848
rect 40184 6808 40190 6820
rect 40770 6808 40776 6820
rect 40828 6848 40834 6860
rect 41156 6857 41184 6888
rect 40957 6851 41015 6857
rect 40957 6848 40969 6851
rect 40828 6820 40969 6848
rect 40828 6808 40834 6820
rect 40957 6817 40969 6820
rect 41003 6817 41015 6851
rect 40957 6811 41015 6817
rect 41141 6851 41199 6857
rect 41141 6817 41153 6851
rect 41187 6817 41199 6851
rect 41141 6811 41199 6817
rect 41230 6808 41236 6860
rect 41288 6848 41294 6860
rect 41693 6851 41751 6857
rect 41693 6848 41705 6851
rect 41288 6820 41705 6848
rect 41288 6808 41294 6820
rect 41693 6817 41705 6820
rect 41739 6817 41751 6851
rect 41693 6811 41751 6817
rect 40862 6740 40868 6792
rect 40920 6740 40926 6792
rect 41601 6783 41659 6789
rect 41601 6780 41613 6783
rect 41386 6752 41613 6780
rect 40310 6721 40316 6724
rect 40037 6715 40095 6721
rect 39224 6684 39988 6712
rect 33744 6616 33916 6644
rect 33744 6604 33750 6616
rect 34146 6604 34152 6656
rect 34204 6604 34210 6656
rect 34974 6604 34980 6656
rect 35032 6644 35038 6656
rect 35897 6647 35955 6653
rect 35897 6644 35909 6647
rect 35032 6616 35909 6644
rect 35032 6604 35038 6616
rect 35897 6613 35909 6616
rect 35943 6613 35955 6647
rect 35897 6607 35955 6613
rect 38381 6647 38439 6653
rect 38381 6613 38393 6647
rect 38427 6644 38439 6647
rect 39133 6647 39191 6653
rect 39133 6644 39145 6647
rect 38427 6616 39145 6644
rect 38427 6613 38439 6616
rect 38381 6607 38439 6613
rect 39133 6613 39145 6616
rect 39179 6644 39191 6647
rect 39224 6644 39252 6684
rect 39179 6616 39252 6644
rect 39301 6647 39359 6653
rect 39179 6613 39191 6616
rect 39133 6607 39191 6613
rect 39301 6613 39313 6647
rect 39347 6644 39359 6647
rect 39666 6644 39672 6656
rect 39347 6616 39672 6644
rect 39347 6613 39359 6616
rect 39301 6607 39359 6613
rect 39666 6604 39672 6616
rect 39724 6604 39730 6656
rect 39960 6644 39988 6684
rect 40037 6681 40049 6715
rect 40083 6681 40095 6715
rect 40037 6675 40095 6681
rect 40253 6715 40316 6721
rect 40253 6681 40265 6715
rect 40299 6681 40316 6715
rect 40253 6675 40316 6681
rect 40310 6672 40316 6675
rect 40368 6672 40374 6724
rect 41386 6712 41414 6752
rect 41601 6749 41613 6752
rect 41647 6749 41659 6783
rect 41601 6743 41659 6749
rect 42245 6783 42303 6789
rect 42245 6749 42257 6783
rect 42291 6780 42303 6783
rect 42610 6780 42616 6792
rect 42291 6752 42616 6780
rect 42291 6749 42303 6752
rect 42245 6743 42303 6749
rect 42610 6740 42616 6752
rect 42668 6740 42674 6792
rect 40420 6684 41414 6712
rect 40420 6656 40448 6684
rect 40126 6644 40132 6656
rect 39960 6616 40132 6644
rect 40126 6604 40132 6616
rect 40184 6604 40190 6656
rect 40402 6604 40408 6656
rect 40460 6604 40466 6656
rect 40678 6604 40684 6656
rect 40736 6644 40742 6656
rect 41141 6647 41199 6653
rect 41141 6644 41153 6647
rect 40736 6616 41153 6644
rect 40736 6604 40742 6616
rect 41141 6613 41153 6616
rect 41187 6613 41199 6647
rect 41141 6607 41199 6613
rect 42242 6604 42248 6656
rect 42300 6644 42306 6656
rect 42337 6647 42395 6653
rect 42337 6644 42349 6647
rect 42300 6616 42349 6644
rect 42300 6604 42306 6616
rect 42337 6613 42349 6616
rect 42383 6613 42395 6647
rect 42337 6607 42395 6613
rect 1104 6554 45051 6576
rect 1104 6502 11896 6554
rect 11948 6502 11960 6554
rect 12012 6502 12024 6554
rect 12076 6502 12088 6554
rect 12140 6502 12152 6554
rect 12204 6502 22843 6554
rect 22895 6502 22907 6554
rect 22959 6502 22971 6554
rect 23023 6502 23035 6554
rect 23087 6502 23099 6554
rect 23151 6502 33790 6554
rect 33842 6502 33854 6554
rect 33906 6502 33918 6554
rect 33970 6502 33982 6554
rect 34034 6502 34046 6554
rect 34098 6502 44737 6554
rect 44789 6502 44801 6554
rect 44853 6502 44865 6554
rect 44917 6502 44929 6554
rect 44981 6502 44993 6554
rect 45045 6502 45051 6554
rect 1104 6480 45051 6502
rect 2866 6400 2872 6452
rect 2924 6400 2930 6452
rect 4709 6443 4767 6449
rect 4709 6409 4721 6443
rect 4755 6409 4767 6443
rect 4709 6403 4767 6409
rect 6840 6412 9260 6440
rect 4724 6372 4752 6403
rect 2746 6344 4752 6372
rect 934 6264 940 6316
rect 992 6304 998 6316
rect 1765 6307 1823 6313
rect 1765 6304 1777 6307
rect 992 6276 1777 6304
rect 992 6264 998 6276
rect 1765 6273 1777 6276
rect 1811 6273 1823 6307
rect 1765 6267 1823 6273
rect 2314 6264 2320 6316
rect 2372 6304 2378 6316
rect 2746 6304 2774 6344
rect 2372 6276 2774 6304
rect 2372 6264 2378 6276
rect 3326 6264 3332 6316
rect 3384 6264 3390 6316
rect 3596 6307 3654 6313
rect 3596 6273 3608 6307
rect 3642 6304 3654 6307
rect 6840 6304 6868 6412
rect 6914 6332 6920 6384
rect 6972 6372 6978 6384
rect 8174 6375 8232 6381
rect 8174 6372 8186 6375
rect 6972 6344 8186 6372
rect 6972 6332 6978 6344
rect 8174 6341 8186 6344
rect 8220 6341 8232 6375
rect 9232 6372 9260 6412
rect 9306 6400 9312 6452
rect 9364 6400 9370 6452
rect 11146 6400 11152 6452
rect 11204 6400 11210 6452
rect 12526 6440 12532 6452
rect 12176 6412 12532 6440
rect 10502 6372 10508 6384
rect 9232 6344 10508 6372
rect 8174 6335 8232 6341
rect 10502 6332 10508 6344
rect 10560 6332 10566 6384
rect 12176 6381 12204 6412
rect 12526 6400 12532 6412
rect 12584 6400 12590 6452
rect 12618 6400 12624 6452
rect 12676 6440 12682 6452
rect 13541 6443 13599 6449
rect 13541 6440 13553 6443
rect 12676 6412 13553 6440
rect 12676 6400 12682 6412
rect 13541 6409 13553 6412
rect 13587 6409 13599 6443
rect 13541 6403 13599 6409
rect 13722 6400 13728 6452
rect 13780 6440 13786 6452
rect 15029 6443 15087 6449
rect 15029 6440 15041 6443
rect 13780 6412 15041 6440
rect 13780 6400 13786 6412
rect 15029 6409 15041 6412
rect 15075 6409 15087 6443
rect 19886 6440 19892 6452
rect 15029 6403 15087 6409
rect 15120 6412 19892 6440
rect 12161 6375 12219 6381
rect 12161 6341 12173 6375
rect 12207 6341 12219 6375
rect 12161 6335 12219 6341
rect 12377 6375 12435 6381
rect 12377 6341 12389 6375
rect 12423 6372 12435 6375
rect 13170 6372 13176 6384
rect 12423 6344 13176 6372
rect 12423 6341 12435 6344
rect 12377 6335 12435 6341
rect 13170 6332 13176 6344
rect 13228 6332 13234 6384
rect 13357 6375 13415 6381
rect 13357 6372 13369 6375
rect 13280 6344 13369 6372
rect 3642 6276 6868 6304
rect 3642 6273 3654 6276
rect 3596 6267 3654 6273
rect 7926 6264 7932 6316
rect 7984 6264 7990 6316
rect 8662 6264 8668 6316
rect 8720 6304 8726 6316
rect 9582 6304 9588 6316
rect 8720 6276 9588 6304
rect 8720 6264 8726 6276
rect 9582 6264 9588 6276
rect 9640 6304 9646 6316
rect 9769 6307 9827 6313
rect 9769 6304 9781 6307
rect 9640 6276 9781 6304
rect 9640 6264 9646 6276
rect 9769 6273 9781 6276
rect 9815 6273 9827 6307
rect 9769 6267 9827 6273
rect 10036 6307 10094 6313
rect 10036 6273 10048 6307
rect 10082 6304 10094 6307
rect 12066 6304 12072 6316
rect 10082 6276 12072 6304
rect 10082 6273 10094 6276
rect 10036 6267 10094 6273
rect 12066 6264 12072 6276
rect 12124 6264 12130 6316
rect 13280 6236 13308 6344
rect 13357 6341 13369 6344
rect 13403 6341 13415 6375
rect 13357 6335 13415 6341
rect 13446 6332 13452 6384
rect 13504 6372 13510 6384
rect 14001 6375 14059 6381
rect 14001 6372 14013 6375
rect 13504 6344 14013 6372
rect 13504 6332 13510 6344
rect 14001 6341 14013 6344
rect 14047 6372 14059 6375
rect 14274 6372 14280 6384
rect 14047 6344 14280 6372
rect 14047 6341 14059 6344
rect 14001 6335 14059 6341
rect 14274 6332 14280 6344
rect 14332 6332 14338 6384
rect 14826 6332 14832 6384
rect 14884 6332 14890 6384
rect 14918 6332 14924 6384
rect 14976 6372 14982 6384
rect 15120 6372 15148 6412
rect 19886 6400 19892 6412
rect 19944 6400 19950 6452
rect 20257 6443 20315 6449
rect 20257 6409 20269 6443
rect 20303 6440 20315 6443
rect 20806 6440 20812 6452
rect 20303 6412 20812 6440
rect 20303 6409 20315 6412
rect 20257 6403 20315 6409
rect 20806 6400 20812 6412
rect 20864 6400 20870 6452
rect 20990 6400 20996 6452
rect 21048 6440 21054 6452
rect 21910 6440 21916 6452
rect 21048 6412 21916 6440
rect 21048 6400 21054 6412
rect 21910 6400 21916 6412
rect 21968 6400 21974 6452
rect 22646 6400 22652 6452
rect 22704 6440 22710 6452
rect 23385 6443 23443 6449
rect 23385 6440 23397 6443
rect 22704 6412 23397 6440
rect 22704 6400 22710 6412
rect 23385 6409 23397 6412
rect 23431 6409 23443 6443
rect 23385 6403 23443 6409
rect 24026 6400 24032 6452
rect 24084 6440 24090 6452
rect 24857 6443 24915 6449
rect 24857 6440 24869 6443
rect 24084 6412 24869 6440
rect 24084 6400 24090 6412
rect 24857 6409 24869 6412
rect 24903 6409 24915 6443
rect 24857 6403 24915 6409
rect 25222 6400 25228 6452
rect 25280 6400 25286 6452
rect 32858 6400 32864 6452
rect 32916 6440 32922 6452
rect 34330 6440 34336 6452
rect 32916 6412 34336 6440
rect 32916 6400 32922 6412
rect 34330 6400 34336 6412
rect 34388 6400 34394 6452
rect 35434 6400 35440 6452
rect 35492 6440 35498 6452
rect 38470 6440 38476 6452
rect 35492 6412 38476 6440
rect 35492 6400 35498 6412
rect 38470 6400 38476 6412
rect 38528 6440 38534 6452
rect 38565 6443 38623 6449
rect 38565 6440 38577 6443
rect 38528 6412 38577 6440
rect 38528 6400 38534 6412
rect 38565 6409 38577 6412
rect 38611 6409 38623 6443
rect 38565 6403 38623 6409
rect 39482 6400 39488 6452
rect 39540 6440 39546 6452
rect 40862 6440 40868 6452
rect 39540 6412 40868 6440
rect 39540 6400 39546 6412
rect 40862 6400 40868 6412
rect 40920 6400 40926 6452
rect 14976 6344 15148 6372
rect 17681 6375 17739 6381
rect 14976 6332 14982 6344
rect 17681 6341 17693 6375
rect 17727 6372 17739 6375
rect 18414 6372 18420 6384
rect 17727 6344 18420 6372
rect 17727 6341 17739 6344
rect 17681 6335 17739 6341
rect 18414 6332 18420 6344
rect 18472 6332 18478 6384
rect 18598 6332 18604 6384
rect 18656 6372 18662 6384
rect 18877 6375 18935 6381
rect 18877 6372 18889 6375
rect 18656 6344 18889 6372
rect 18656 6332 18662 6344
rect 18877 6341 18889 6344
rect 18923 6372 18935 6375
rect 18923 6344 20944 6372
rect 18923 6341 18935 6344
rect 18877 6335 18935 6341
rect 14090 6264 14096 6316
rect 14148 6304 14154 6316
rect 14185 6307 14243 6313
rect 14185 6304 14197 6307
rect 14148 6276 14197 6304
rect 14148 6264 14154 6276
rect 14185 6273 14197 6276
rect 14231 6273 14243 6307
rect 14185 6267 14243 6273
rect 18782 6264 18788 6316
rect 18840 6304 18846 6316
rect 18840 6276 19656 6304
rect 18840 6264 18846 6276
rect 13354 6236 13360 6248
rect 13280 6208 13360 6236
rect 13354 6196 13360 6208
rect 13412 6196 13418 6248
rect 17770 6196 17776 6248
rect 17828 6196 17834 6248
rect 17957 6239 18015 6245
rect 17957 6205 17969 6239
rect 18003 6236 18015 6239
rect 18322 6236 18328 6248
rect 18003 6208 18328 6236
rect 18003 6205 18015 6208
rect 17957 6199 18015 6205
rect 18322 6196 18328 6208
rect 18380 6196 18386 6248
rect 18966 6196 18972 6248
rect 19024 6196 19030 6248
rect 19150 6196 19156 6248
rect 19208 6196 19214 6248
rect 19628 6236 19656 6276
rect 19702 6264 19708 6316
rect 19760 6264 19766 6316
rect 19886 6264 19892 6316
rect 19944 6264 19950 6316
rect 19978 6264 19984 6316
rect 20036 6264 20042 6316
rect 20916 6313 20944 6344
rect 21450 6332 21456 6384
rect 21508 6372 21514 6384
rect 22250 6375 22308 6381
rect 22250 6372 22262 6375
rect 21508 6344 22262 6372
rect 21508 6332 21514 6344
rect 22250 6341 22262 6344
rect 22296 6341 22308 6375
rect 22250 6335 22308 6341
rect 20073 6307 20131 6313
rect 20073 6273 20085 6307
rect 20119 6273 20131 6307
rect 20073 6267 20131 6273
rect 20901 6307 20959 6313
rect 20901 6273 20913 6307
rect 20947 6273 20959 6307
rect 20901 6267 20959 6273
rect 20088 6236 20116 6267
rect 21542 6264 21548 6316
rect 21600 6304 21606 6316
rect 22005 6307 22063 6313
rect 22005 6304 22017 6307
rect 21600 6276 22017 6304
rect 21600 6264 21606 6276
rect 22005 6273 22017 6276
rect 22051 6273 22063 6307
rect 22005 6267 22063 6273
rect 24213 6307 24271 6313
rect 24213 6273 24225 6307
rect 24259 6304 24271 6307
rect 25240 6304 25268 6400
rect 27709 6375 27767 6381
rect 27709 6372 27721 6375
rect 24259 6276 25268 6304
rect 25332 6344 27721 6372
rect 24259 6273 24271 6276
rect 24213 6267 24271 6273
rect 25332 6248 25360 6344
rect 27709 6341 27721 6344
rect 27755 6341 27767 6375
rect 27709 6335 27767 6341
rect 27982 6332 27988 6384
rect 28040 6372 28046 6384
rect 28782 6375 28840 6381
rect 28782 6372 28794 6375
rect 28040 6344 28794 6372
rect 28040 6332 28046 6344
rect 28782 6341 28794 6344
rect 28828 6341 28840 6375
rect 28782 6335 28840 6341
rect 32769 6375 32827 6381
rect 32769 6341 32781 6375
rect 32815 6372 32827 6375
rect 36262 6372 36268 6384
rect 32815 6344 35112 6372
rect 32815 6341 32827 6344
rect 32769 6335 32827 6341
rect 27617 6307 27675 6313
rect 27617 6273 27629 6307
rect 27663 6304 27675 6307
rect 27890 6304 27896 6316
rect 27663 6276 27896 6304
rect 27663 6273 27675 6276
rect 27617 6267 27675 6273
rect 27890 6264 27896 6276
rect 27948 6264 27954 6316
rect 31481 6307 31539 6313
rect 31481 6273 31493 6307
rect 31527 6273 31539 6307
rect 31481 6267 31539 6273
rect 31665 6307 31723 6313
rect 31665 6273 31677 6307
rect 31711 6273 31723 6307
rect 31665 6267 31723 6273
rect 31757 6307 31815 6313
rect 31757 6273 31769 6307
rect 31803 6304 31815 6307
rect 31803 6276 32168 6304
rect 31803 6273 31815 6276
rect 31757 6267 31815 6273
rect 19628 6208 20116 6236
rect 20346 6196 20352 6248
rect 20404 6236 20410 6248
rect 20993 6239 21051 6245
rect 20993 6236 21005 6239
rect 20404 6208 21005 6236
rect 20404 6196 20410 6208
rect 20993 6205 21005 6208
rect 21039 6236 21051 6239
rect 21174 6236 21180 6248
rect 21039 6208 21180 6236
rect 21039 6205 21051 6208
rect 20993 6199 21051 6205
rect 21174 6196 21180 6208
rect 21232 6196 21238 6248
rect 25314 6196 25320 6248
rect 25372 6196 25378 6248
rect 25501 6239 25559 6245
rect 25501 6205 25513 6239
rect 25547 6236 25559 6239
rect 26142 6236 26148 6248
rect 25547 6208 26148 6236
rect 25547 6205 25559 6208
rect 25501 6199 25559 6205
rect 11698 6128 11704 6180
rect 11756 6168 11762 6180
rect 12526 6168 12532 6180
rect 11756 6140 12532 6168
rect 11756 6128 11762 6140
rect 12526 6128 12532 6140
rect 12584 6128 12590 6180
rect 12986 6128 12992 6180
rect 13044 6128 13050 6180
rect 14369 6171 14427 6177
rect 14369 6168 14381 6171
rect 13372 6140 14381 6168
rect 12345 6103 12403 6109
rect 12345 6069 12357 6103
rect 12391 6100 12403 6103
rect 13170 6100 13176 6112
rect 12391 6072 13176 6100
rect 12391 6069 12403 6072
rect 12345 6063 12403 6069
rect 13170 6060 13176 6072
rect 13228 6060 13234 6112
rect 13372 6109 13400 6140
rect 14369 6137 14381 6140
rect 14415 6137 14427 6171
rect 14369 6131 14427 6137
rect 14642 6128 14648 6180
rect 14700 6168 14706 6180
rect 20806 6168 20812 6180
rect 14700 6140 20812 6168
rect 14700 6128 14706 6140
rect 20806 6128 20812 6140
rect 20864 6128 20870 6180
rect 20898 6128 20904 6180
rect 20956 6168 20962 6180
rect 21269 6171 21327 6177
rect 21269 6168 21281 6171
rect 20956 6140 21281 6168
rect 20956 6128 20962 6140
rect 21269 6137 21281 6140
rect 21315 6137 21327 6171
rect 24305 6171 24363 6177
rect 24305 6168 24317 6171
rect 21269 6131 21327 6137
rect 23216 6140 24317 6168
rect 13357 6103 13415 6109
rect 13357 6069 13369 6103
rect 13403 6069 13415 6103
rect 13357 6063 13415 6069
rect 14090 6060 14096 6112
rect 14148 6100 14154 6112
rect 14918 6100 14924 6112
rect 14148 6072 14924 6100
rect 14148 6060 14154 6072
rect 14918 6060 14924 6072
rect 14976 6100 14982 6112
rect 15013 6103 15071 6109
rect 15013 6100 15025 6103
rect 14976 6072 15025 6100
rect 14976 6060 14982 6072
rect 15013 6069 15025 6072
rect 15059 6069 15071 6103
rect 15013 6063 15071 6069
rect 15197 6103 15255 6109
rect 15197 6069 15209 6103
rect 15243 6100 15255 6103
rect 15286 6100 15292 6112
rect 15243 6072 15292 6100
rect 15243 6069 15255 6072
rect 15197 6063 15255 6069
rect 15286 6060 15292 6072
rect 15344 6060 15350 6112
rect 16022 6060 16028 6112
rect 16080 6100 16086 6112
rect 17313 6103 17371 6109
rect 17313 6100 17325 6103
rect 16080 6072 17325 6100
rect 16080 6060 16086 6072
rect 17313 6069 17325 6072
rect 17359 6069 17371 6103
rect 17313 6063 17371 6069
rect 18509 6103 18567 6109
rect 18509 6069 18521 6103
rect 18555 6100 18567 6103
rect 19242 6100 19248 6112
rect 18555 6072 19248 6100
rect 18555 6069 18567 6072
rect 18509 6063 18567 6069
rect 19242 6060 19248 6072
rect 19300 6060 19306 6112
rect 19702 6060 19708 6112
rect 19760 6100 19766 6112
rect 23216 6100 23244 6140
rect 24305 6137 24317 6140
rect 24351 6137 24363 6171
rect 24305 6131 24363 6137
rect 24394 6128 24400 6180
rect 24452 6168 24458 6180
rect 25516 6168 25544 6199
rect 26142 6196 26148 6208
rect 26200 6196 26206 6248
rect 27801 6239 27859 6245
rect 27801 6205 27813 6239
rect 27847 6236 27859 6239
rect 27982 6236 27988 6248
rect 27847 6208 27988 6236
rect 27847 6205 27859 6208
rect 27801 6199 27859 6205
rect 27982 6196 27988 6208
rect 28040 6196 28046 6248
rect 28537 6239 28595 6245
rect 28537 6205 28549 6239
rect 28583 6205 28595 6239
rect 28537 6199 28595 6205
rect 24452 6140 25544 6168
rect 24452 6128 24458 6140
rect 26786 6128 26792 6180
rect 26844 6168 26850 6180
rect 28166 6168 28172 6180
rect 26844 6140 28172 6168
rect 26844 6128 26850 6140
rect 28166 6128 28172 6140
rect 28224 6168 28230 6180
rect 28552 6168 28580 6199
rect 28224 6140 28580 6168
rect 31496 6168 31524 6267
rect 31680 6236 31708 6267
rect 31938 6236 31944 6248
rect 31680 6208 31944 6236
rect 31938 6196 31944 6208
rect 31996 6196 32002 6248
rect 32140 6236 32168 6276
rect 32214 6264 32220 6316
rect 32272 6304 32278 6316
rect 33042 6304 33048 6316
rect 32272 6276 33048 6304
rect 32272 6264 32278 6276
rect 33042 6264 33048 6276
rect 33100 6264 33106 6316
rect 33134 6264 33140 6316
rect 33192 6264 33198 6316
rect 33229 6307 33287 6313
rect 33229 6273 33241 6307
rect 33275 6273 33287 6307
rect 33229 6267 33287 6273
rect 33244 6236 33272 6267
rect 33410 6264 33416 6316
rect 33468 6264 33474 6316
rect 34054 6264 34060 6316
rect 34112 6264 34118 6316
rect 34149 6307 34207 6313
rect 34149 6273 34161 6307
rect 34195 6273 34207 6307
rect 34149 6267 34207 6273
rect 33873 6239 33931 6245
rect 33873 6236 33885 6239
rect 32140 6208 33180 6236
rect 33244 6208 33885 6236
rect 32858 6168 32864 6180
rect 31496 6140 32864 6168
rect 28224 6128 28230 6140
rect 32858 6128 32864 6140
rect 32916 6128 32922 6180
rect 33152 6168 33180 6208
rect 33873 6205 33885 6208
rect 33919 6205 33931 6239
rect 33873 6199 33931 6205
rect 33962 6196 33968 6248
rect 34020 6236 34026 6248
rect 34164 6236 34192 6267
rect 34238 6264 34244 6316
rect 34296 6304 34302 6316
rect 34425 6307 34483 6313
rect 34425 6304 34437 6307
rect 34296 6276 34437 6304
rect 34296 6264 34302 6276
rect 34425 6273 34437 6276
rect 34471 6273 34483 6307
rect 34425 6267 34483 6273
rect 34020 6208 34192 6236
rect 34020 6196 34026 6208
rect 34330 6196 34336 6248
rect 34388 6196 34394 6248
rect 34440 6236 34468 6267
rect 34974 6264 34980 6316
rect 35032 6264 35038 6316
rect 35084 6313 35112 6344
rect 35176 6344 36268 6372
rect 35176 6313 35204 6344
rect 36262 6332 36268 6344
rect 36320 6332 36326 6384
rect 38930 6332 38936 6384
rect 38988 6372 38994 6384
rect 38988 6344 39620 6372
rect 38988 6332 38994 6344
rect 35069 6307 35127 6313
rect 35069 6273 35081 6307
rect 35115 6273 35127 6307
rect 35069 6267 35127 6273
rect 35161 6307 35219 6313
rect 35161 6273 35173 6307
rect 35207 6273 35219 6307
rect 35161 6267 35219 6273
rect 35894 6264 35900 6316
rect 35952 6264 35958 6316
rect 36078 6264 36084 6316
rect 36136 6264 36142 6316
rect 38473 6307 38531 6313
rect 38473 6273 38485 6307
rect 38519 6304 38531 6307
rect 38519 6276 39436 6304
rect 38519 6273 38531 6276
rect 38473 6267 38531 6273
rect 38930 6236 38936 6248
rect 34440 6208 38936 6236
rect 38930 6196 38936 6208
rect 38988 6196 38994 6248
rect 39408 6245 39436 6276
rect 39482 6264 39488 6316
rect 39540 6264 39546 6316
rect 39592 6313 39620 6344
rect 40218 6332 40224 6384
rect 40276 6372 40282 6384
rect 40494 6372 40500 6384
rect 40276 6344 40500 6372
rect 40276 6332 40282 6344
rect 40494 6332 40500 6344
rect 40552 6332 40558 6384
rect 42705 6375 42763 6381
rect 42705 6372 42717 6375
rect 41814 6344 42717 6372
rect 42705 6341 42717 6344
rect 42751 6341 42763 6375
rect 42705 6335 42763 6341
rect 39577 6307 39635 6313
rect 39577 6273 39589 6307
rect 39623 6273 39635 6307
rect 39577 6267 39635 6273
rect 40034 6264 40040 6316
rect 40092 6304 40098 6316
rect 40313 6307 40371 6313
rect 40313 6304 40325 6307
rect 40092 6276 40325 6304
rect 40092 6264 40098 6276
rect 40313 6273 40325 6276
rect 40359 6273 40371 6307
rect 40313 6267 40371 6273
rect 42610 6264 42616 6316
rect 42668 6264 42674 6316
rect 39301 6239 39359 6245
rect 39301 6205 39313 6239
rect 39347 6205 39359 6239
rect 39301 6199 39359 6205
rect 39393 6239 39451 6245
rect 39393 6205 39405 6239
rect 39439 6205 39451 6239
rect 39393 6199 39451 6205
rect 33318 6168 33324 6180
rect 33152 6140 33324 6168
rect 33318 6128 33324 6140
rect 33376 6128 33382 6180
rect 34256 6140 36032 6168
rect 19760 6072 23244 6100
rect 19760 6060 19766 6072
rect 26326 6060 26332 6112
rect 26384 6100 26390 6112
rect 27249 6103 27307 6109
rect 27249 6100 27261 6103
rect 26384 6072 27261 6100
rect 26384 6060 26390 6072
rect 27249 6069 27261 6072
rect 27295 6069 27307 6103
rect 27249 6063 27307 6069
rect 29917 6103 29975 6109
rect 29917 6069 29929 6103
rect 29963 6100 29975 6103
rect 30098 6100 30104 6112
rect 29963 6072 30104 6100
rect 29963 6069 29975 6072
rect 29917 6063 29975 6069
rect 30098 6060 30104 6072
rect 30156 6060 30162 6112
rect 32030 6060 32036 6112
rect 32088 6100 32094 6112
rect 32674 6100 32680 6112
rect 32088 6072 32680 6100
rect 32088 6060 32094 6072
rect 32674 6060 32680 6072
rect 32732 6100 32738 6112
rect 34256 6100 34284 6140
rect 36004 6112 36032 6140
rect 32732 6072 34284 6100
rect 32732 6060 32738 6072
rect 35342 6060 35348 6112
rect 35400 6060 35406 6112
rect 35986 6060 35992 6112
rect 36044 6060 36050 6112
rect 39114 6060 39120 6112
rect 39172 6060 39178 6112
rect 39316 6100 39344 6199
rect 39408 6168 39436 6199
rect 40586 6196 40592 6248
rect 40644 6196 40650 6248
rect 39408 6140 40264 6168
rect 40236 6112 40264 6140
rect 40126 6100 40132 6112
rect 39316 6072 40132 6100
rect 40126 6060 40132 6072
rect 40184 6060 40190 6112
rect 40218 6060 40224 6112
rect 40276 6100 40282 6112
rect 42061 6103 42119 6109
rect 42061 6100 42073 6103
rect 40276 6072 42073 6100
rect 40276 6060 40282 6072
rect 42061 6069 42073 6072
rect 42107 6069 42119 6103
rect 42061 6063 42119 6069
rect 1104 6010 44896 6032
rect 1104 5958 6423 6010
rect 6475 5958 6487 6010
rect 6539 5958 6551 6010
rect 6603 5958 6615 6010
rect 6667 5958 6679 6010
rect 6731 5958 17370 6010
rect 17422 5958 17434 6010
rect 17486 5958 17498 6010
rect 17550 5958 17562 6010
rect 17614 5958 17626 6010
rect 17678 5958 28317 6010
rect 28369 5958 28381 6010
rect 28433 5958 28445 6010
rect 28497 5958 28509 6010
rect 28561 5958 28573 6010
rect 28625 5958 39264 6010
rect 39316 5958 39328 6010
rect 39380 5958 39392 6010
rect 39444 5958 39456 6010
rect 39508 5958 39520 6010
rect 39572 5958 44896 6010
rect 1104 5936 44896 5958
rect 3234 5856 3240 5908
rect 3292 5856 3298 5908
rect 5258 5856 5264 5908
rect 5316 5896 5322 5908
rect 5353 5899 5411 5905
rect 5353 5896 5365 5899
rect 5316 5868 5365 5896
rect 5316 5856 5322 5868
rect 5353 5865 5365 5868
rect 5399 5865 5411 5899
rect 5353 5859 5411 5865
rect 9582 5856 9588 5908
rect 9640 5896 9646 5908
rect 11701 5899 11759 5905
rect 11701 5896 11713 5899
rect 9640 5868 11713 5896
rect 9640 5856 9646 5868
rect 11701 5865 11713 5868
rect 11747 5896 11759 5899
rect 12250 5896 12256 5908
rect 11747 5868 12256 5896
rect 11747 5865 11759 5868
rect 11701 5859 11759 5865
rect 12250 5856 12256 5868
rect 12308 5856 12314 5908
rect 12986 5856 12992 5908
rect 13044 5896 13050 5908
rect 13722 5896 13728 5908
rect 13044 5868 13728 5896
rect 13044 5856 13050 5868
rect 13722 5856 13728 5868
rect 13780 5896 13786 5908
rect 14369 5899 14427 5905
rect 14369 5896 14381 5899
rect 13780 5868 14381 5896
rect 13780 5856 13786 5868
rect 14369 5865 14381 5868
rect 14415 5865 14427 5899
rect 14369 5859 14427 5865
rect 14458 5856 14464 5908
rect 14516 5856 14522 5908
rect 15286 5856 15292 5908
rect 15344 5896 15350 5908
rect 18233 5899 18291 5905
rect 15344 5868 18184 5896
rect 15344 5856 15350 5868
rect 12526 5788 12532 5840
rect 12584 5828 12590 5840
rect 14182 5828 14188 5840
rect 12584 5800 14188 5828
rect 12584 5788 12590 5800
rect 14182 5788 14188 5800
rect 14240 5788 14246 5840
rect 3970 5720 3976 5772
rect 4028 5720 4034 5772
rect 5810 5720 5816 5772
rect 5868 5760 5874 5772
rect 5868 5732 9628 5760
rect 5868 5720 5874 5732
rect 9600 5704 9628 5732
rect 13354 5720 13360 5772
rect 13412 5760 13418 5772
rect 14553 5763 14611 5769
rect 14553 5760 14565 5763
rect 13412 5732 14565 5760
rect 13412 5720 13418 5732
rect 14553 5729 14565 5732
rect 14599 5760 14611 5763
rect 14642 5760 14648 5772
rect 14599 5732 14648 5760
rect 14599 5729 14611 5732
rect 14553 5723 14611 5729
rect 14642 5720 14648 5732
rect 14700 5720 14706 5772
rect 16485 5763 16543 5769
rect 16485 5729 16497 5763
rect 16531 5760 16543 5763
rect 17126 5760 17132 5772
rect 16531 5732 17132 5760
rect 16531 5729 16543 5732
rect 16485 5723 16543 5729
rect 17126 5720 17132 5732
rect 17184 5720 17190 5772
rect 18156 5760 18184 5868
rect 18233 5865 18245 5899
rect 18279 5896 18291 5899
rect 18414 5896 18420 5908
rect 18279 5868 18420 5896
rect 18279 5865 18291 5868
rect 18233 5859 18291 5865
rect 18414 5856 18420 5868
rect 18472 5856 18478 5908
rect 20898 5856 20904 5908
rect 20956 5896 20962 5908
rect 21542 5896 21548 5908
rect 20956 5868 21548 5896
rect 20956 5856 20962 5868
rect 18322 5788 18328 5840
rect 18380 5828 18386 5840
rect 19150 5828 19156 5840
rect 18380 5800 19156 5828
rect 18380 5788 18386 5800
rect 19150 5788 19156 5800
rect 19208 5828 19214 5840
rect 19208 5800 20576 5828
rect 19208 5788 19214 5800
rect 18156 5732 18828 5760
rect 2130 5652 2136 5704
rect 2188 5692 2194 5704
rect 2777 5695 2835 5701
rect 2777 5692 2789 5695
rect 2188 5664 2789 5692
rect 2188 5652 2194 5664
rect 2777 5661 2789 5664
rect 2823 5661 2835 5695
rect 2777 5655 2835 5661
rect 3421 5695 3479 5701
rect 3421 5661 3433 5695
rect 3467 5692 3479 5695
rect 5166 5692 5172 5704
rect 3467 5664 5172 5692
rect 3467 5661 3479 5664
rect 3421 5655 3479 5661
rect 5166 5652 5172 5664
rect 5224 5652 5230 5704
rect 5994 5652 6000 5704
rect 6052 5652 6058 5704
rect 9582 5652 9588 5704
rect 9640 5652 9646 5704
rect 9769 5695 9827 5701
rect 9769 5661 9781 5695
rect 9815 5692 9827 5695
rect 10042 5692 10048 5704
rect 9815 5664 10048 5692
rect 9815 5661 9827 5664
rect 9769 5655 9827 5661
rect 10042 5652 10048 5664
rect 10100 5652 10106 5704
rect 10410 5652 10416 5704
rect 10468 5652 10474 5704
rect 13170 5652 13176 5704
rect 13228 5692 13234 5704
rect 14277 5695 14335 5701
rect 14277 5692 14289 5695
rect 13228 5664 14289 5692
rect 13228 5652 13234 5664
rect 14277 5661 14289 5664
rect 14323 5692 14335 5695
rect 14826 5692 14832 5704
rect 14323 5664 14832 5692
rect 14323 5661 14335 5664
rect 14277 5655 14335 5661
rect 14826 5652 14832 5664
rect 14884 5652 14890 5704
rect 16022 5652 16028 5704
rect 16080 5652 16086 5704
rect 18690 5652 18696 5704
rect 18748 5652 18754 5704
rect 18800 5692 18828 5732
rect 20346 5720 20352 5772
rect 20404 5720 20410 5772
rect 20548 5760 20576 5800
rect 21284 5769 21312 5868
rect 21542 5856 21548 5868
rect 21600 5856 21606 5908
rect 21910 5856 21916 5908
rect 21968 5896 21974 5908
rect 24394 5896 24400 5908
rect 21968 5868 24400 5896
rect 21968 5856 21974 5868
rect 24394 5856 24400 5868
rect 24452 5856 24458 5908
rect 29730 5856 29736 5908
rect 29788 5856 29794 5908
rect 31938 5856 31944 5908
rect 31996 5896 32002 5908
rect 32490 5896 32496 5908
rect 31996 5868 32496 5896
rect 31996 5856 32002 5868
rect 32490 5856 32496 5868
rect 32548 5856 32554 5908
rect 32677 5899 32735 5905
rect 32677 5865 32689 5899
rect 32723 5896 32735 5899
rect 33410 5896 33416 5908
rect 32723 5868 33416 5896
rect 32723 5865 32735 5868
rect 32677 5859 32735 5865
rect 33410 5856 33416 5868
rect 33468 5856 33474 5908
rect 34057 5899 34115 5905
rect 34057 5865 34069 5899
rect 34103 5896 34115 5899
rect 34146 5896 34152 5908
rect 34103 5868 34152 5896
rect 34103 5865 34115 5868
rect 34057 5859 34115 5865
rect 34146 5856 34152 5868
rect 34204 5856 34210 5908
rect 34422 5856 34428 5908
rect 34480 5896 34486 5908
rect 34977 5899 35035 5905
rect 34977 5896 34989 5899
rect 34480 5868 34989 5896
rect 34480 5856 34486 5868
rect 34977 5865 34989 5868
rect 35023 5865 35035 5899
rect 34977 5859 35035 5865
rect 35894 5856 35900 5908
rect 35952 5896 35958 5908
rect 39666 5896 39672 5908
rect 35952 5868 39672 5896
rect 35952 5856 35958 5868
rect 27890 5788 27896 5840
rect 27948 5828 27954 5840
rect 28169 5831 28227 5837
rect 28169 5828 28181 5831
rect 27948 5800 28181 5828
rect 27948 5788 27954 5800
rect 28169 5797 28181 5800
rect 28215 5828 28227 5831
rect 33594 5828 33600 5840
rect 28215 5800 33600 5828
rect 28215 5797 28227 5800
rect 28169 5791 28227 5797
rect 21269 5763 21327 5769
rect 20548 5732 21128 5760
rect 18800 5664 20024 5692
rect 4218 5627 4276 5633
rect 4218 5624 4230 5627
rect 2608 5596 4230 5624
rect 2608 5565 2636 5596
rect 4218 5593 4230 5596
rect 4264 5593 4276 5627
rect 4218 5587 4276 5593
rect 16758 5584 16764 5636
rect 16816 5584 16822 5636
rect 18785 5627 18843 5633
rect 18785 5624 18797 5627
rect 17986 5596 18797 5624
rect 18785 5593 18797 5596
rect 18831 5593 18843 5627
rect 19996 5624 20024 5664
rect 20364 5688 20392 5720
rect 20441 5695 20499 5701
rect 20441 5688 20453 5695
rect 20364 5661 20453 5688
rect 20487 5661 20499 5695
rect 20364 5660 20499 5661
rect 20441 5655 20499 5660
rect 20530 5652 20536 5704
rect 20588 5652 20594 5704
rect 20622 5652 20628 5704
rect 20680 5652 20686 5704
rect 20809 5695 20867 5701
rect 20809 5661 20821 5695
rect 20855 5692 20867 5695
rect 20990 5692 20996 5704
rect 20855 5664 20996 5692
rect 20855 5661 20867 5664
rect 20809 5655 20867 5661
rect 20990 5652 20996 5664
rect 21048 5652 21054 5704
rect 21100 5692 21128 5732
rect 21269 5729 21281 5763
rect 21315 5729 21327 5763
rect 21269 5723 21327 5729
rect 24578 5720 24584 5772
rect 24636 5760 24642 5772
rect 26786 5760 26792 5772
rect 24636 5732 26792 5760
rect 24636 5720 24642 5732
rect 26786 5720 26792 5732
rect 26844 5720 26850 5772
rect 27982 5720 27988 5772
rect 28040 5760 28046 5772
rect 30285 5763 30343 5769
rect 30285 5760 30297 5763
rect 28040 5732 30297 5760
rect 28040 5720 28046 5732
rect 30285 5729 30297 5732
rect 30331 5760 30343 5763
rect 30466 5760 30472 5772
rect 30331 5732 30472 5760
rect 30331 5729 30343 5732
rect 30285 5723 30343 5729
rect 30466 5720 30472 5732
rect 30524 5720 30530 5772
rect 33336 5769 33364 5800
rect 33594 5788 33600 5800
rect 33652 5788 33658 5840
rect 33686 5788 33692 5840
rect 33744 5788 33750 5840
rect 35621 5831 35679 5837
rect 35621 5828 35633 5831
rect 34072 5800 35633 5828
rect 33321 5763 33379 5769
rect 30576 5732 33180 5760
rect 21910 5692 21916 5704
rect 21100 5664 21916 5692
rect 21910 5652 21916 5664
rect 21968 5652 21974 5704
rect 26326 5652 26332 5704
rect 26384 5652 26390 5704
rect 27430 5652 27436 5704
rect 27488 5692 27494 5704
rect 28813 5695 28871 5701
rect 28813 5692 28825 5695
rect 27488 5664 28825 5692
rect 27488 5652 27494 5664
rect 28813 5661 28825 5664
rect 28859 5661 28871 5695
rect 28813 5655 28871 5661
rect 30098 5652 30104 5704
rect 30156 5692 30162 5704
rect 30576 5692 30604 5732
rect 30156 5664 30604 5692
rect 31389 5695 31447 5701
rect 30156 5652 30162 5664
rect 31389 5661 31401 5695
rect 31435 5692 31447 5695
rect 31938 5692 31944 5704
rect 31435 5664 31944 5692
rect 31435 5661 31447 5664
rect 31389 5655 31447 5661
rect 31938 5652 31944 5664
rect 31996 5652 32002 5704
rect 32030 5652 32036 5704
rect 32088 5652 32094 5704
rect 32214 5652 32220 5704
rect 32272 5652 32278 5704
rect 32858 5695 32916 5701
rect 32858 5661 32870 5695
rect 32904 5692 32916 5695
rect 32950 5692 32956 5704
rect 32904 5664 32956 5692
rect 32904 5661 32916 5664
rect 32858 5655 32916 5661
rect 32950 5652 32956 5664
rect 33008 5652 33014 5704
rect 20165 5627 20223 5633
rect 19996 5596 20116 5624
rect 18785 5587 18843 5593
rect 2593 5559 2651 5565
rect 2593 5525 2605 5559
rect 2639 5525 2651 5559
rect 2593 5519 2651 5525
rect 6181 5559 6239 5565
rect 6181 5525 6193 5559
rect 6227 5556 6239 5559
rect 7742 5556 7748 5568
rect 6227 5528 7748 5556
rect 6227 5525 6239 5528
rect 6181 5519 6239 5525
rect 7742 5516 7748 5528
rect 7800 5516 7806 5568
rect 9950 5516 9956 5568
rect 10008 5516 10014 5568
rect 15841 5559 15899 5565
rect 15841 5525 15853 5559
rect 15887 5556 15899 5559
rect 16574 5556 16580 5568
rect 15887 5528 16580 5556
rect 15887 5525 15899 5528
rect 15841 5519 15899 5525
rect 16574 5516 16580 5528
rect 16632 5516 16638 5568
rect 20088 5556 20116 5596
rect 20165 5593 20177 5627
rect 20211 5624 20223 5627
rect 21514 5627 21572 5633
rect 21514 5624 21526 5627
rect 20211 5596 21526 5624
rect 20211 5593 20223 5596
rect 20165 5587 20223 5593
rect 21514 5593 21526 5596
rect 21560 5593 21572 5627
rect 27034 5627 27092 5633
rect 27034 5624 27046 5627
rect 21514 5587 21572 5593
rect 26160 5596 27046 5624
rect 20438 5556 20444 5568
rect 20088 5528 20444 5556
rect 20438 5516 20444 5528
rect 20496 5556 20502 5568
rect 20990 5556 20996 5568
rect 20496 5528 20996 5556
rect 20496 5516 20502 5528
rect 20990 5516 20996 5528
rect 21048 5516 21054 5568
rect 21174 5516 21180 5568
rect 21232 5556 21238 5568
rect 26160 5565 26188 5596
rect 27034 5593 27046 5596
rect 27080 5593 27092 5627
rect 27034 5587 27092 5593
rect 30190 5584 30196 5636
rect 30248 5584 30254 5636
rect 31481 5627 31539 5633
rect 31481 5593 31493 5627
rect 31527 5624 31539 5627
rect 33152 5624 33180 5732
rect 33321 5729 33333 5763
rect 33367 5729 33379 5763
rect 33704 5760 33732 5788
rect 34072 5760 34100 5800
rect 35621 5797 35633 5800
rect 35667 5797 35679 5831
rect 35621 5791 35679 5797
rect 33321 5723 33379 5729
rect 33612 5732 34100 5760
rect 34149 5763 34207 5769
rect 33229 5695 33287 5701
rect 33229 5661 33241 5695
rect 33275 5692 33287 5695
rect 33612 5692 33640 5732
rect 34149 5729 34161 5763
rect 34195 5760 34207 5763
rect 35342 5760 35348 5772
rect 34195 5732 35348 5760
rect 34195 5729 34207 5732
rect 34149 5723 34207 5729
rect 35342 5720 35348 5732
rect 35400 5720 35406 5772
rect 33275 5664 33640 5692
rect 33275 5661 33287 5664
rect 33229 5655 33287 5661
rect 33686 5652 33692 5704
rect 33744 5692 33750 5704
rect 34885 5695 34943 5701
rect 34885 5692 34897 5695
rect 33744 5664 34897 5692
rect 33744 5652 33750 5664
rect 34885 5661 34897 5664
rect 34931 5661 34943 5695
rect 34885 5655 34943 5661
rect 35529 5695 35587 5701
rect 35529 5661 35541 5695
rect 35575 5661 35587 5695
rect 35529 5655 35587 5661
rect 33781 5627 33839 5633
rect 33781 5624 33793 5627
rect 31527 5596 33088 5624
rect 33152 5596 33793 5624
rect 31527 5593 31539 5596
rect 31481 5587 31539 5593
rect 22649 5559 22707 5565
rect 22649 5556 22661 5559
rect 21232 5528 22661 5556
rect 21232 5516 21238 5528
rect 22649 5525 22661 5528
rect 22695 5525 22707 5559
rect 22649 5519 22707 5525
rect 26145 5559 26203 5565
rect 26145 5525 26157 5559
rect 26191 5525 26203 5559
rect 26145 5519 26203 5525
rect 28258 5516 28264 5568
rect 28316 5556 28322 5568
rect 28629 5559 28687 5565
rect 28629 5556 28641 5559
rect 28316 5528 28641 5556
rect 28316 5516 28322 5528
rect 28629 5525 28641 5528
rect 28675 5525 28687 5559
rect 28629 5519 28687 5525
rect 32122 5516 32128 5568
rect 32180 5516 32186 5568
rect 32766 5516 32772 5568
rect 32824 5556 32830 5568
rect 32861 5559 32919 5565
rect 32861 5556 32873 5559
rect 32824 5528 32873 5556
rect 32824 5516 32830 5528
rect 32861 5525 32873 5528
rect 32907 5525 32919 5559
rect 33060 5556 33088 5596
rect 33781 5593 33793 5596
rect 33827 5624 33839 5627
rect 34054 5624 34060 5636
rect 33827 5596 34060 5624
rect 33827 5593 33839 5596
rect 33781 5587 33839 5593
rect 34054 5584 34060 5596
rect 34112 5584 34118 5636
rect 34146 5584 34152 5636
rect 34204 5624 34210 5636
rect 34241 5627 34299 5633
rect 34241 5624 34253 5627
rect 34204 5596 34253 5624
rect 34204 5584 34210 5596
rect 34241 5593 34253 5596
rect 34287 5593 34299 5627
rect 34241 5587 34299 5593
rect 33873 5559 33931 5565
rect 33873 5556 33885 5559
rect 33060 5528 33885 5556
rect 32861 5519 32919 5525
rect 33873 5525 33885 5528
rect 33919 5556 33931 5559
rect 33962 5556 33968 5568
rect 33919 5528 33968 5556
rect 33919 5525 33931 5528
rect 33873 5519 33931 5525
rect 33962 5516 33968 5528
rect 34020 5516 34026 5568
rect 35544 5556 35572 5655
rect 36556 5633 36584 5868
rect 39666 5856 39672 5868
rect 39724 5856 39730 5908
rect 40126 5856 40132 5908
rect 40184 5896 40190 5908
rect 40402 5896 40408 5908
rect 40184 5868 40408 5896
rect 40184 5856 40190 5868
rect 40402 5856 40408 5868
rect 40460 5856 40466 5908
rect 40494 5856 40500 5908
rect 40552 5896 40558 5908
rect 40862 5896 40868 5908
rect 40552 5868 40868 5896
rect 40552 5856 40558 5868
rect 40862 5856 40868 5868
rect 40920 5896 40926 5908
rect 42613 5899 42671 5905
rect 42613 5896 42625 5899
rect 40920 5868 42625 5896
rect 40920 5856 40926 5868
rect 42613 5865 42625 5868
rect 42659 5865 42671 5899
rect 42613 5859 42671 5865
rect 39022 5788 39028 5840
rect 39080 5828 39086 5840
rect 39485 5831 39543 5837
rect 39485 5828 39497 5831
rect 39080 5800 39497 5828
rect 39080 5788 39086 5800
rect 39485 5797 39497 5800
rect 39531 5797 39543 5831
rect 39485 5791 39543 5797
rect 40034 5788 40040 5840
rect 40092 5828 40098 5840
rect 40092 5800 40908 5828
rect 40092 5788 40098 5800
rect 37458 5720 37464 5772
rect 37516 5760 37522 5772
rect 37737 5763 37795 5769
rect 37737 5760 37749 5763
rect 37516 5732 37749 5760
rect 37516 5720 37522 5732
rect 37737 5729 37749 5732
rect 37783 5729 37795 5763
rect 40218 5760 40224 5772
rect 37737 5723 37795 5729
rect 40052 5732 40224 5760
rect 40052 5701 40080 5732
rect 40218 5720 40224 5732
rect 40276 5720 40282 5772
rect 40310 5720 40316 5772
rect 40368 5720 40374 5772
rect 40880 5769 40908 5800
rect 40865 5763 40923 5769
rect 40865 5729 40877 5763
rect 40911 5729 40923 5763
rect 40865 5723 40923 5729
rect 40037 5695 40095 5701
rect 40037 5661 40049 5695
rect 40083 5661 40095 5695
rect 40037 5655 40095 5661
rect 40126 5652 40132 5704
rect 40184 5692 40190 5704
rect 40328 5692 40356 5720
rect 40184 5664 40356 5692
rect 40184 5652 40190 5664
rect 42242 5652 42248 5704
rect 42300 5652 42306 5704
rect 44082 5652 44088 5704
rect 44140 5652 44146 5704
rect 36541 5627 36599 5633
rect 36541 5593 36553 5627
rect 36587 5593 36599 5627
rect 36541 5587 36599 5593
rect 36725 5627 36783 5633
rect 36725 5593 36737 5627
rect 36771 5624 36783 5627
rect 37182 5624 37188 5636
rect 36771 5596 37188 5624
rect 36771 5593 36783 5596
rect 36725 5587 36783 5593
rect 36078 5556 36084 5568
rect 35544 5528 36084 5556
rect 36078 5516 36084 5528
rect 36136 5556 36142 5568
rect 36740 5556 36768 5587
rect 37182 5584 37188 5596
rect 37240 5584 37246 5636
rect 38010 5584 38016 5636
rect 38068 5584 38074 5636
rect 38654 5584 38660 5636
rect 38712 5584 38718 5636
rect 41138 5584 41144 5636
rect 41196 5584 41202 5636
rect 36136 5528 36768 5556
rect 36136 5516 36142 5528
rect 36906 5516 36912 5568
rect 36964 5516 36970 5568
rect 40313 5559 40371 5565
rect 40313 5525 40325 5559
rect 40359 5556 40371 5559
rect 41046 5556 41052 5568
rect 40359 5528 41052 5556
rect 40359 5525 40371 5528
rect 40313 5519 40371 5525
rect 41046 5516 41052 5528
rect 41104 5516 41110 5568
rect 44269 5559 44327 5565
rect 44269 5525 44281 5559
rect 44315 5556 44327 5559
rect 45002 5556 45008 5568
rect 44315 5528 45008 5556
rect 44315 5525 44327 5528
rect 44269 5519 44327 5525
rect 45002 5516 45008 5528
rect 45060 5516 45066 5568
rect 1104 5466 45051 5488
rect 1104 5414 11896 5466
rect 11948 5414 11960 5466
rect 12012 5414 12024 5466
rect 12076 5414 12088 5466
rect 12140 5414 12152 5466
rect 12204 5414 22843 5466
rect 22895 5414 22907 5466
rect 22959 5414 22971 5466
rect 23023 5414 23035 5466
rect 23087 5414 23099 5466
rect 23151 5414 33790 5466
rect 33842 5414 33854 5466
rect 33906 5414 33918 5466
rect 33970 5414 33982 5466
rect 34034 5414 34046 5466
rect 34098 5414 44737 5466
rect 44789 5414 44801 5466
rect 44853 5414 44865 5466
rect 44917 5414 44929 5466
rect 44981 5414 44993 5466
rect 45045 5414 45051 5466
rect 1104 5392 45051 5414
rect 5350 5312 5356 5364
rect 5408 5312 5414 5364
rect 13633 5355 13691 5361
rect 13633 5321 13645 5355
rect 13679 5352 13691 5355
rect 14090 5352 14096 5364
rect 13679 5324 14096 5352
rect 13679 5321 13691 5324
rect 13633 5315 13691 5321
rect 14090 5312 14096 5324
rect 14148 5312 14154 5364
rect 15470 5312 15476 5364
rect 15528 5352 15534 5364
rect 15528 5324 18552 5352
rect 15528 5312 15534 5324
rect 9582 5284 9588 5296
rect 9232 5256 9588 5284
rect 3970 5176 3976 5228
rect 4028 5176 4034 5228
rect 4246 5225 4252 5228
rect 4240 5216 4252 5225
rect 4080 5188 4252 5216
rect 934 5108 940 5160
rect 992 5148 998 5160
rect 1581 5151 1639 5157
rect 1581 5148 1593 5151
rect 992 5120 1593 5148
rect 992 5108 998 5120
rect 1581 5117 1593 5120
rect 1627 5117 1639 5151
rect 1581 5111 1639 5117
rect 1857 5151 1915 5157
rect 1857 5117 1869 5151
rect 1903 5148 1915 5151
rect 4080 5148 4108 5188
rect 4240 5179 4252 5188
rect 4246 5176 4252 5179
rect 4304 5176 4310 5228
rect 9232 5225 9260 5256
rect 9582 5244 9588 5256
rect 9640 5284 9646 5296
rect 9640 5256 14780 5284
rect 9640 5244 9646 5256
rect 14752 5228 14780 5256
rect 9217 5219 9275 5225
rect 9217 5185 9229 5219
rect 9263 5185 9275 5219
rect 9217 5179 9275 5185
rect 9306 5176 9312 5228
rect 9364 5216 9370 5228
rect 9401 5219 9459 5225
rect 9401 5216 9413 5219
rect 9364 5188 9413 5216
rect 9364 5176 9370 5188
rect 9401 5185 9413 5188
rect 9447 5185 9459 5219
rect 9401 5179 9459 5185
rect 12250 5176 12256 5228
rect 12308 5176 12314 5228
rect 12520 5219 12578 5225
rect 12520 5185 12532 5219
rect 12566 5216 12578 5219
rect 13078 5216 13084 5228
rect 12566 5188 13084 5216
rect 12566 5185 12578 5188
rect 12520 5179 12578 5185
rect 13078 5176 13084 5188
rect 13136 5176 13142 5228
rect 14090 5176 14096 5228
rect 14148 5176 14154 5228
rect 14734 5176 14740 5228
rect 14792 5216 14798 5228
rect 15488 5225 15516 5312
rect 17126 5284 17132 5296
rect 16868 5256 17132 5284
rect 16868 5225 16896 5256
rect 17126 5244 17132 5256
rect 17184 5244 17190 5296
rect 18414 5284 18420 5296
rect 18354 5256 18420 5284
rect 18414 5244 18420 5256
rect 18472 5244 18478 5296
rect 18524 5284 18552 5324
rect 18598 5312 18604 5364
rect 18656 5312 18662 5364
rect 21085 5355 21143 5361
rect 21085 5321 21097 5355
rect 21131 5352 21143 5355
rect 21818 5352 21824 5364
rect 21131 5324 21824 5352
rect 21131 5321 21143 5324
rect 21085 5315 21143 5321
rect 21818 5312 21824 5324
rect 21876 5312 21882 5364
rect 24394 5312 24400 5364
rect 24452 5312 24458 5364
rect 28166 5312 28172 5364
rect 28224 5352 28230 5364
rect 29917 5355 29975 5361
rect 29917 5352 29929 5355
rect 28224 5324 29929 5352
rect 28224 5312 28230 5324
rect 29917 5321 29929 5324
rect 29963 5352 29975 5355
rect 31202 5352 31208 5364
rect 29963 5324 31208 5352
rect 29963 5321 29975 5324
rect 29917 5315 29975 5321
rect 31202 5312 31208 5324
rect 31260 5312 31266 5364
rect 32858 5312 32864 5364
rect 32916 5352 32922 5364
rect 34146 5352 34152 5364
rect 32916 5324 34152 5352
rect 32916 5312 32922 5324
rect 34146 5312 34152 5324
rect 34204 5312 34210 5364
rect 34606 5312 34612 5364
rect 34664 5352 34670 5364
rect 35069 5355 35127 5361
rect 35069 5352 35081 5355
rect 34664 5324 35081 5352
rect 34664 5312 34670 5324
rect 35069 5321 35081 5324
rect 35115 5352 35127 5355
rect 35434 5352 35440 5364
rect 35115 5324 35440 5352
rect 35115 5321 35127 5324
rect 35069 5315 35127 5321
rect 35434 5312 35440 5324
rect 35492 5312 35498 5364
rect 36199 5355 36257 5361
rect 36199 5321 36211 5355
rect 36245 5352 36257 5355
rect 36906 5352 36912 5364
rect 36245 5324 36912 5352
rect 36245 5321 36257 5324
rect 36199 5315 36257 5321
rect 36906 5312 36912 5324
rect 36964 5312 36970 5364
rect 38683 5355 38741 5361
rect 38683 5321 38695 5355
rect 38729 5352 38741 5355
rect 39114 5352 39120 5364
rect 38729 5324 39120 5352
rect 38729 5321 38741 5324
rect 38683 5315 38741 5321
rect 39114 5312 39120 5324
rect 39172 5312 39178 5364
rect 40494 5312 40500 5364
rect 40552 5312 40558 5364
rect 40586 5312 40592 5364
rect 40644 5352 40650 5364
rect 41141 5355 41199 5361
rect 41141 5352 41153 5355
rect 40644 5324 41153 5352
rect 40644 5312 40650 5324
rect 41141 5321 41153 5324
rect 41187 5321 41199 5355
rect 41141 5315 41199 5321
rect 24578 5284 24584 5296
rect 18524 5256 22094 5284
rect 15289 5219 15347 5225
rect 15289 5216 15301 5219
rect 14792 5188 15301 5216
rect 14792 5176 14798 5188
rect 15289 5185 15301 5188
rect 15335 5185 15347 5219
rect 15289 5179 15347 5185
rect 15473 5219 15531 5225
rect 15473 5185 15485 5219
rect 15519 5185 15531 5219
rect 15473 5179 15531 5185
rect 16853 5219 16911 5225
rect 16853 5185 16865 5219
rect 16899 5185 16911 5219
rect 16853 5179 16911 5185
rect 19242 5176 19248 5228
rect 19300 5176 19306 5228
rect 20990 5176 20996 5228
rect 21048 5176 21054 5228
rect 21174 5176 21180 5228
rect 21232 5176 21238 5228
rect 1903 5120 4108 5148
rect 1903 5117 1915 5120
rect 1857 5111 1915 5117
rect 14182 5108 14188 5160
rect 14240 5108 14246 5160
rect 14369 5151 14427 5157
rect 14369 5117 14381 5151
rect 14415 5148 14427 5151
rect 14642 5148 14648 5160
rect 14415 5120 14648 5148
rect 14415 5117 14427 5120
rect 14369 5111 14427 5117
rect 14642 5108 14648 5120
rect 14700 5108 14706 5160
rect 17129 5151 17187 5157
rect 17129 5117 17141 5151
rect 17175 5148 17187 5151
rect 17175 5120 19104 5148
rect 17175 5117 17187 5120
rect 17129 5111 17187 5117
rect 19076 5089 19104 5120
rect 19061 5083 19119 5089
rect 19061 5049 19073 5083
rect 19107 5049 19119 5083
rect 19061 5043 19119 5049
rect 9585 5015 9643 5021
rect 9585 4981 9597 5015
rect 9631 5012 9643 5015
rect 13538 5012 13544 5024
rect 9631 4984 13544 5012
rect 9631 4981 9643 4984
rect 9585 4975 9643 4981
rect 13538 4972 13544 4984
rect 13596 4972 13602 5024
rect 14274 4972 14280 5024
rect 14332 4972 14338 5024
rect 15194 4972 15200 5024
rect 15252 5012 15258 5024
rect 15657 5015 15715 5021
rect 15657 5012 15669 5015
rect 15252 4984 15669 5012
rect 15252 4972 15258 4984
rect 15657 4981 15669 4984
rect 15703 4981 15715 5015
rect 22066 5012 22094 5256
rect 23032 5256 24584 5284
rect 23032 5225 23060 5256
rect 24578 5244 24584 5256
rect 24636 5244 24642 5296
rect 28629 5287 28687 5293
rect 28629 5253 28641 5287
rect 28675 5284 28687 5287
rect 28718 5284 28724 5296
rect 28675 5256 28724 5284
rect 28675 5253 28687 5256
rect 28629 5247 28687 5253
rect 28718 5244 28724 5256
rect 28776 5284 28782 5296
rect 33781 5287 33839 5293
rect 33781 5284 33793 5287
rect 28776 5256 33793 5284
rect 28776 5244 28782 5256
rect 33781 5253 33793 5256
rect 33827 5253 33839 5287
rect 33781 5247 33839 5253
rect 35989 5287 36047 5293
rect 35989 5253 36001 5287
rect 36035 5253 36047 5287
rect 38473 5287 38531 5293
rect 38473 5284 38485 5287
rect 35989 5247 36047 5253
rect 36280 5256 38485 5284
rect 23290 5225 23296 5228
rect 23017 5219 23075 5225
rect 23017 5185 23029 5219
rect 23063 5185 23075 5219
rect 23017 5179 23075 5185
rect 23284 5179 23296 5225
rect 23290 5176 23296 5179
rect 23348 5176 23354 5228
rect 32122 5176 32128 5228
rect 32180 5216 32186 5228
rect 32401 5219 32459 5225
rect 32401 5216 32413 5219
rect 32180 5188 32413 5216
rect 32180 5176 32186 5188
rect 32401 5185 32413 5188
rect 32447 5185 32459 5219
rect 32401 5179 32459 5185
rect 32493 5219 32551 5225
rect 32493 5185 32505 5219
rect 32539 5185 32551 5219
rect 32493 5179 32551 5185
rect 32214 5108 32220 5160
rect 32272 5148 32278 5160
rect 32508 5148 32536 5179
rect 32674 5176 32680 5228
rect 32732 5176 32738 5228
rect 32769 5219 32827 5225
rect 32769 5185 32781 5219
rect 32815 5185 32827 5219
rect 32769 5179 32827 5185
rect 32272 5120 32536 5148
rect 32272 5108 32278 5120
rect 32490 5040 32496 5092
rect 32548 5080 32554 5092
rect 32784 5080 32812 5179
rect 32858 5176 32864 5228
rect 32916 5176 32922 5228
rect 33318 5176 33324 5228
rect 33376 5216 33382 5228
rect 36004 5216 36032 5247
rect 36280 5228 36308 5256
rect 38473 5253 38485 5256
rect 38519 5284 38531 5287
rect 40126 5284 40132 5296
rect 38519 5256 40132 5284
rect 38519 5253 38531 5256
rect 38473 5247 38531 5253
rect 40126 5244 40132 5256
rect 40184 5244 40190 5296
rect 40313 5287 40371 5293
rect 40313 5253 40325 5287
rect 40359 5284 40371 5287
rect 40678 5284 40684 5296
rect 40359 5256 40684 5284
rect 40359 5253 40371 5256
rect 40313 5247 40371 5253
rect 40678 5244 40684 5256
rect 40736 5244 40742 5296
rect 40788 5256 41276 5284
rect 40788 5228 40816 5256
rect 36262 5216 36268 5228
rect 33376 5188 36268 5216
rect 33376 5176 33382 5188
rect 36262 5176 36268 5188
rect 36320 5176 36326 5228
rect 37366 5176 37372 5228
rect 37424 5216 37430 5228
rect 37829 5219 37887 5225
rect 37829 5216 37841 5219
rect 37424 5188 37841 5216
rect 37424 5176 37430 5188
rect 37829 5185 37841 5188
rect 37875 5185 37887 5219
rect 37829 5179 37887 5185
rect 37921 5219 37979 5225
rect 37921 5185 37933 5219
rect 37967 5216 37979 5219
rect 38654 5216 38660 5228
rect 37967 5188 38660 5216
rect 37967 5185 37979 5188
rect 37921 5179 37979 5185
rect 38654 5176 38660 5188
rect 38712 5176 38718 5228
rect 39485 5219 39543 5225
rect 39485 5185 39497 5219
rect 39531 5216 39543 5219
rect 39666 5216 39672 5228
rect 39531 5188 39672 5216
rect 39531 5185 39543 5188
rect 39485 5179 39543 5185
rect 39666 5176 39672 5188
rect 39724 5176 39730 5228
rect 40589 5219 40647 5225
rect 40589 5185 40601 5219
rect 40635 5216 40647 5219
rect 40770 5216 40776 5228
rect 40635 5188 40776 5216
rect 40635 5185 40647 5188
rect 40589 5179 40647 5185
rect 40770 5176 40776 5188
rect 40828 5176 40834 5228
rect 41046 5176 41052 5228
rect 41104 5176 41110 5228
rect 41248 5225 41276 5256
rect 41233 5219 41291 5225
rect 41233 5185 41245 5219
rect 41279 5185 41291 5219
rect 41233 5179 41291 5185
rect 42978 5176 42984 5228
rect 43036 5176 43042 5228
rect 32548 5052 32812 5080
rect 32548 5040 32554 5052
rect 35894 5040 35900 5092
rect 35952 5080 35958 5092
rect 36357 5083 36415 5089
rect 36357 5080 36369 5083
rect 35952 5052 36369 5080
rect 35952 5040 35958 5052
rect 36357 5049 36369 5052
rect 36403 5049 36415 5083
rect 39301 5083 39359 5089
rect 39301 5080 39313 5083
rect 36357 5043 36415 5049
rect 38672 5052 39313 5080
rect 27338 5012 27344 5024
rect 22066 4984 27344 5012
rect 15657 4975 15715 4981
rect 27338 4972 27344 4984
rect 27396 4972 27402 5024
rect 31478 4972 31484 5024
rect 31536 5012 31542 5024
rect 32401 5015 32459 5021
rect 32401 5012 32413 5015
rect 31536 4984 32413 5012
rect 31536 4972 31542 4984
rect 32401 4981 32413 4984
rect 32447 4981 32459 5015
rect 32401 4975 32459 4981
rect 35986 4972 35992 5024
rect 36044 5012 36050 5024
rect 38672 5021 38700 5052
rect 39301 5049 39313 5052
rect 39347 5049 39359 5083
rect 39301 5043 39359 5049
rect 40313 5083 40371 5089
rect 40313 5049 40325 5083
rect 40359 5080 40371 5083
rect 41138 5080 41144 5092
rect 40359 5052 41144 5080
rect 40359 5049 40371 5052
rect 40313 5043 40371 5049
rect 41138 5040 41144 5052
rect 41196 5040 41202 5092
rect 36173 5015 36231 5021
rect 36173 5012 36185 5015
rect 36044 4984 36185 5012
rect 36044 4972 36050 4984
rect 36173 4981 36185 4984
rect 36219 4981 36231 5015
rect 36173 4975 36231 4981
rect 38657 5015 38715 5021
rect 38657 4981 38669 5015
rect 38703 4981 38715 5015
rect 38657 4975 38715 4981
rect 38838 4972 38844 5024
rect 38896 4972 38902 5024
rect 42797 5015 42855 5021
rect 42797 4981 42809 5015
rect 42843 5012 42855 5015
rect 44082 5012 44088 5024
rect 42843 4984 44088 5012
rect 42843 4981 42855 4984
rect 42797 4975 42855 4981
rect 44082 4972 44088 4984
rect 44140 4972 44146 5024
rect 1104 4922 44896 4944
rect 1104 4870 6423 4922
rect 6475 4870 6487 4922
rect 6539 4870 6551 4922
rect 6603 4870 6615 4922
rect 6667 4870 6679 4922
rect 6731 4870 17370 4922
rect 17422 4870 17434 4922
rect 17486 4870 17498 4922
rect 17550 4870 17562 4922
rect 17614 4870 17626 4922
rect 17678 4870 28317 4922
rect 28369 4870 28381 4922
rect 28433 4870 28445 4922
rect 28497 4870 28509 4922
rect 28561 4870 28573 4922
rect 28625 4870 39264 4922
rect 39316 4870 39328 4922
rect 39380 4870 39392 4922
rect 39444 4870 39456 4922
rect 39508 4870 39520 4922
rect 39572 4870 44896 4922
rect 1104 4848 44896 4870
rect 4246 4768 4252 4820
rect 4304 4808 4310 4820
rect 4304 4780 13124 4808
rect 4304 4768 4310 4780
rect 13096 4740 13124 4780
rect 13170 4768 13176 4820
rect 13228 4768 13234 4820
rect 18414 4768 18420 4820
rect 18472 4768 18478 4820
rect 18984 4780 26648 4808
rect 18984 4752 19012 4780
rect 18966 4740 18972 4752
rect 13096 4712 18972 4740
rect 18966 4700 18972 4712
rect 19024 4700 19030 4752
rect 23017 4743 23075 4749
rect 23017 4740 23029 4743
rect 22066 4712 23029 4740
rect 4893 4675 4951 4681
rect 4893 4641 4905 4675
rect 4939 4672 4951 4675
rect 5810 4672 5816 4684
rect 4939 4644 5816 4672
rect 4939 4641 4951 4644
rect 4893 4635 4951 4641
rect 5810 4632 5816 4644
rect 5868 4632 5874 4684
rect 20530 4632 20536 4684
rect 20588 4632 20594 4684
rect 20806 4632 20812 4684
rect 20864 4672 20870 4684
rect 22066 4672 22094 4712
rect 23017 4709 23029 4712
rect 23063 4709 23075 4743
rect 23017 4703 23075 4709
rect 20864 4644 22094 4672
rect 22281 4675 22339 4681
rect 20864 4632 20870 4644
rect 22281 4641 22293 4675
rect 22327 4672 22339 4675
rect 22741 4675 22799 4681
rect 22741 4672 22753 4675
rect 22327 4644 22753 4672
rect 22327 4641 22339 4644
rect 22281 4635 22339 4641
rect 22741 4641 22753 4644
rect 22787 4641 22799 4675
rect 22741 4635 22799 4641
rect 5077 4607 5135 4613
rect 5077 4573 5089 4607
rect 5123 4604 5135 4607
rect 5258 4604 5264 4616
rect 5123 4576 5264 4604
rect 5123 4573 5135 4576
rect 5077 4567 5135 4573
rect 5258 4564 5264 4576
rect 5316 4564 5322 4616
rect 11793 4607 11851 4613
rect 11793 4573 11805 4607
rect 11839 4604 11851 4607
rect 11839 4576 12296 4604
rect 11839 4573 11851 4576
rect 11793 4567 11851 4573
rect 12268 4548 12296 4576
rect 15194 4564 15200 4616
rect 15252 4564 15258 4616
rect 15654 4564 15660 4616
rect 15712 4564 15718 4616
rect 17954 4564 17960 4616
rect 18012 4604 18018 4616
rect 18325 4607 18383 4613
rect 18325 4604 18337 4607
rect 18012 4576 18337 4604
rect 18012 4564 18018 4576
rect 18325 4573 18337 4576
rect 18371 4604 18383 4607
rect 18690 4604 18696 4616
rect 18371 4576 18696 4604
rect 18371 4573 18383 4576
rect 18325 4567 18383 4573
rect 18690 4564 18696 4576
rect 18748 4604 18754 4616
rect 19429 4607 19487 4613
rect 19429 4604 19441 4607
rect 18748 4576 19441 4604
rect 18748 4564 18754 4576
rect 19429 4573 19441 4576
rect 19475 4573 19487 4607
rect 19429 4567 19487 4573
rect 11606 4496 11612 4548
rect 11664 4536 11670 4548
rect 12038 4539 12096 4545
rect 12038 4536 12050 4539
rect 11664 4508 12050 4536
rect 11664 4496 11670 4508
rect 12038 4505 12050 4508
rect 12084 4505 12096 4539
rect 12038 4499 12096 4505
rect 12250 4496 12256 4548
rect 12308 4496 12314 4548
rect 17126 4496 17132 4548
rect 17184 4536 17190 4548
rect 17405 4539 17463 4545
rect 17405 4536 17417 4539
rect 17184 4508 17417 4536
rect 17184 4496 17190 4508
rect 17405 4505 17417 4508
rect 17451 4536 17463 4539
rect 17862 4536 17868 4548
rect 17451 4508 17868 4536
rect 17451 4505 17463 4508
rect 17405 4499 17463 4505
rect 17862 4496 17868 4508
rect 17920 4496 17926 4548
rect 19444 4536 19472 4567
rect 20714 4536 20720 4548
rect 19444 4508 20720 4536
rect 20714 4496 20720 4508
rect 20772 4496 20778 4548
rect 22094 4536 22100 4548
rect 22034 4508 22100 4536
rect 22094 4496 22100 4508
rect 22152 4496 22158 4548
rect 26620 4536 26648 4780
rect 27798 4768 27804 4820
rect 27856 4808 27862 4820
rect 28537 4811 28595 4817
rect 28537 4808 28549 4811
rect 27856 4780 28549 4808
rect 27856 4768 27862 4780
rect 28537 4777 28549 4780
rect 28583 4808 28595 4811
rect 32953 4811 33011 4817
rect 28583 4780 32904 4808
rect 28583 4777 28595 4780
rect 28537 4771 28595 4777
rect 32876 4740 32904 4780
rect 32953 4777 32965 4811
rect 32999 4808 33011 4811
rect 33686 4808 33692 4820
rect 32999 4780 33692 4808
rect 32999 4777 33011 4780
rect 32953 4771 33011 4777
rect 33686 4768 33692 4780
rect 33744 4768 33750 4820
rect 37182 4768 37188 4820
rect 37240 4768 37246 4820
rect 38010 4768 38016 4820
rect 38068 4808 38074 4820
rect 38381 4811 38439 4817
rect 38381 4808 38393 4811
rect 38068 4780 38393 4808
rect 38068 4768 38074 4780
rect 38381 4777 38393 4780
rect 38427 4777 38439 4811
rect 38381 4771 38439 4777
rect 33134 4740 33140 4752
rect 32876 4712 33140 4740
rect 33134 4700 33140 4712
rect 33192 4700 33198 4752
rect 33318 4700 33324 4752
rect 33376 4740 33382 4752
rect 33376 4712 33454 4740
rect 33376 4700 33382 4712
rect 26786 4632 26792 4684
rect 26844 4672 26850 4684
rect 27157 4675 27215 4681
rect 27157 4672 27169 4675
rect 26844 4644 27169 4672
rect 26844 4632 26850 4644
rect 27157 4641 27169 4644
rect 27203 4641 27215 4675
rect 27157 4635 27215 4641
rect 31202 4632 31208 4684
rect 31260 4632 31266 4684
rect 31478 4632 31484 4684
rect 31536 4632 31542 4684
rect 33426 4681 33454 4712
rect 33413 4675 33471 4681
rect 33413 4641 33425 4675
rect 33459 4641 33471 4675
rect 33413 4635 33471 4641
rect 35434 4632 35440 4684
rect 35492 4632 35498 4684
rect 27424 4607 27482 4613
rect 27424 4573 27436 4607
rect 27470 4604 27482 4607
rect 28166 4604 28172 4616
rect 27470 4576 28172 4604
rect 27470 4573 27482 4576
rect 27424 4567 27482 4573
rect 28166 4564 28172 4576
rect 28224 4564 28230 4616
rect 32858 4564 32864 4616
rect 32916 4604 32922 4616
rect 33781 4607 33839 4613
rect 33781 4604 33793 4607
rect 32916 4576 33793 4604
rect 32916 4564 32922 4576
rect 33781 4573 33793 4576
rect 33827 4573 33839 4607
rect 33781 4567 33839 4573
rect 33870 4564 33876 4616
rect 33928 4564 33934 4616
rect 37366 4564 37372 4616
rect 37424 4604 37430 4616
rect 37645 4607 37703 4613
rect 37645 4604 37657 4607
rect 37424 4576 37657 4604
rect 37424 4564 37430 4576
rect 37645 4573 37657 4576
rect 37691 4573 37703 4607
rect 37645 4567 37703 4573
rect 38565 4607 38623 4613
rect 38565 4573 38577 4607
rect 38611 4604 38623 4607
rect 38838 4604 38844 4616
rect 38611 4576 38844 4604
rect 38611 4573 38623 4576
rect 38565 4567 38623 4573
rect 38838 4564 38844 4576
rect 38896 4564 38902 4616
rect 44082 4564 44088 4616
rect 44140 4564 44146 4616
rect 27890 4536 27896 4548
rect 26620 4508 27896 4536
rect 27890 4496 27896 4508
rect 27948 4496 27954 4548
rect 33502 4536 33508 4548
rect 32706 4508 33508 4536
rect 33502 4496 33508 4508
rect 33560 4496 33566 4548
rect 35066 4496 35072 4548
rect 35124 4536 35130 4548
rect 35713 4539 35771 4545
rect 35713 4536 35725 4539
rect 35124 4508 35725 4536
rect 35124 4496 35130 4508
rect 35713 4505 35725 4508
rect 35759 4505 35771 4539
rect 37737 4539 37795 4545
rect 37737 4536 37749 4539
rect 36938 4508 37749 4536
rect 35713 4499 35771 4505
rect 37737 4505 37749 4508
rect 37783 4505 37795 4539
rect 37737 4499 37795 4505
rect 5261 4471 5319 4477
rect 5261 4437 5273 4471
rect 5307 4468 5319 4471
rect 5902 4468 5908 4480
rect 5307 4440 5908 4468
rect 5307 4437 5319 4440
rect 5261 4431 5319 4437
rect 5902 4428 5908 4440
rect 5960 4428 5966 4480
rect 14826 4428 14832 4480
rect 14884 4468 14890 4480
rect 15013 4471 15071 4477
rect 15013 4468 15025 4471
rect 14884 4440 15025 4468
rect 14884 4428 14890 4440
rect 15013 4437 15025 4440
rect 15059 4437 15071 4471
rect 15013 4431 15071 4437
rect 19426 4428 19432 4480
rect 19484 4468 19490 4480
rect 19521 4471 19579 4477
rect 19521 4468 19533 4471
rect 19484 4440 19533 4468
rect 19484 4428 19490 4440
rect 19521 4437 19533 4440
rect 19567 4437 19579 4471
rect 19521 4431 19579 4437
rect 23198 4428 23204 4480
rect 23256 4428 23262 4480
rect 33134 4428 33140 4480
rect 33192 4468 33198 4480
rect 33689 4471 33747 4477
rect 33689 4468 33701 4471
rect 33192 4440 33701 4468
rect 33192 4428 33198 4440
rect 33689 4437 33701 4440
rect 33735 4437 33747 4471
rect 33689 4431 33747 4437
rect 44266 4428 44272 4480
rect 44324 4428 44330 4480
rect 1104 4378 45051 4400
rect 1104 4326 11896 4378
rect 11948 4326 11960 4378
rect 12012 4326 12024 4378
rect 12076 4326 12088 4378
rect 12140 4326 12152 4378
rect 12204 4326 22843 4378
rect 22895 4326 22907 4378
rect 22959 4326 22971 4378
rect 23023 4326 23035 4378
rect 23087 4326 23099 4378
rect 23151 4326 33790 4378
rect 33842 4326 33854 4378
rect 33906 4326 33918 4378
rect 33970 4326 33982 4378
rect 34034 4326 34046 4378
rect 34098 4326 44737 4378
rect 44789 4326 44801 4378
rect 44853 4326 44865 4378
rect 44917 4326 44929 4378
rect 44981 4326 44993 4378
rect 45045 4326 45051 4378
rect 1104 4304 45051 4326
rect 13078 4224 13084 4276
rect 13136 4224 13142 4276
rect 13538 4224 13544 4276
rect 13596 4264 13602 4276
rect 42978 4264 42984 4276
rect 13596 4236 42984 4264
rect 13596 4224 13602 4236
rect 42978 4224 42984 4236
rect 43036 4224 43042 4276
rect 14826 4156 14832 4208
rect 14884 4156 14890 4208
rect 17586 4196 17592 4208
rect 16054 4168 17592 4196
rect 17586 4156 17592 4168
rect 17644 4156 17650 4208
rect 19426 4156 19432 4208
rect 19484 4156 19490 4208
rect 20714 4156 20720 4208
rect 20772 4196 20778 4208
rect 23934 4196 23940 4208
rect 20772 4168 23940 4196
rect 20772 4156 20778 4168
rect 12989 4131 13047 4137
rect 12989 4097 13001 4131
rect 13035 4097 13047 4131
rect 12989 4091 13047 4097
rect 13173 4131 13231 4137
rect 13173 4097 13185 4131
rect 13219 4128 13231 4131
rect 13219 4100 14504 4128
rect 13219 4097 13231 4100
rect 13173 4091 13231 4097
rect 13004 4060 13032 4091
rect 14274 4060 14280 4072
rect 13004 4032 14280 4060
rect 14274 4020 14280 4032
rect 14332 4020 14338 4072
rect 14476 3992 14504 4100
rect 16758 4088 16764 4140
rect 16816 4128 16822 4140
rect 16853 4131 16911 4137
rect 16853 4128 16865 4131
rect 16816 4100 16865 4128
rect 16816 4088 16822 4100
rect 16853 4097 16865 4100
rect 16899 4097 16911 4131
rect 16853 4091 16911 4097
rect 17497 4131 17555 4137
rect 17497 4097 17509 4131
rect 17543 4128 17555 4131
rect 17954 4128 17960 4140
rect 17543 4100 17960 4128
rect 17543 4097 17555 4100
rect 17497 4091 17555 4097
rect 17954 4088 17960 4100
rect 18012 4088 18018 4140
rect 22020 4137 22048 4168
rect 23934 4156 23940 4168
rect 23992 4156 23998 4208
rect 27798 4156 27804 4208
rect 27856 4156 27862 4208
rect 32416 4168 33272 4196
rect 22005 4131 22063 4137
rect 22005 4097 22017 4131
rect 22051 4097 22063 4131
rect 22005 4091 22063 4097
rect 22094 4088 22100 4140
rect 22152 4088 22158 4140
rect 22925 4131 22983 4137
rect 22925 4097 22937 4131
rect 22971 4128 22983 4131
rect 23198 4128 23204 4140
rect 22971 4100 23204 4128
rect 22971 4097 22983 4100
rect 22925 4091 22983 4097
rect 23198 4088 23204 4100
rect 23256 4088 23262 4140
rect 27890 4088 27896 4140
rect 27948 4088 27954 4140
rect 31573 4131 31631 4137
rect 31573 4097 31585 4131
rect 31619 4128 31631 4131
rect 32416 4128 32444 4168
rect 31619 4100 32444 4128
rect 32493 4131 32551 4137
rect 31619 4097 31631 4100
rect 31573 4091 31631 4097
rect 32493 4097 32505 4131
rect 32539 4128 32551 4131
rect 33134 4128 33140 4140
rect 32539 4100 33140 4128
rect 32539 4097 32551 4100
rect 32493 4091 32551 4097
rect 14550 4020 14556 4072
rect 14608 4020 14614 4072
rect 15286 4060 15292 4072
rect 14660 4032 15292 4060
rect 14660 3992 14688 4032
rect 15286 4020 15292 4032
rect 15344 4020 15350 4072
rect 17862 4020 17868 4072
rect 17920 4060 17926 4072
rect 18141 4063 18199 4069
rect 18141 4060 18153 4063
rect 17920 4032 18153 4060
rect 17920 4020 17926 4032
rect 18141 4029 18153 4032
rect 18187 4029 18199 4063
rect 18417 4063 18475 4069
rect 18417 4060 18429 4063
rect 18141 4023 18199 4029
rect 18248 4032 18429 4060
rect 14476 3964 14688 3992
rect 16301 3995 16359 4001
rect 16301 3961 16313 3995
rect 16347 3992 16359 3995
rect 18248 3992 18276 4032
rect 18417 4029 18429 4032
rect 18463 4029 18475 4063
rect 18417 4023 18475 4029
rect 19889 4063 19947 4069
rect 19889 4029 19901 4063
rect 19935 4060 19947 4063
rect 20806 4060 20812 4072
rect 19935 4032 20812 4060
rect 19935 4029 19947 4032
rect 19889 4023 19947 4029
rect 20806 4020 20812 4032
rect 20864 4020 20870 4072
rect 27982 4020 27988 4072
rect 28040 4020 28046 4072
rect 16347 3964 18276 3992
rect 22741 3995 22799 4001
rect 16347 3961 16359 3964
rect 16301 3955 16359 3961
rect 22741 3961 22753 3995
rect 22787 3992 22799 3995
rect 23290 3992 23296 4004
rect 22787 3964 23296 3992
rect 22787 3961 22799 3964
rect 22741 3955 22799 3961
rect 23290 3952 23296 3964
rect 23348 3952 23354 4004
rect 27430 3952 27436 4004
rect 27488 3952 27494 4004
rect 15838 3884 15844 3936
rect 15896 3924 15902 3936
rect 16945 3927 17003 3933
rect 16945 3924 16957 3927
rect 15896 3896 16957 3924
rect 15896 3884 15902 3896
rect 16945 3893 16957 3896
rect 16991 3893 17003 3927
rect 16945 3887 17003 3893
rect 17586 3884 17592 3936
rect 17644 3884 17650 3936
rect 23750 3884 23756 3936
rect 23808 3924 23814 3936
rect 31018 3924 31024 3936
rect 23808 3896 31024 3924
rect 23808 3884 23814 3896
rect 31018 3884 31024 3896
rect 31076 3924 31082 3936
rect 31588 3924 31616 4091
rect 33134 4088 33140 4100
rect 33192 4088 33198 4140
rect 33244 4128 33272 4168
rect 38194 4156 38200 4208
rect 38252 4156 38258 4208
rect 33413 4131 33471 4137
rect 33413 4128 33425 4131
rect 33244 4100 33425 4128
rect 33413 4097 33425 4100
rect 33459 4097 33471 4131
rect 33413 4091 33471 4097
rect 32122 4020 32128 4072
rect 32180 4060 32186 4072
rect 32677 4063 32735 4069
rect 32677 4060 32689 4063
rect 32180 4032 32689 4060
rect 32180 4020 32186 4032
rect 32677 4029 32689 4032
rect 32723 4029 32735 4063
rect 32677 4023 32735 4029
rect 32769 4063 32827 4069
rect 32769 4029 32781 4063
rect 32815 4029 32827 4063
rect 33428 4060 33456 4091
rect 33502 4088 33508 4140
rect 33560 4088 33566 4140
rect 35253 4131 35311 4137
rect 35253 4097 35265 4131
rect 35299 4128 35311 4131
rect 35894 4128 35900 4140
rect 35299 4100 35900 4128
rect 35299 4097 35311 4100
rect 35253 4091 35311 4097
rect 35894 4088 35900 4100
rect 35952 4088 35958 4140
rect 36354 4088 36360 4140
rect 36412 4088 36418 4140
rect 37366 4128 37372 4140
rect 36648 4100 37372 4128
rect 33428 4032 36216 4060
rect 32769 4023 32827 4029
rect 31938 3952 31944 4004
rect 31996 3992 32002 4004
rect 32784 3992 32812 4023
rect 32858 3992 32864 4004
rect 31996 3964 32864 3992
rect 31996 3952 32002 3964
rect 32858 3952 32864 3964
rect 32916 3952 32922 4004
rect 35066 3952 35072 4004
rect 35124 3952 35130 4004
rect 36188 3992 36216 4032
rect 36262 4020 36268 4072
rect 36320 4020 36326 4072
rect 36648 3992 36676 4100
rect 37366 4088 37372 4100
rect 37424 4088 37430 4140
rect 37458 4088 37464 4140
rect 37516 4088 37522 4140
rect 37737 4063 37795 4069
rect 37737 4060 37749 4063
rect 36740 4032 37749 4060
rect 36740 4001 36768 4032
rect 37737 4029 37749 4032
rect 37783 4029 37795 4063
rect 37737 4023 37795 4029
rect 36188 3964 36676 3992
rect 36725 3995 36783 4001
rect 36725 3961 36737 3995
rect 36771 3961 36783 3995
rect 36725 3955 36783 3961
rect 31076 3896 31616 3924
rect 31076 3884 31082 3896
rect 31662 3884 31668 3936
rect 31720 3884 31726 3936
rect 32030 3884 32036 3936
rect 32088 3924 32094 3936
rect 32309 3927 32367 3933
rect 32309 3924 32321 3927
rect 32088 3896 32321 3924
rect 32088 3884 32094 3896
rect 32309 3893 32321 3896
rect 32355 3893 32367 3927
rect 32309 3887 32367 3893
rect 36354 3884 36360 3936
rect 36412 3924 36418 3936
rect 39209 3927 39267 3933
rect 39209 3924 39221 3927
rect 36412 3896 39221 3924
rect 36412 3884 36418 3896
rect 39209 3893 39221 3896
rect 39255 3924 39267 3927
rect 44082 3924 44088 3936
rect 39255 3896 44088 3924
rect 39255 3893 39267 3896
rect 39209 3887 39267 3893
rect 44082 3884 44088 3896
rect 44140 3884 44146 3936
rect 1104 3834 44896 3856
rect 1104 3782 6423 3834
rect 6475 3782 6487 3834
rect 6539 3782 6551 3834
rect 6603 3782 6615 3834
rect 6667 3782 6679 3834
rect 6731 3782 17370 3834
rect 17422 3782 17434 3834
rect 17486 3782 17498 3834
rect 17550 3782 17562 3834
rect 17614 3782 17626 3834
rect 17678 3782 28317 3834
rect 28369 3782 28381 3834
rect 28433 3782 28445 3834
rect 28497 3782 28509 3834
rect 28561 3782 28573 3834
rect 28625 3782 39264 3834
rect 39316 3782 39328 3834
rect 39380 3782 39392 3834
rect 39444 3782 39456 3834
rect 39508 3782 39520 3834
rect 39572 3782 44896 3834
rect 1104 3760 44896 3782
rect 9950 3680 9956 3732
rect 10008 3720 10014 3732
rect 26878 3720 26884 3732
rect 10008 3692 26884 3720
rect 10008 3680 10014 3692
rect 26878 3680 26884 3692
rect 26936 3680 26942 3732
rect 31376 3723 31434 3729
rect 31376 3689 31388 3723
rect 31422 3720 31434 3723
rect 32030 3720 32036 3732
rect 31422 3692 32036 3720
rect 31422 3689 31434 3692
rect 31376 3683 31434 3689
rect 32030 3680 32036 3692
rect 32088 3680 32094 3732
rect 32858 3680 32864 3732
rect 32916 3680 32922 3732
rect 37553 3723 37611 3729
rect 37553 3689 37565 3723
rect 37599 3720 37611 3723
rect 38194 3720 38200 3732
rect 37599 3692 38200 3720
rect 37599 3689 37611 3692
rect 37553 3683 37611 3689
rect 38194 3680 38200 3692
rect 38252 3680 38258 3732
rect 22373 3655 22431 3661
rect 22373 3621 22385 3655
rect 22419 3652 22431 3655
rect 23750 3652 23756 3664
rect 22419 3624 23756 3652
rect 22419 3621 22431 3624
rect 22373 3615 22431 3621
rect 23750 3612 23756 3624
rect 23808 3612 23814 3664
rect 23382 3544 23388 3596
rect 23440 3584 23446 3596
rect 33502 3584 33508 3596
rect 23440 3556 33508 3584
rect 23440 3544 23446 3556
rect 33502 3544 33508 3556
rect 33560 3544 33566 3596
rect 934 3476 940 3528
rect 992 3516 998 3528
rect 1765 3519 1823 3525
rect 1765 3516 1777 3519
rect 992 3488 1777 3516
rect 992 3476 998 3488
rect 1765 3485 1777 3488
rect 1811 3485 1823 3519
rect 1765 3479 1823 3485
rect 5902 3476 5908 3528
rect 5960 3476 5966 3528
rect 14550 3476 14556 3528
rect 14608 3476 14614 3528
rect 14826 3476 14832 3528
rect 14884 3516 14890 3528
rect 15657 3519 15715 3525
rect 15657 3516 15669 3519
rect 14884 3488 15669 3516
rect 14884 3476 14890 3488
rect 15657 3485 15669 3488
rect 15703 3485 15715 3519
rect 15657 3479 15715 3485
rect 16669 3519 16727 3525
rect 16669 3485 16681 3519
rect 16715 3516 16727 3519
rect 16942 3516 16948 3528
rect 16715 3488 16948 3516
rect 16715 3485 16727 3488
rect 16669 3479 16727 3485
rect 16942 3476 16948 3488
rect 17000 3476 17006 3528
rect 17034 3476 17040 3528
rect 17092 3476 17098 3528
rect 17862 3476 17868 3528
rect 17920 3516 17926 3528
rect 19429 3519 19487 3525
rect 19429 3516 19441 3519
rect 17920 3488 19441 3516
rect 17920 3476 17926 3488
rect 19429 3485 19441 3488
rect 19475 3516 19487 3519
rect 20530 3516 20536 3528
rect 19475 3488 20536 3516
rect 19475 3485 19487 3488
rect 19429 3479 19487 3485
rect 20530 3476 20536 3488
rect 20588 3476 20594 3528
rect 31110 3476 31116 3528
rect 31168 3476 31174 3528
rect 37366 3476 37372 3528
rect 37424 3516 37430 3528
rect 37461 3519 37519 3525
rect 37461 3516 37473 3519
rect 37424 3488 37473 3516
rect 37424 3476 37430 3488
rect 37461 3485 37473 3488
rect 37507 3485 37519 3519
rect 37461 3479 37519 3485
rect 44361 3519 44419 3525
rect 44361 3485 44373 3519
rect 44407 3516 44419 3519
rect 44634 3516 44640 3528
rect 44407 3488 44640 3516
rect 44407 3485 44419 3488
rect 44361 3479 44419 3485
rect 44634 3476 44640 3488
rect 44692 3476 44698 3528
rect 14568 3448 14596 3476
rect 16574 3448 16580 3460
rect 14568 3420 16580 3448
rect 16574 3408 16580 3420
rect 16632 3408 16638 3460
rect 18463 3451 18521 3457
rect 17328 3420 17434 3448
rect 5718 3340 5724 3392
rect 5776 3340 5782 3392
rect 14458 3340 14464 3392
rect 14516 3380 14522 3392
rect 14645 3383 14703 3389
rect 14645 3380 14657 3383
rect 14516 3352 14657 3380
rect 14516 3340 14522 3352
rect 14645 3349 14657 3352
rect 14691 3349 14703 3383
rect 14645 3343 14703 3349
rect 17034 3340 17040 3392
rect 17092 3380 17098 3392
rect 17328 3380 17356 3420
rect 18463 3417 18475 3451
rect 18509 3448 18521 3451
rect 18874 3448 18880 3460
rect 18509 3420 18880 3448
rect 18509 3417 18521 3420
rect 18463 3411 18521 3417
rect 18874 3408 18880 3420
rect 18932 3408 18938 3460
rect 22094 3408 22100 3460
rect 22152 3408 22158 3460
rect 31662 3408 31668 3460
rect 31720 3448 31726 3460
rect 36354 3448 36360 3460
rect 31720 3420 31878 3448
rect 32784 3420 36360 3448
rect 31720 3408 31726 3420
rect 17092 3352 17356 3380
rect 17092 3340 17098 3352
rect 18598 3340 18604 3392
rect 18656 3380 18662 3392
rect 19521 3383 19579 3389
rect 19521 3380 19533 3383
rect 18656 3352 19533 3380
rect 18656 3340 18662 3352
rect 19521 3349 19533 3352
rect 19567 3349 19579 3383
rect 19521 3343 19579 3349
rect 30282 3340 30288 3392
rect 30340 3380 30346 3392
rect 32784 3380 32812 3420
rect 36354 3408 36360 3420
rect 36412 3408 36418 3460
rect 30340 3352 32812 3380
rect 30340 3340 30346 3352
rect 1104 3290 45051 3312
rect 1104 3238 11896 3290
rect 11948 3238 11960 3290
rect 12012 3238 12024 3290
rect 12076 3238 12088 3290
rect 12140 3238 12152 3290
rect 12204 3238 22843 3290
rect 22895 3238 22907 3290
rect 22959 3238 22971 3290
rect 23023 3238 23035 3290
rect 23087 3238 23099 3290
rect 23151 3238 33790 3290
rect 33842 3238 33854 3290
rect 33906 3238 33918 3290
rect 33970 3238 33982 3290
rect 34034 3238 34046 3290
rect 34098 3238 44737 3290
rect 44789 3238 44801 3290
rect 44853 3238 44865 3290
rect 44917 3238 44929 3290
rect 44981 3238 44993 3290
rect 45045 3238 45051 3290
rect 1104 3216 45051 3238
rect 9677 3179 9735 3185
rect 9677 3145 9689 3179
rect 9723 3176 9735 3179
rect 16255 3179 16313 3185
rect 9723 3148 12434 3176
rect 9723 3145 9735 3148
rect 9677 3139 9735 3145
rect 7742 3000 7748 3052
rect 7800 3000 7806 3052
rect 9398 3000 9404 3052
rect 9456 3040 9462 3052
rect 9493 3043 9551 3049
rect 9493 3040 9505 3043
rect 9456 3012 9505 3040
rect 9456 3000 9462 3012
rect 9493 3009 9505 3012
rect 9539 3009 9551 3043
rect 12406 3040 12434 3148
rect 16255 3145 16267 3179
rect 16301 3176 16313 3179
rect 16850 3176 16856 3188
rect 16301 3148 16856 3176
rect 16301 3145 16313 3148
rect 16255 3139 16313 3145
rect 16850 3136 16856 3148
rect 16908 3136 16914 3188
rect 16942 3136 16948 3188
rect 17000 3136 17006 3188
rect 17589 3179 17647 3185
rect 17589 3145 17601 3179
rect 17635 3176 17647 3179
rect 20303 3179 20361 3185
rect 17635 3148 19196 3176
rect 17635 3145 17647 3148
rect 17589 3139 17647 3145
rect 15838 3068 15844 3120
rect 15896 3068 15902 3120
rect 16574 3068 16580 3120
rect 16632 3108 16638 3120
rect 17862 3108 17868 3120
rect 16632 3080 17868 3108
rect 16632 3068 16638 3080
rect 14001 3043 14059 3049
rect 14001 3040 14013 3043
rect 12406 3012 14013 3040
rect 9493 3003 9551 3009
rect 14001 3009 14013 3012
rect 14047 3009 14059 3043
rect 14001 3003 14059 3009
rect 14458 3000 14464 3052
rect 14516 3000 14522 3052
rect 14826 3000 14832 3052
rect 14884 3000 14890 3052
rect 16868 3049 16896 3080
rect 17862 3068 17868 3080
rect 17920 3068 17926 3120
rect 19168 3108 19196 3148
rect 20303 3145 20315 3179
rect 20349 3176 20361 3179
rect 22094 3176 22100 3188
rect 20349 3148 22100 3176
rect 20349 3145 20361 3148
rect 20303 3139 20361 3145
rect 22094 3136 22100 3148
rect 22152 3136 22158 3188
rect 26878 3136 26884 3188
rect 26936 3176 26942 3188
rect 33873 3179 33931 3185
rect 33873 3176 33885 3179
rect 26936 3148 33885 3176
rect 26936 3136 26942 3148
rect 33873 3145 33885 3148
rect 33919 3145 33931 3179
rect 33873 3139 33931 3145
rect 44177 3179 44235 3185
rect 44177 3145 44189 3179
rect 44223 3176 44235 3179
rect 44450 3176 44456 3188
rect 44223 3148 44456 3176
rect 44223 3145 44235 3148
rect 44177 3139 44235 3145
rect 19168 3080 19274 3108
rect 16853 3043 16911 3049
rect 16853 3009 16865 3043
rect 16899 3009 16911 3043
rect 16853 3003 16911 3009
rect 17497 3043 17555 3049
rect 17497 3009 17509 3043
rect 17543 3009 17555 3043
rect 17497 3003 17555 3009
rect 18509 3043 18567 3049
rect 18509 3009 18521 3043
rect 18555 3040 18567 3043
rect 18598 3040 18604 3052
rect 18555 3012 18604 3040
rect 18555 3009 18567 3012
rect 18509 3003 18567 3009
rect 16758 2932 16764 2984
rect 16816 2972 16822 2984
rect 17512 2972 17540 3003
rect 18598 3000 18604 3012
rect 18656 3000 18662 3052
rect 18874 3000 18880 3052
rect 18932 3000 18938 3052
rect 22462 3000 22468 3052
rect 22520 3000 22526 3052
rect 33888 3040 33916 3139
rect 44450 3136 44456 3148
rect 44508 3136 44514 3188
rect 34241 3043 34299 3049
rect 34241 3040 34253 3043
rect 33888 3012 34253 3040
rect 34241 3009 34253 3012
rect 34287 3009 34299 3043
rect 34241 3003 34299 3009
rect 44361 3043 44419 3049
rect 44361 3009 44373 3043
rect 44407 3040 44419 3043
rect 45094 3040 45100 3052
rect 44407 3012 45100 3040
rect 44407 3009 44419 3012
rect 44361 3003 44419 3009
rect 45094 3000 45100 3012
rect 45152 3000 45158 3052
rect 16816 2944 17540 2972
rect 16816 2932 16822 2944
rect 934 2796 940 2848
rect 992 2836 998 2848
rect 1765 2839 1823 2845
rect 1765 2836 1777 2839
rect 992 2808 1777 2836
rect 992 2796 998 2808
rect 1765 2805 1777 2808
rect 1811 2805 1823 2839
rect 1765 2799 1823 2805
rect 7561 2839 7619 2845
rect 7561 2805 7573 2839
rect 7607 2836 7619 2839
rect 9582 2836 9588 2848
rect 7607 2808 9588 2836
rect 7607 2805 7619 2808
rect 7561 2799 7619 2805
rect 9582 2796 9588 2808
rect 9640 2796 9646 2848
rect 13817 2839 13875 2845
rect 13817 2805 13829 2839
rect 13863 2836 13875 2839
rect 14182 2836 14188 2848
rect 13863 2808 14188 2836
rect 13863 2805 13875 2808
rect 13817 2799 13875 2805
rect 14182 2796 14188 2808
rect 14240 2796 14246 2848
rect 22281 2839 22339 2845
rect 22281 2805 22293 2839
rect 22327 2836 22339 2839
rect 22646 2836 22652 2848
rect 22327 2808 22652 2836
rect 22327 2805 22339 2808
rect 22281 2799 22339 2805
rect 22646 2796 22652 2808
rect 22704 2796 22710 2848
rect 34425 2839 34483 2845
rect 34425 2805 34437 2839
rect 34471 2836 34483 2839
rect 35526 2836 35532 2848
rect 34471 2808 35532 2836
rect 34471 2805 34483 2808
rect 34425 2799 34483 2805
rect 35526 2796 35532 2808
rect 35584 2796 35590 2848
rect 1104 2746 44896 2768
rect 1104 2694 6423 2746
rect 6475 2694 6487 2746
rect 6539 2694 6551 2746
rect 6603 2694 6615 2746
rect 6667 2694 6679 2746
rect 6731 2694 17370 2746
rect 17422 2694 17434 2746
rect 17486 2694 17498 2746
rect 17550 2694 17562 2746
rect 17614 2694 17626 2746
rect 17678 2694 28317 2746
rect 28369 2694 28381 2746
rect 28433 2694 28445 2746
rect 28497 2694 28509 2746
rect 28561 2694 28573 2746
rect 28625 2694 39264 2746
rect 39316 2694 39328 2746
rect 39380 2694 39392 2746
rect 39444 2694 39456 2746
rect 39508 2694 39520 2746
rect 39572 2694 44896 2746
rect 1104 2672 44896 2694
rect 16945 2635 17003 2641
rect 16945 2601 16957 2635
rect 16991 2632 17003 2635
rect 17126 2632 17132 2644
rect 16991 2604 17132 2632
rect 16991 2601 17003 2604
rect 16945 2595 17003 2601
rect 17126 2592 17132 2604
rect 17184 2592 17190 2644
rect 27338 2592 27344 2644
rect 27396 2592 27402 2644
rect 37461 2635 37519 2641
rect 37461 2601 37473 2635
rect 37507 2632 37519 2635
rect 38102 2632 38108 2644
rect 37507 2604 38108 2632
rect 37507 2601 37519 2604
rect 37461 2595 37519 2601
rect 38102 2592 38108 2604
rect 38160 2592 38166 2644
rect 43438 2592 43444 2644
rect 43496 2592 43502 2644
rect 30190 2524 30196 2576
rect 30248 2564 30254 2576
rect 42889 2567 42947 2573
rect 42889 2564 42901 2567
rect 30248 2536 42901 2564
rect 30248 2524 30254 2536
rect 42889 2533 42901 2536
rect 42935 2533 42947 2567
rect 42889 2527 42947 2533
rect 14 2456 20 2508
rect 72 2496 78 2508
rect 2409 2499 2467 2505
rect 2409 2496 2421 2499
rect 72 2468 2421 2496
rect 72 2456 78 2468
rect 2409 2465 2421 2468
rect 2455 2465 2467 2499
rect 2409 2459 2467 2465
rect 12802 2456 12808 2508
rect 12860 2496 12866 2508
rect 13173 2499 13231 2505
rect 13173 2496 13185 2499
rect 12860 2468 13185 2496
rect 12860 2456 12866 2468
rect 13173 2465 13185 2468
rect 13219 2465 13231 2499
rect 17773 2499 17831 2505
rect 17773 2496 17785 2499
rect 13173 2459 13231 2465
rect 16868 2468 17785 2496
rect 1302 2388 1308 2440
rect 1360 2428 1366 2440
rect 1765 2431 1823 2437
rect 1765 2428 1777 2431
rect 1360 2400 1777 2428
rect 1360 2388 1366 2400
rect 1765 2397 1777 2400
rect 1811 2397 1823 2431
rect 1765 2391 1823 2397
rect 4154 2388 4160 2440
rect 4212 2388 4218 2440
rect 4522 2388 4528 2440
rect 4580 2428 4586 2440
rect 4801 2431 4859 2437
rect 4801 2428 4813 2431
rect 4580 2400 4813 2428
rect 4580 2388 4586 2400
rect 4801 2397 4813 2400
rect 4847 2397 4859 2431
rect 4801 2391 4859 2397
rect 5718 2388 5724 2440
rect 5776 2428 5782 2440
rect 6549 2431 6607 2437
rect 6549 2428 6561 2431
rect 5776 2400 6561 2428
rect 5776 2388 5782 2400
rect 6549 2397 6561 2400
rect 6595 2397 6607 2431
rect 6549 2391 6607 2397
rect 7742 2388 7748 2440
rect 7800 2428 7806 2440
rect 8021 2431 8079 2437
rect 8021 2428 8033 2431
rect 7800 2400 8033 2428
rect 7800 2388 7806 2400
rect 8021 2397 8033 2400
rect 8067 2397 8079 2431
rect 8021 2391 8079 2397
rect 9582 2388 9588 2440
rect 9640 2428 9646 2440
rect 9769 2431 9827 2437
rect 9769 2428 9781 2431
rect 9640 2400 9781 2428
rect 9640 2388 9646 2400
rect 9769 2397 9781 2400
rect 9815 2397 9827 2431
rect 9769 2391 9827 2397
rect 11054 2388 11060 2440
rect 11112 2428 11118 2440
rect 11885 2431 11943 2437
rect 11885 2428 11897 2431
rect 11112 2400 11897 2428
rect 11112 2388 11118 2400
rect 11885 2397 11897 2400
rect 11931 2397 11943 2431
rect 11885 2391 11943 2397
rect 12894 2388 12900 2440
rect 12952 2388 12958 2440
rect 15657 2431 15715 2437
rect 15657 2397 15669 2431
rect 15703 2428 15715 2431
rect 16114 2428 16120 2440
rect 15703 2400 16120 2428
rect 15703 2397 15715 2400
rect 15657 2391 15715 2397
rect 16114 2388 16120 2400
rect 16172 2388 16178 2440
rect 16758 2388 16764 2440
rect 16816 2428 16822 2440
rect 16868 2437 16896 2468
rect 17773 2465 17785 2468
rect 17819 2465 17831 2499
rect 17773 2459 17831 2465
rect 32582 2456 32588 2508
rect 32640 2456 32646 2508
rect 16853 2431 16911 2437
rect 16853 2428 16865 2431
rect 16816 2400 16865 2428
rect 16816 2388 16822 2400
rect 16853 2397 16865 2400
rect 16899 2397 16911 2431
rect 16853 2391 16911 2397
rect 17402 2388 17408 2440
rect 17460 2428 17466 2440
rect 17497 2431 17555 2437
rect 17497 2428 17509 2431
rect 17460 2400 17509 2428
rect 17460 2388 17466 2400
rect 17497 2397 17509 2400
rect 17543 2397 17555 2431
rect 17497 2391 17555 2397
rect 19334 2388 19340 2440
rect 19392 2428 19398 2440
rect 19613 2431 19671 2437
rect 19613 2428 19625 2431
rect 19392 2400 19625 2428
rect 19392 2388 19398 2400
rect 19613 2397 19625 2400
rect 19659 2397 19671 2431
rect 19613 2391 19671 2397
rect 20714 2388 20720 2440
rect 20772 2428 20778 2440
rect 20901 2431 20959 2437
rect 20901 2428 20913 2431
rect 20772 2400 20913 2428
rect 20772 2388 20778 2400
rect 20901 2397 20913 2400
rect 20947 2397 20959 2431
rect 20901 2391 20959 2397
rect 22646 2388 22652 2440
rect 22704 2388 22710 2440
rect 23842 2388 23848 2440
rect 23900 2428 23906 2440
rect 24765 2431 24823 2437
rect 24765 2428 24777 2431
rect 23900 2400 24777 2428
rect 23900 2388 23906 2400
rect 24765 2397 24777 2400
rect 24811 2397 24823 2431
rect 24765 2391 24823 2397
rect 25774 2388 25780 2440
rect 25832 2428 25838 2440
rect 26053 2431 26111 2437
rect 26053 2428 26065 2431
rect 25832 2400 26065 2428
rect 25832 2388 25838 2400
rect 26053 2397 26065 2400
rect 26099 2397 26111 2431
rect 26053 2391 26111 2397
rect 27062 2388 27068 2440
rect 27120 2428 27126 2440
rect 27157 2431 27215 2437
rect 27157 2428 27169 2431
rect 27120 2400 27169 2428
rect 27120 2388 27126 2400
rect 27157 2397 27169 2400
rect 27203 2397 27215 2431
rect 27157 2391 27215 2397
rect 28994 2388 29000 2440
rect 29052 2428 29058 2440
rect 29917 2431 29975 2437
rect 29917 2428 29929 2431
rect 29052 2400 29929 2428
rect 29052 2388 29058 2400
rect 29917 2397 29929 2400
rect 29963 2397 29975 2431
rect 29917 2391 29975 2397
rect 30374 2388 30380 2440
rect 30432 2428 30438 2440
rect 30561 2431 30619 2437
rect 30561 2428 30573 2431
rect 30432 2400 30573 2428
rect 30432 2388 30438 2400
rect 30561 2397 30573 2400
rect 30607 2397 30619 2431
rect 30561 2391 30619 2397
rect 32214 2388 32220 2440
rect 32272 2428 32278 2440
rect 32309 2431 32367 2437
rect 32309 2428 32321 2431
rect 32272 2400 32321 2428
rect 32272 2388 32278 2400
rect 32309 2397 32321 2400
rect 32355 2397 32367 2431
rect 32309 2391 32367 2397
rect 35526 2388 35532 2440
rect 35584 2388 35590 2440
rect 37642 2388 37648 2440
rect 37700 2388 37706 2440
rect 38654 2388 38660 2440
rect 38712 2428 38718 2440
rect 38933 2431 38991 2437
rect 38933 2428 38945 2431
rect 38712 2400 38945 2428
rect 38712 2388 38718 2400
rect 38933 2397 38945 2400
rect 38979 2397 38991 2431
rect 38933 2391 38991 2397
rect 40034 2388 40040 2440
rect 40092 2428 40098 2440
rect 40221 2431 40279 2437
rect 40221 2428 40233 2431
rect 40092 2400 40233 2428
rect 40092 2388 40098 2400
rect 40221 2397 40233 2400
rect 40267 2397 40279 2431
rect 40221 2391 40279 2397
rect 43625 2431 43683 2437
rect 43625 2397 43637 2431
rect 43671 2428 43683 2431
rect 43806 2428 43812 2440
rect 43671 2400 43812 2428
rect 43671 2397 43683 2400
rect 43625 2391 43683 2397
rect 43806 2388 43812 2400
rect 43864 2388 43870 2440
rect 44082 2388 44088 2440
rect 44140 2388 44146 2440
rect 41874 2320 41880 2372
rect 41932 2360 41938 2372
rect 42705 2363 42763 2369
rect 42705 2360 42717 2363
rect 41932 2332 42717 2360
rect 41932 2320 41938 2332
rect 42705 2329 42717 2332
rect 42751 2329 42763 2363
rect 42705 2323 42763 2329
rect 6454 2252 6460 2304
rect 6512 2292 6518 2304
rect 6733 2295 6791 2301
rect 6733 2292 6745 2295
rect 6512 2264 6745 2292
rect 6512 2252 6518 2264
rect 6733 2261 6745 2264
rect 6779 2261 6791 2295
rect 6733 2255 6791 2261
rect 9674 2252 9680 2304
rect 9732 2292 9738 2304
rect 9953 2295 10011 2301
rect 9953 2292 9965 2295
rect 9732 2264 9965 2292
rect 9732 2252 9738 2264
rect 9953 2261 9965 2264
rect 9999 2261 10011 2295
rect 9953 2255 10011 2261
rect 22554 2252 22560 2304
rect 22612 2292 22618 2304
rect 22833 2295 22891 2301
rect 22833 2292 22845 2295
rect 22612 2264 22845 2292
rect 22612 2252 22618 2264
rect 22833 2261 22845 2264
rect 22879 2261 22891 2295
rect 22833 2255 22891 2261
rect 25869 2295 25927 2301
rect 25869 2261 25881 2295
rect 25915 2292 25927 2295
rect 31846 2292 31852 2304
rect 25915 2264 31852 2292
rect 25915 2261 25927 2264
rect 25869 2255 25927 2261
rect 31846 2252 31852 2264
rect 31904 2252 31910 2304
rect 35434 2252 35440 2304
rect 35492 2292 35498 2304
rect 35713 2295 35771 2301
rect 35713 2292 35725 2295
rect 35492 2264 35725 2292
rect 35492 2252 35498 2264
rect 35713 2261 35725 2264
rect 35759 2261 35771 2295
rect 35713 2255 35771 2261
rect 44266 2252 44272 2304
rect 44324 2252 44330 2304
rect 1104 2202 45051 2224
rect 1104 2150 11896 2202
rect 11948 2150 11960 2202
rect 12012 2150 12024 2202
rect 12076 2150 12088 2202
rect 12140 2150 12152 2202
rect 12204 2150 22843 2202
rect 22895 2150 22907 2202
rect 22959 2150 22971 2202
rect 23023 2150 23035 2202
rect 23087 2150 23099 2202
rect 23151 2150 33790 2202
rect 33842 2150 33854 2202
rect 33906 2150 33918 2202
rect 33970 2150 33982 2202
rect 34034 2150 34046 2202
rect 34098 2150 44737 2202
rect 44789 2150 44801 2202
rect 44853 2150 44865 2202
rect 44917 2150 44929 2202
rect 44981 2150 44993 2202
rect 45045 2150 45051 2202
rect 1104 2128 45051 2150
rect 3234 892 3240 944
rect 3292 932 3298 944
rect 4154 932 4160 944
rect 3292 904 4160 932
rect 3292 892 3298 904
rect 4154 892 4160 904
rect 4212 892 4218 944
rect 36722 892 36728 944
rect 36780 932 36786 944
rect 37642 932 37648 944
rect 36780 904 37648 932
rect 36780 892 36786 904
rect 37642 892 37648 904
rect 37700 892 37706 944
<< via1 >>
rect 34152 19048 34204 19100
rect 35072 19048 35124 19100
rect 41880 19048 41932 19100
rect 42800 19048 42852 19100
rect 43720 17960 43772 18012
rect 45008 17960 45060 18012
rect 11896 17382 11948 17434
rect 11960 17382 12012 17434
rect 12024 17382 12076 17434
rect 12088 17382 12140 17434
rect 12152 17382 12204 17434
rect 22843 17382 22895 17434
rect 22907 17382 22959 17434
rect 22971 17382 23023 17434
rect 23035 17382 23087 17434
rect 23099 17382 23151 17434
rect 33790 17382 33842 17434
rect 33854 17382 33906 17434
rect 33918 17382 33970 17434
rect 33982 17382 34034 17434
rect 34046 17382 34098 17434
rect 44737 17382 44789 17434
rect 44801 17382 44853 17434
rect 44865 17382 44917 17434
rect 44929 17382 44981 17434
rect 44993 17382 45045 17434
rect 17408 17280 17460 17332
rect 20720 17280 20772 17332
rect 40592 17280 40644 17332
rect 44272 17323 44324 17332
rect 44272 17289 44281 17323
rect 44281 17289 44315 17323
rect 44315 17289 44324 17323
rect 44272 17280 44324 17289
rect 1308 17212 1360 17264
rect 3240 17255 3292 17264
rect 3240 17221 3249 17255
rect 3249 17221 3283 17255
rect 3283 17221 3292 17255
rect 3240 17212 3292 17221
rect 4528 17212 4580 17264
rect 11060 17212 11112 17264
rect 16120 17255 16172 17264
rect 16120 17221 16129 17255
rect 16129 17221 16163 17255
rect 16163 17221 16172 17255
rect 16120 17212 16172 17221
rect 32220 17212 32272 17264
rect 38660 17212 38712 17264
rect 940 17144 992 17196
rect 6460 17144 6512 17196
rect 7748 17144 7800 17196
rect 9680 17144 9732 17196
rect 12900 17144 12952 17196
rect 14188 17144 14240 17196
rect 16580 17144 16632 17196
rect 19340 17144 19392 17196
rect 20720 17187 20772 17196
rect 20720 17153 20729 17187
rect 20729 17153 20763 17187
rect 20763 17153 20772 17187
rect 20720 17144 20772 17153
rect 22560 17144 22612 17196
rect 23848 17144 23900 17196
rect 25780 17144 25832 17196
rect 27712 17144 27764 17196
rect 29000 17144 29052 17196
rect 30932 17144 30984 17196
rect 35072 17187 35124 17196
rect 35072 17153 35081 17187
rect 35081 17153 35115 17187
rect 35115 17153 35124 17187
rect 35072 17144 35124 17153
rect 35440 17144 35492 17196
rect 37372 17144 37424 17196
rect 40684 17187 40736 17196
rect 40684 17153 40693 17187
rect 40693 17153 40727 17187
rect 40727 17153 40736 17187
rect 40684 17144 40736 17153
rect 42800 17187 42852 17196
rect 42800 17153 42809 17187
rect 42809 17153 42843 17187
rect 42843 17153 42852 17187
rect 42800 17144 42852 17153
rect 43812 17144 43864 17196
rect 44088 17187 44140 17196
rect 44088 17153 44097 17187
rect 44097 17153 44131 17187
rect 44131 17153 44140 17187
rect 44088 17144 44140 17153
rect 1860 17051 1912 17060
rect 1860 17017 1869 17051
rect 1869 17017 1903 17051
rect 1903 17017 1912 17051
rect 1860 17008 1912 17017
rect 4068 17008 4120 17060
rect 13084 17008 13136 17060
rect 16304 17051 16356 17060
rect 16304 17017 16313 17051
rect 16313 17017 16347 17051
rect 16347 17017 16356 17051
rect 16304 17008 16356 17017
rect 2504 16983 2556 16992
rect 2504 16949 2513 16983
rect 2513 16949 2547 16983
rect 2547 16949 2556 16983
rect 2504 16940 2556 16949
rect 4804 16983 4856 16992
rect 4804 16949 4813 16983
rect 4813 16949 4847 16983
rect 4847 16949 4856 16983
rect 4804 16940 4856 16949
rect 9956 16940 10008 16992
rect 23296 16940 23348 16992
rect 30932 16940 30984 16992
rect 32220 16940 32272 16992
rect 34888 16983 34940 16992
rect 34888 16949 34897 16983
rect 34897 16949 34931 16983
rect 34931 16949 34940 16983
rect 34888 16940 34940 16949
rect 38936 16983 38988 16992
rect 38936 16949 38945 16983
rect 38945 16949 38979 16983
rect 38979 16949 38988 16983
rect 38936 16940 38988 16949
rect 6423 16838 6475 16890
rect 6487 16838 6539 16890
rect 6551 16838 6603 16890
rect 6615 16838 6667 16890
rect 6679 16838 6731 16890
rect 17370 16838 17422 16890
rect 17434 16838 17486 16890
rect 17498 16838 17550 16890
rect 17562 16838 17614 16890
rect 17626 16838 17678 16890
rect 28317 16838 28369 16890
rect 28381 16838 28433 16890
rect 28445 16838 28497 16890
rect 28509 16838 28561 16890
rect 28573 16838 28625 16890
rect 39264 16838 39316 16890
rect 39328 16838 39380 16890
rect 39392 16838 39444 16890
rect 39456 16838 39508 16890
rect 39520 16838 39572 16890
rect 2504 16736 2556 16788
rect 34796 16736 34848 16788
rect 43720 16779 43772 16788
rect 43720 16745 43729 16779
rect 43729 16745 43763 16779
rect 43763 16745 43772 16779
rect 43720 16736 43772 16745
rect 45100 16736 45152 16788
rect 1952 16600 2004 16652
rect 20 16532 72 16584
rect 14188 16532 14240 16584
rect 27620 16532 27672 16584
rect 20720 16396 20772 16448
rect 40684 16396 40736 16448
rect 11896 16294 11948 16346
rect 11960 16294 12012 16346
rect 12024 16294 12076 16346
rect 12088 16294 12140 16346
rect 12152 16294 12204 16346
rect 22843 16294 22895 16346
rect 22907 16294 22959 16346
rect 22971 16294 23023 16346
rect 23035 16294 23087 16346
rect 23099 16294 23151 16346
rect 33790 16294 33842 16346
rect 33854 16294 33906 16346
rect 33918 16294 33970 16346
rect 33982 16294 34034 16346
rect 34046 16294 34098 16346
rect 44737 16294 44789 16346
rect 44801 16294 44853 16346
rect 44865 16294 44917 16346
rect 44929 16294 44981 16346
rect 44993 16294 45045 16346
rect 44088 16192 44140 16244
rect 1032 16056 1084 16108
rect 6828 15852 6880 15904
rect 44364 15895 44416 15904
rect 44364 15861 44373 15895
rect 44373 15861 44407 15895
rect 44407 15861 44416 15895
rect 44364 15852 44416 15861
rect 6423 15750 6475 15802
rect 6487 15750 6539 15802
rect 6551 15750 6603 15802
rect 6615 15750 6667 15802
rect 6679 15750 6731 15802
rect 17370 15750 17422 15802
rect 17434 15750 17486 15802
rect 17498 15750 17550 15802
rect 17562 15750 17614 15802
rect 17626 15750 17678 15802
rect 28317 15750 28369 15802
rect 28381 15750 28433 15802
rect 28445 15750 28497 15802
rect 28509 15750 28561 15802
rect 28573 15750 28625 15802
rect 39264 15750 39316 15802
rect 39328 15750 39380 15802
rect 39392 15750 39444 15802
rect 39456 15750 39508 15802
rect 39520 15750 39572 15802
rect 32956 15648 33008 15700
rect 2964 15444 3016 15496
rect 32680 15376 32732 15428
rect 940 15308 992 15360
rect 31760 15308 31812 15360
rect 32496 15351 32548 15360
rect 32496 15317 32505 15351
rect 32505 15317 32539 15351
rect 32539 15317 32548 15351
rect 32496 15308 32548 15317
rect 11896 15206 11948 15258
rect 11960 15206 12012 15258
rect 12024 15206 12076 15258
rect 12088 15206 12140 15258
rect 12152 15206 12204 15258
rect 22843 15206 22895 15258
rect 22907 15206 22959 15258
rect 22971 15206 23023 15258
rect 23035 15206 23087 15258
rect 23099 15206 23151 15258
rect 33790 15206 33842 15258
rect 33854 15206 33906 15258
rect 33918 15206 33970 15258
rect 33982 15206 34034 15258
rect 34046 15206 34098 15258
rect 44737 15206 44789 15258
rect 44801 15206 44853 15258
rect 44865 15206 44917 15258
rect 44929 15206 44981 15258
rect 44993 15206 45045 15258
rect 23296 15147 23348 15156
rect 23296 15113 23305 15147
rect 23305 15113 23339 15147
rect 23339 15113 23348 15147
rect 23296 15104 23348 15113
rect 34888 15104 34940 15156
rect 18880 15036 18932 15088
rect 26240 15079 26292 15088
rect 26240 15045 26249 15079
rect 26249 15045 26283 15079
rect 26283 15045 26292 15079
rect 26240 15036 26292 15045
rect 32220 15036 32272 15088
rect 33508 15036 33560 15088
rect 18144 14943 18196 14952
rect 18144 14909 18153 14943
rect 18153 14909 18187 14943
rect 18187 14909 18196 14943
rect 18144 14900 18196 14909
rect 20076 14900 20128 14952
rect 32496 14968 32548 15020
rect 26608 14900 26660 14952
rect 18420 14764 18472 14816
rect 31576 14875 31628 14884
rect 31576 14841 31585 14875
rect 31585 14841 31619 14875
rect 31619 14841 31628 14875
rect 31576 14832 31628 14841
rect 31852 14900 31904 14952
rect 32312 14943 32364 14952
rect 32312 14909 32321 14943
rect 32321 14909 32355 14943
rect 32355 14909 32364 14943
rect 32312 14900 32364 14909
rect 32680 14943 32732 14952
rect 32680 14909 32689 14943
rect 32689 14909 32723 14943
rect 32723 14909 32732 14943
rect 32680 14900 32732 14909
rect 32956 14900 33008 14952
rect 33600 15011 33652 15020
rect 33600 14977 33609 15011
rect 33609 14977 33643 15011
rect 33643 14977 33652 15011
rect 33600 14968 33652 14977
rect 33968 15036 34020 15088
rect 37832 15036 37884 15088
rect 32588 14832 32640 14884
rect 20444 14764 20496 14816
rect 22836 14807 22888 14816
rect 22836 14773 22845 14807
rect 22845 14773 22879 14807
rect 22879 14773 22888 14807
rect 22836 14764 22888 14773
rect 25136 14764 25188 14816
rect 31392 14764 31444 14816
rect 32220 14764 32272 14816
rect 34520 14832 34572 14884
rect 36544 15011 36596 15020
rect 36544 14977 36553 15011
rect 36553 14977 36587 15011
rect 36587 14977 36596 15011
rect 36544 14968 36596 14977
rect 36912 14968 36964 15020
rect 32772 14764 32824 14816
rect 33416 14807 33468 14816
rect 33416 14773 33425 14807
rect 33425 14773 33459 14807
rect 33459 14773 33468 14807
rect 33416 14764 33468 14773
rect 34888 14764 34940 14816
rect 36636 14764 36688 14816
rect 37464 14807 37516 14816
rect 37464 14773 37473 14807
rect 37473 14773 37507 14807
rect 37507 14773 37516 14807
rect 37464 14764 37516 14773
rect 37832 14764 37884 14816
rect 38936 14764 38988 14816
rect 6423 14662 6475 14714
rect 6487 14662 6539 14714
rect 6551 14662 6603 14714
rect 6615 14662 6667 14714
rect 6679 14662 6731 14714
rect 17370 14662 17422 14714
rect 17434 14662 17486 14714
rect 17498 14662 17550 14714
rect 17562 14662 17614 14714
rect 17626 14662 17678 14714
rect 28317 14662 28369 14714
rect 28381 14662 28433 14714
rect 28445 14662 28497 14714
rect 28509 14662 28561 14714
rect 28573 14662 28625 14714
rect 39264 14662 39316 14714
rect 39328 14662 39380 14714
rect 39392 14662 39444 14714
rect 39456 14662 39508 14714
rect 39520 14662 39572 14714
rect 1952 14560 2004 14612
rect 18880 14492 18932 14544
rect 18144 14424 18196 14476
rect 27252 14560 27304 14612
rect 30288 14560 30340 14612
rect 32680 14560 32732 14612
rect 33600 14560 33652 14612
rect 42708 14560 42760 14612
rect 36452 14492 36504 14544
rect 9864 14399 9916 14408
rect 9864 14365 9873 14399
rect 9873 14365 9907 14399
rect 9907 14365 9916 14399
rect 9864 14356 9916 14365
rect 9956 14356 10008 14408
rect 13360 14288 13412 14340
rect 18696 14399 18748 14408
rect 18696 14365 18705 14399
rect 18705 14365 18739 14399
rect 18739 14365 18748 14399
rect 32956 14424 33008 14476
rect 18696 14356 18748 14365
rect 22560 14356 22612 14408
rect 29184 14356 29236 14408
rect 31392 14356 31444 14408
rect 33508 14356 33560 14408
rect 34888 14399 34940 14408
rect 34888 14365 34897 14399
rect 34897 14365 34931 14399
rect 34931 14365 34940 14399
rect 34888 14356 34940 14365
rect 35164 14356 35216 14408
rect 36820 14399 36872 14408
rect 36820 14365 36829 14399
rect 36829 14365 36863 14399
rect 36863 14365 36872 14399
rect 36820 14356 36872 14365
rect 37464 14356 37516 14408
rect 40960 14399 41012 14408
rect 40960 14365 40969 14399
rect 40969 14365 41003 14399
rect 41003 14365 41012 14399
rect 40960 14356 41012 14365
rect 11244 14263 11296 14272
rect 11244 14229 11253 14263
rect 11253 14229 11287 14263
rect 11287 14229 11296 14263
rect 11244 14220 11296 14229
rect 11336 14220 11388 14272
rect 14372 14220 14424 14272
rect 18052 14263 18104 14272
rect 18052 14229 18061 14263
rect 18061 14229 18095 14263
rect 18095 14229 18104 14263
rect 18052 14220 18104 14229
rect 20168 14288 20220 14340
rect 20260 14288 20312 14340
rect 18420 14220 18472 14272
rect 19524 14263 19576 14272
rect 19524 14229 19533 14263
rect 19533 14229 19567 14263
rect 19567 14229 19576 14263
rect 19524 14220 19576 14229
rect 26424 14331 26476 14340
rect 26424 14297 26458 14331
rect 26458 14297 26476 14331
rect 26424 14288 26476 14297
rect 26516 14288 26568 14340
rect 32312 14288 32364 14340
rect 22376 14220 22428 14272
rect 22836 14220 22888 14272
rect 27528 14263 27580 14272
rect 27528 14229 27537 14263
rect 27537 14229 27571 14263
rect 27571 14229 27580 14263
rect 27528 14220 27580 14229
rect 32680 14263 32732 14272
rect 32680 14229 32689 14263
rect 32689 14229 32723 14263
rect 32723 14229 32732 14263
rect 32680 14220 32732 14229
rect 33232 14220 33284 14272
rect 36544 14288 36596 14340
rect 36360 14263 36412 14272
rect 36360 14229 36369 14263
rect 36369 14229 36403 14263
rect 36403 14229 36412 14263
rect 36360 14220 36412 14229
rect 40500 14220 40552 14272
rect 42984 14399 43036 14408
rect 42984 14365 42993 14399
rect 42993 14365 43027 14399
rect 43027 14365 43036 14399
rect 42984 14356 43036 14365
rect 41972 14263 42024 14272
rect 41972 14229 41981 14263
rect 41981 14229 42015 14263
rect 42015 14229 42024 14263
rect 41972 14220 42024 14229
rect 44272 14263 44324 14272
rect 44272 14229 44281 14263
rect 44281 14229 44315 14263
rect 44315 14229 44324 14263
rect 44272 14220 44324 14229
rect 11896 14118 11948 14170
rect 11960 14118 12012 14170
rect 12024 14118 12076 14170
rect 12088 14118 12140 14170
rect 12152 14118 12204 14170
rect 22843 14118 22895 14170
rect 22907 14118 22959 14170
rect 22971 14118 23023 14170
rect 23035 14118 23087 14170
rect 23099 14118 23151 14170
rect 33790 14118 33842 14170
rect 33854 14118 33906 14170
rect 33918 14118 33970 14170
rect 33982 14118 34034 14170
rect 34046 14118 34098 14170
rect 44737 14118 44789 14170
rect 44801 14118 44853 14170
rect 44865 14118 44917 14170
rect 44929 14118 44981 14170
rect 44993 14118 45045 14170
rect 6828 14016 6880 14068
rect 5540 13948 5592 14000
rect 5356 13923 5408 13932
rect 5356 13889 5365 13923
rect 5365 13889 5399 13923
rect 5399 13889 5408 13923
rect 5356 13880 5408 13889
rect 6920 13923 6972 13932
rect 6920 13889 6929 13923
rect 6929 13889 6963 13923
rect 6963 13889 6972 13923
rect 16304 14016 16356 14068
rect 17960 14016 18012 14068
rect 20076 14059 20128 14068
rect 20076 14025 20085 14059
rect 20085 14025 20119 14059
rect 20119 14025 20128 14059
rect 20076 14016 20128 14025
rect 20168 14016 20220 14068
rect 14648 13948 14700 14000
rect 6920 13880 6972 13889
rect 13360 13923 13412 13932
rect 13360 13889 13394 13923
rect 13394 13889 13412 13923
rect 13360 13880 13412 13889
rect 17224 13923 17276 13932
rect 17224 13889 17233 13923
rect 17233 13889 17267 13923
rect 17267 13889 17276 13923
rect 17224 13880 17276 13889
rect 18144 13948 18196 14000
rect 19524 13948 19576 14000
rect 20444 13991 20496 14000
rect 20444 13957 20453 13991
rect 20453 13957 20487 13991
rect 20487 13957 20496 13991
rect 20444 13948 20496 13957
rect 25136 14059 25188 14068
rect 25136 14025 25145 14059
rect 25145 14025 25179 14059
rect 25179 14025 25188 14059
rect 25136 14016 25188 14025
rect 20260 13923 20312 13932
rect 20260 13889 20269 13923
rect 20269 13889 20303 13923
rect 20303 13889 20312 13923
rect 20260 13880 20312 13889
rect 20628 13880 20680 13932
rect 21180 13923 21232 13932
rect 21180 13889 21189 13923
rect 21189 13889 21223 13923
rect 21223 13889 21232 13923
rect 21180 13880 21232 13889
rect 22468 13923 22520 13932
rect 22468 13889 22477 13923
rect 22477 13889 22511 13923
rect 22511 13889 22520 13923
rect 22468 13880 22520 13889
rect 22560 13880 22612 13932
rect 27436 14016 27488 14068
rect 27528 14016 27580 14068
rect 31576 14059 31628 14068
rect 31576 14025 31591 14059
rect 31591 14025 31625 14059
rect 31625 14025 31628 14059
rect 31576 14016 31628 14025
rect 33508 14016 33560 14068
rect 34796 14016 34848 14068
rect 36268 14016 36320 14068
rect 36452 14016 36504 14068
rect 36636 14059 36688 14068
rect 36636 14025 36645 14059
rect 36645 14025 36679 14059
rect 36679 14025 36688 14059
rect 36636 14016 36688 14025
rect 36912 14059 36964 14068
rect 36912 14025 36921 14059
rect 36921 14025 36955 14059
rect 36955 14025 36964 14059
rect 36912 14016 36964 14025
rect 37280 14016 37332 14068
rect 940 13812 992 13864
rect 11336 13812 11388 13864
rect 11428 13812 11480 13864
rect 18512 13812 18564 13864
rect 20812 13812 20864 13864
rect 21272 13812 21324 13864
rect 26332 13880 26384 13932
rect 26516 13948 26568 14000
rect 27160 13880 27212 13932
rect 27528 13923 27580 13932
rect 27528 13889 27537 13923
rect 27537 13889 27571 13923
rect 27571 13889 27580 13923
rect 27528 13880 27580 13889
rect 29184 13948 29236 14000
rect 30288 13948 30340 14000
rect 1860 13744 1912 13796
rect 27620 13812 27672 13864
rect 5632 13676 5684 13728
rect 12440 13719 12492 13728
rect 12440 13685 12449 13719
rect 12449 13685 12483 13719
rect 12483 13685 12492 13719
rect 12440 13676 12492 13685
rect 14464 13719 14516 13728
rect 14464 13685 14473 13719
rect 14473 13685 14507 13719
rect 14507 13685 14516 13719
rect 14464 13676 14516 13685
rect 19984 13676 20036 13728
rect 24768 13719 24820 13728
rect 24768 13685 24777 13719
rect 24777 13685 24811 13719
rect 24811 13685 24820 13719
rect 24768 13676 24820 13685
rect 26976 13676 27028 13728
rect 27436 13744 27488 13796
rect 29920 13812 29972 13864
rect 30564 13923 30616 13932
rect 30564 13889 30573 13923
rect 30573 13889 30607 13923
rect 30607 13889 30616 13923
rect 30564 13880 30616 13889
rect 32680 13948 32732 14000
rect 30840 13923 30892 13932
rect 30840 13889 30849 13923
rect 30849 13889 30883 13923
rect 30883 13889 30892 13923
rect 30840 13880 30892 13889
rect 31760 13923 31812 13932
rect 31760 13889 31769 13923
rect 31769 13889 31803 13923
rect 31803 13889 31812 13923
rect 31760 13880 31812 13889
rect 33692 13948 33744 14000
rect 32956 13880 33008 13932
rect 33416 13880 33468 13932
rect 31760 13744 31812 13796
rect 29920 13676 29972 13728
rect 32680 13676 32732 13728
rect 36360 13948 36412 14000
rect 37648 13991 37700 14000
rect 34796 13923 34848 13932
rect 34796 13889 34805 13923
rect 34805 13889 34839 13923
rect 34839 13889 34848 13923
rect 34796 13880 34848 13889
rect 35440 13923 35492 13932
rect 35440 13889 35449 13923
rect 35449 13889 35483 13923
rect 35483 13889 35492 13923
rect 35440 13880 35492 13889
rect 37648 13957 37657 13991
rect 37657 13957 37691 13991
rect 37691 13957 37700 13991
rect 37648 13948 37700 13957
rect 37556 13880 37608 13932
rect 41972 13948 42024 14000
rect 36360 13812 36412 13864
rect 36452 13812 36504 13864
rect 38384 13923 38436 13932
rect 38384 13889 38393 13923
rect 38393 13889 38427 13923
rect 38427 13889 38436 13923
rect 38384 13880 38436 13889
rect 38936 13812 38988 13864
rect 36084 13744 36136 13796
rect 36820 13744 36872 13796
rect 40592 13744 40644 13796
rect 36636 13676 36688 13728
rect 37464 13719 37516 13728
rect 37464 13685 37473 13719
rect 37473 13685 37507 13719
rect 37507 13685 37516 13719
rect 37464 13676 37516 13685
rect 42064 13719 42116 13728
rect 42064 13685 42073 13719
rect 42073 13685 42107 13719
rect 42107 13685 42116 13719
rect 42064 13676 42116 13685
rect 6423 13574 6475 13626
rect 6487 13574 6539 13626
rect 6551 13574 6603 13626
rect 6615 13574 6667 13626
rect 6679 13574 6731 13626
rect 17370 13574 17422 13626
rect 17434 13574 17486 13626
rect 17498 13574 17550 13626
rect 17562 13574 17614 13626
rect 17626 13574 17678 13626
rect 28317 13574 28369 13626
rect 28381 13574 28433 13626
rect 28445 13574 28497 13626
rect 28509 13574 28561 13626
rect 28573 13574 28625 13626
rect 39264 13574 39316 13626
rect 39328 13574 39380 13626
rect 39392 13574 39444 13626
rect 39456 13574 39508 13626
rect 39520 13574 39572 13626
rect 14648 13515 14700 13524
rect 14648 13481 14657 13515
rect 14657 13481 14691 13515
rect 14691 13481 14700 13515
rect 14648 13472 14700 13481
rect 18512 13472 18564 13524
rect 20444 13472 20496 13524
rect 8576 13404 8628 13456
rect 20260 13404 20312 13456
rect 21180 13472 21232 13524
rect 26332 13515 26384 13524
rect 26332 13481 26341 13515
rect 26341 13481 26375 13515
rect 26375 13481 26384 13515
rect 26332 13472 26384 13481
rect 26424 13472 26476 13524
rect 30840 13472 30892 13524
rect 32128 13515 32180 13524
rect 32128 13481 32137 13515
rect 32137 13481 32171 13515
rect 32171 13481 32180 13515
rect 32128 13472 32180 13481
rect 33416 13472 33468 13524
rect 37280 13472 37332 13524
rect 42708 13472 42760 13524
rect 5080 13311 5132 13320
rect 5080 13277 5089 13311
rect 5089 13277 5123 13311
rect 5123 13277 5132 13311
rect 5080 13268 5132 13277
rect 7564 13379 7616 13388
rect 7564 13345 7573 13379
rect 7573 13345 7607 13379
rect 7607 13345 7616 13379
rect 7564 13336 7616 13345
rect 11060 13336 11112 13388
rect 11428 13379 11480 13388
rect 11428 13345 11437 13379
rect 11437 13345 11471 13379
rect 11471 13345 11480 13379
rect 11428 13336 11480 13345
rect 18144 13336 18196 13388
rect 20720 13379 20772 13388
rect 20720 13345 20729 13379
rect 20729 13345 20763 13379
rect 20763 13345 20772 13379
rect 20720 13336 20772 13345
rect 5632 13268 5684 13320
rect 11244 13268 11296 13320
rect 14372 13311 14424 13320
rect 14372 13277 14381 13311
rect 14381 13277 14415 13311
rect 14415 13277 14424 13311
rect 14372 13268 14424 13277
rect 14464 13311 14516 13320
rect 14464 13277 14473 13311
rect 14473 13277 14507 13311
rect 14507 13277 14516 13311
rect 14464 13268 14516 13277
rect 11796 13200 11848 13252
rect 7380 13175 7432 13184
rect 7380 13141 7389 13175
rect 7389 13141 7423 13175
rect 7423 13141 7432 13175
rect 7380 13132 7432 13141
rect 10324 13132 10376 13184
rect 11704 13132 11756 13184
rect 12808 13175 12860 13184
rect 12808 13141 12817 13175
rect 12817 13141 12851 13175
rect 12851 13141 12860 13175
rect 12808 13132 12860 13141
rect 17960 13200 18012 13252
rect 19984 13311 20036 13320
rect 19984 13277 19993 13311
rect 19993 13277 20027 13311
rect 20027 13277 20036 13311
rect 19984 13268 20036 13277
rect 20628 13268 20680 13320
rect 21548 13336 21600 13388
rect 22008 13336 22060 13388
rect 21456 13311 21508 13320
rect 21456 13277 21465 13311
rect 21465 13277 21499 13311
rect 21499 13277 21508 13311
rect 21456 13268 21508 13277
rect 22284 13268 22336 13320
rect 30288 13404 30340 13456
rect 22652 13336 22704 13388
rect 26332 13336 26384 13388
rect 30564 13404 30616 13456
rect 31484 13404 31536 13456
rect 31760 13404 31812 13456
rect 32404 13404 32456 13456
rect 24584 13311 24636 13320
rect 24584 13277 24593 13311
rect 24593 13277 24627 13311
rect 24627 13277 24636 13311
rect 24584 13268 24636 13277
rect 26976 13311 27028 13320
rect 26976 13277 26985 13311
rect 26985 13277 27019 13311
rect 27019 13277 27028 13311
rect 26976 13268 27028 13277
rect 27160 13268 27212 13320
rect 28908 13311 28960 13320
rect 28908 13277 28917 13311
rect 28917 13277 28951 13311
rect 28951 13277 28960 13311
rect 28908 13268 28960 13277
rect 29920 13311 29972 13320
rect 29920 13277 29929 13311
rect 29929 13277 29963 13311
rect 29963 13277 29972 13311
rect 29920 13268 29972 13277
rect 30932 13379 30984 13388
rect 30932 13345 30941 13379
rect 30941 13345 30975 13379
rect 30975 13345 30984 13379
rect 30932 13336 30984 13345
rect 30564 13268 30616 13320
rect 32680 13311 32732 13320
rect 32680 13277 32688 13311
rect 32688 13277 32722 13311
rect 32722 13277 32732 13311
rect 32680 13268 32732 13277
rect 32772 13311 32824 13320
rect 32772 13277 32781 13311
rect 32781 13277 32815 13311
rect 32815 13277 32824 13311
rect 32772 13268 32824 13277
rect 33140 13268 33192 13320
rect 36084 13379 36136 13388
rect 36084 13345 36093 13379
rect 36093 13345 36127 13379
rect 36127 13345 36136 13379
rect 36084 13336 36136 13345
rect 36820 13336 36872 13388
rect 18052 13132 18104 13184
rect 20720 13200 20772 13252
rect 22652 13200 22704 13252
rect 20996 13175 21048 13184
rect 20996 13141 21005 13175
rect 21005 13141 21039 13175
rect 21039 13141 21048 13175
rect 20996 13132 21048 13141
rect 26884 13200 26936 13252
rect 30932 13200 30984 13252
rect 31852 13200 31904 13252
rect 32404 13243 32456 13252
rect 32404 13209 32413 13243
rect 32413 13209 32447 13243
rect 32447 13209 32456 13243
rect 32404 13200 32456 13209
rect 32496 13243 32548 13252
rect 32496 13209 32505 13243
rect 32505 13209 32539 13243
rect 32539 13209 32548 13243
rect 32496 13200 32548 13209
rect 35716 13200 35768 13252
rect 36268 13311 36320 13320
rect 36268 13277 36277 13311
rect 36277 13277 36311 13311
rect 36311 13277 36320 13311
rect 36268 13268 36320 13277
rect 37464 13268 37516 13320
rect 40500 13311 40552 13320
rect 40500 13277 40509 13311
rect 40509 13277 40543 13311
rect 40543 13277 40552 13311
rect 40500 13268 40552 13277
rect 40592 13268 40644 13320
rect 41972 13336 42024 13388
rect 42064 13268 42116 13320
rect 40132 13200 40184 13252
rect 41052 13200 41104 13252
rect 41696 13200 41748 13252
rect 32680 13132 32732 13184
rect 36452 13175 36504 13184
rect 36452 13141 36461 13175
rect 36461 13141 36495 13175
rect 36495 13141 36504 13175
rect 36452 13132 36504 13141
rect 38384 13132 38436 13184
rect 38660 13132 38712 13184
rect 40408 13175 40460 13184
rect 40408 13141 40417 13175
rect 40417 13141 40451 13175
rect 40451 13141 40460 13175
rect 40408 13132 40460 13141
rect 42340 13175 42392 13184
rect 42340 13141 42349 13175
rect 42349 13141 42383 13175
rect 42383 13141 42392 13175
rect 42340 13132 42392 13141
rect 11896 13030 11948 13082
rect 11960 13030 12012 13082
rect 12024 13030 12076 13082
rect 12088 13030 12140 13082
rect 12152 13030 12204 13082
rect 22843 13030 22895 13082
rect 22907 13030 22959 13082
rect 22971 13030 23023 13082
rect 23035 13030 23087 13082
rect 23099 13030 23151 13082
rect 33790 13030 33842 13082
rect 33854 13030 33906 13082
rect 33918 13030 33970 13082
rect 33982 13030 34034 13082
rect 34046 13030 34098 13082
rect 44737 13030 44789 13082
rect 44801 13030 44853 13082
rect 44865 13030 44917 13082
rect 44929 13030 44981 13082
rect 44993 13030 45045 13082
rect 5356 12928 5408 12980
rect 11704 12971 11756 12980
rect 11704 12937 11713 12971
rect 11713 12937 11747 12971
rect 11747 12937 11756 12971
rect 11704 12928 11756 12937
rect 14556 12971 14608 12980
rect 14556 12937 14565 12971
rect 14565 12937 14599 12971
rect 14599 12937 14608 12971
rect 14556 12928 14608 12937
rect 3148 12835 3200 12844
rect 3148 12801 3157 12835
rect 3157 12801 3191 12835
rect 3191 12801 3200 12835
rect 3148 12792 3200 12801
rect 3976 12792 4028 12844
rect 4344 12835 4396 12844
rect 4344 12801 4378 12835
rect 4378 12801 4396 12835
rect 4344 12792 4396 12801
rect 4804 12792 4856 12844
rect 5080 12724 5132 12776
rect 8576 12835 8628 12844
rect 8576 12801 8585 12835
rect 8585 12801 8619 12835
rect 8619 12801 8628 12835
rect 8576 12792 8628 12801
rect 9864 12860 9916 12912
rect 11428 12860 11480 12912
rect 20812 12928 20864 12980
rect 10048 12835 10100 12844
rect 10048 12801 10082 12835
rect 10082 12801 10100 12835
rect 10048 12792 10100 12801
rect 11152 12792 11204 12844
rect 13820 12792 13872 12844
rect 17224 12792 17276 12844
rect 12348 12767 12400 12776
rect 12348 12733 12357 12767
rect 12357 12733 12391 12767
rect 12391 12733 12400 12767
rect 12348 12724 12400 12733
rect 13176 12767 13228 12776
rect 13176 12733 13185 12767
rect 13185 12733 13219 12767
rect 13219 12733 13228 12767
rect 13176 12724 13228 12733
rect 18144 12792 18196 12844
rect 18512 12835 18564 12844
rect 18512 12801 18521 12835
rect 18521 12801 18555 12835
rect 18555 12801 18564 12835
rect 18512 12792 18564 12801
rect 20904 12835 20956 12844
rect 20904 12801 20913 12835
rect 20913 12801 20947 12835
rect 20947 12801 20956 12835
rect 20904 12792 20956 12801
rect 22192 12928 22244 12980
rect 22468 12928 22520 12980
rect 27160 12928 27212 12980
rect 31944 12928 31996 12980
rect 33048 12928 33100 12980
rect 21088 12835 21140 12844
rect 21088 12801 21097 12835
rect 21097 12801 21131 12835
rect 21131 12801 21140 12835
rect 21088 12792 21140 12801
rect 17960 12724 18012 12776
rect 20812 12724 20864 12776
rect 22008 12835 22060 12844
rect 22008 12801 22017 12835
rect 22017 12801 22051 12835
rect 22051 12801 22060 12835
rect 22008 12792 22060 12801
rect 25228 12792 25280 12844
rect 25964 12792 26016 12844
rect 29184 12835 29236 12844
rect 29184 12801 29193 12835
rect 29193 12801 29227 12835
rect 29227 12801 29236 12835
rect 29184 12792 29236 12801
rect 29460 12835 29512 12844
rect 29460 12801 29494 12835
rect 29494 12801 29512 12835
rect 29460 12792 29512 12801
rect 2780 12588 2832 12640
rect 7748 12588 7800 12640
rect 11152 12631 11204 12640
rect 11152 12597 11161 12631
rect 11161 12597 11195 12631
rect 11195 12597 11204 12631
rect 11152 12588 11204 12597
rect 14096 12588 14148 12640
rect 14372 12588 14424 12640
rect 21272 12656 21324 12708
rect 20628 12588 20680 12640
rect 21456 12724 21508 12776
rect 21548 12656 21600 12708
rect 22192 12724 22244 12776
rect 24676 12724 24728 12776
rect 31484 12903 31536 12912
rect 31484 12869 31493 12903
rect 31493 12869 31527 12903
rect 31527 12869 31536 12903
rect 31484 12860 31536 12869
rect 33232 12860 33284 12912
rect 33416 12903 33468 12912
rect 33416 12869 33425 12903
rect 33425 12869 33459 12903
rect 33459 12869 33468 12903
rect 33416 12860 33468 12869
rect 31576 12835 31628 12844
rect 31576 12801 31585 12835
rect 31585 12801 31619 12835
rect 31619 12801 31628 12835
rect 31576 12792 31628 12801
rect 32588 12792 32640 12844
rect 32680 12835 32732 12844
rect 32680 12801 32689 12835
rect 32689 12801 32723 12835
rect 32723 12801 32732 12835
rect 32680 12792 32732 12801
rect 37556 12928 37608 12980
rect 36176 12860 36228 12912
rect 36360 12860 36412 12912
rect 40040 12928 40092 12980
rect 40316 12928 40368 12980
rect 40500 12928 40552 12980
rect 41052 12928 41104 12980
rect 35624 12835 35676 12844
rect 35624 12801 35633 12835
rect 35633 12801 35667 12835
rect 35667 12801 35676 12835
rect 35624 12792 35676 12801
rect 35716 12792 35768 12844
rect 36268 12835 36320 12844
rect 36268 12801 36277 12835
rect 36277 12801 36311 12835
rect 36311 12801 36320 12835
rect 36268 12792 36320 12801
rect 36452 12835 36504 12844
rect 36452 12801 36461 12835
rect 36461 12801 36495 12835
rect 36495 12801 36504 12835
rect 36452 12792 36504 12801
rect 36636 12835 36688 12844
rect 36636 12801 36645 12835
rect 36645 12801 36679 12835
rect 36679 12801 36688 12835
rect 36636 12792 36688 12801
rect 37648 12835 37700 12844
rect 37648 12801 37657 12835
rect 37657 12801 37691 12835
rect 37691 12801 37700 12835
rect 37648 12792 37700 12801
rect 32496 12724 32548 12776
rect 22284 12656 22336 12708
rect 23112 12656 23164 12708
rect 32128 12656 32180 12708
rect 33508 12656 33560 12708
rect 22100 12588 22152 12640
rect 22652 12588 22704 12640
rect 30564 12631 30616 12640
rect 30564 12597 30573 12631
rect 30573 12597 30607 12631
rect 30607 12597 30616 12631
rect 30564 12588 30616 12597
rect 31944 12588 31996 12640
rect 36084 12656 36136 12708
rect 37924 12835 37976 12844
rect 37924 12801 37933 12835
rect 37933 12801 37967 12835
rect 37967 12801 37976 12835
rect 37924 12792 37976 12801
rect 38660 12792 38712 12844
rect 39764 12860 39816 12912
rect 42064 12928 42116 12980
rect 39396 12767 39448 12776
rect 39396 12733 39405 12767
rect 39405 12733 39439 12767
rect 39439 12733 39448 12767
rect 39396 12724 39448 12733
rect 37372 12588 37424 12640
rect 38568 12656 38620 12708
rect 40132 12724 40184 12776
rect 41512 12835 41564 12844
rect 41512 12801 41521 12835
rect 41521 12801 41555 12835
rect 41555 12801 41564 12835
rect 41512 12792 41564 12801
rect 42340 12792 42392 12844
rect 40132 12588 40184 12640
rect 40960 12588 41012 12640
rect 41696 12724 41748 12776
rect 41880 12767 41932 12776
rect 41880 12733 41889 12767
rect 41889 12733 41923 12767
rect 41923 12733 41932 12767
rect 41880 12724 41932 12733
rect 41604 12588 41656 12640
rect 45008 12588 45060 12640
rect 6423 12486 6475 12538
rect 6487 12486 6539 12538
rect 6551 12486 6603 12538
rect 6615 12486 6667 12538
rect 6679 12486 6731 12538
rect 17370 12486 17422 12538
rect 17434 12486 17486 12538
rect 17498 12486 17550 12538
rect 17562 12486 17614 12538
rect 17626 12486 17678 12538
rect 28317 12486 28369 12538
rect 28381 12486 28433 12538
rect 28445 12486 28497 12538
rect 28509 12486 28561 12538
rect 28573 12486 28625 12538
rect 39264 12486 39316 12538
rect 39328 12486 39380 12538
rect 39392 12486 39444 12538
rect 39456 12486 39508 12538
rect 39520 12486 39572 12538
rect 2964 12427 3016 12436
rect 2964 12393 2973 12427
rect 2973 12393 3007 12427
rect 3007 12393 3016 12427
rect 2964 12384 3016 12393
rect 7380 12427 7432 12436
rect 7380 12393 7389 12427
rect 7389 12393 7423 12427
rect 7423 12393 7432 12427
rect 7380 12384 7432 12393
rect 10048 12384 10100 12436
rect 11060 12384 11112 12436
rect 11796 12384 11848 12436
rect 13820 12384 13872 12436
rect 20720 12384 20772 12436
rect 21916 12384 21968 12436
rect 3424 12180 3476 12232
rect 5080 12180 5132 12232
rect 9680 12248 9732 12300
rect 12348 12316 12400 12368
rect 20904 12316 20956 12368
rect 7564 12180 7616 12232
rect 7748 12223 7800 12232
rect 7748 12189 7757 12223
rect 7757 12189 7791 12223
rect 7791 12189 7800 12223
rect 7748 12180 7800 12189
rect 10324 12223 10376 12232
rect 10324 12189 10333 12223
rect 10333 12189 10367 12223
rect 10367 12189 10376 12223
rect 10324 12180 10376 12189
rect 11428 12180 11480 12232
rect 14556 12180 14608 12232
rect 17224 12248 17276 12300
rect 18512 12248 18564 12300
rect 17500 12180 17552 12232
rect 17960 12180 18012 12232
rect 18696 12223 18748 12232
rect 18696 12189 18705 12223
rect 18705 12189 18739 12223
rect 18739 12189 18748 12223
rect 18696 12180 18748 12189
rect 21824 12223 21876 12232
rect 21824 12189 21833 12223
rect 21833 12189 21867 12223
rect 21867 12189 21876 12223
rect 21824 12180 21876 12189
rect 22100 12248 22152 12300
rect 25872 12384 25924 12436
rect 26884 12427 26936 12436
rect 26884 12393 26893 12427
rect 26893 12393 26927 12427
rect 26927 12393 26936 12427
rect 26884 12384 26936 12393
rect 31208 12384 31260 12436
rect 33324 12384 33376 12436
rect 35348 12384 35400 12436
rect 35532 12384 35584 12436
rect 29552 12316 29604 12368
rect 31760 12316 31812 12368
rect 24584 12291 24636 12300
rect 24584 12257 24593 12291
rect 24593 12257 24627 12291
rect 24627 12257 24636 12291
rect 24584 12248 24636 12257
rect 24860 12248 24912 12300
rect 26516 12248 26568 12300
rect 28908 12248 28960 12300
rect 32128 12248 32180 12300
rect 6000 12112 6052 12164
rect 4252 12087 4304 12096
rect 4252 12053 4261 12087
rect 4261 12053 4295 12087
rect 4295 12053 4304 12087
rect 4252 12044 4304 12053
rect 4620 12087 4672 12096
rect 4620 12053 4629 12087
rect 4629 12053 4663 12087
rect 4663 12053 4672 12087
rect 4620 12044 4672 12053
rect 8208 12112 8260 12164
rect 12440 12112 12492 12164
rect 7380 12044 7432 12096
rect 11152 12044 11204 12096
rect 13360 12087 13412 12096
rect 13360 12053 13369 12087
rect 13369 12053 13403 12087
rect 13403 12053 13412 12087
rect 13360 12044 13412 12053
rect 17132 12044 17184 12096
rect 21916 12155 21968 12164
rect 21916 12121 21925 12155
rect 21925 12121 21959 12155
rect 21959 12121 21968 12155
rect 21916 12112 21968 12121
rect 22100 12155 22152 12164
rect 22100 12121 22135 12155
rect 22135 12121 22152 12155
rect 23112 12223 23164 12232
rect 23112 12189 23121 12223
rect 23121 12189 23155 12223
rect 23155 12189 23164 12223
rect 23112 12180 23164 12189
rect 26148 12180 26200 12232
rect 29736 12223 29788 12232
rect 29736 12189 29745 12223
rect 29745 12189 29779 12223
rect 29779 12189 29788 12223
rect 29736 12180 29788 12189
rect 22100 12112 22152 12121
rect 21456 12044 21508 12096
rect 22744 12044 22796 12096
rect 25504 12112 25556 12164
rect 29644 12112 29696 12164
rect 30932 12112 30984 12164
rect 25136 12044 25188 12096
rect 31208 12087 31260 12096
rect 31208 12053 31217 12087
rect 31217 12053 31251 12087
rect 31251 12053 31260 12087
rect 31208 12044 31260 12053
rect 31760 12223 31812 12232
rect 31760 12189 31769 12223
rect 31769 12189 31803 12223
rect 31803 12189 31812 12223
rect 31760 12180 31812 12189
rect 31944 12223 31996 12232
rect 31944 12189 31953 12223
rect 31953 12189 31987 12223
rect 31987 12189 31996 12223
rect 31944 12180 31996 12189
rect 33048 12316 33100 12368
rect 35256 12316 35308 12368
rect 35808 12316 35860 12368
rect 32496 12248 32548 12300
rect 32128 12155 32180 12164
rect 32128 12121 32137 12155
rect 32137 12121 32171 12155
rect 32171 12121 32180 12155
rect 32128 12112 32180 12121
rect 33232 12180 33284 12232
rect 35992 12248 36044 12300
rect 36268 12384 36320 12436
rect 37924 12384 37976 12436
rect 38016 12316 38068 12368
rect 38660 12316 38712 12368
rect 39212 12316 39264 12368
rect 40224 12316 40276 12368
rect 32772 12155 32824 12164
rect 32772 12121 32781 12155
rect 32781 12121 32815 12155
rect 32815 12121 32824 12155
rect 32772 12112 32824 12121
rect 35256 12155 35308 12164
rect 35256 12121 35265 12155
rect 35265 12121 35299 12155
rect 35299 12121 35308 12155
rect 35256 12112 35308 12121
rect 35716 12112 35768 12164
rect 33140 12087 33192 12096
rect 33140 12053 33149 12087
rect 33149 12053 33183 12087
rect 33183 12053 33192 12087
rect 33140 12044 33192 12053
rect 35164 12044 35216 12096
rect 35624 12087 35676 12096
rect 35624 12053 35633 12087
rect 35633 12053 35667 12087
rect 35667 12053 35676 12087
rect 35624 12044 35676 12053
rect 36176 12180 36228 12232
rect 36636 12180 36688 12232
rect 37280 12223 37332 12232
rect 37280 12189 37289 12223
rect 37289 12189 37323 12223
rect 37323 12189 37332 12223
rect 37280 12180 37332 12189
rect 37372 12223 37424 12232
rect 37372 12189 37381 12223
rect 37381 12189 37415 12223
rect 37415 12189 37424 12223
rect 37372 12180 37424 12189
rect 37924 12180 37976 12232
rect 37740 12112 37792 12164
rect 38108 12180 38160 12232
rect 38752 12180 38804 12232
rect 40040 12248 40092 12300
rect 40408 12248 40460 12300
rect 38660 12112 38712 12164
rect 39120 12223 39172 12232
rect 39120 12189 39129 12223
rect 39129 12189 39163 12223
rect 39163 12189 39172 12223
rect 39120 12180 39172 12189
rect 39212 12223 39264 12232
rect 39212 12189 39221 12223
rect 39221 12189 39255 12223
rect 39255 12189 39264 12223
rect 39212 12180 39264 12189
rect 41696 12248 41748 12300
rect 39028 12112 39080 12164
rect 38108 12044 38160 12096
rect 38384 12087 38436 12096
rect 38384 12053 38393 12087
rect 38393 12053 38427 12087
rect 38427 12053 38436 12087
rect 38384 12044 38436 12053
rect 38844 12087 38896 12096
rect 38844 12053 38853 12087
rect 38853 12053 38887 12087
rect 38887 12053 38896 12087
rect 38844 12044 38896 12053
rect 39120 12044 39172 12096
rect 40316 12112 40368 12164
rect 41420 12180 41472 12232
rect 41972 12180 42024 12232
rect 42248 12223 42300 12232
rect 42248 12189 42257 12223
rect 42257 12189 42291 12223
rect 42291 12189 42300 12223
rect 42248 12180 42300 12189
rect 41512 12112 41564 12164
rect 40868 12087 40920 12096
rect 40868 12053 40877 12087
rect 40877 12053 40911 12087
rect 40911 12053 40920 12087
rect 40868 12044 40920 12053
rect 41696 12044 41748 12096
rect 11896 11942 11948 11994
rect 11960 11942 12012 11994
rect 12024 11942 12076 11994
rect 12088 11942 12140 11994
rect 12152 11942 12204 11994
rect 22843 11942 22895 11994
rect 22907 11942 22959 11994
rect 22971 11942 23023 11994
rect 23035 11942 23087 11994
rect 23099 11942 23151 11994
rect 33790 11942 33842 11994
rect 33854 11942 33906 11994
rect 33918 11942 33970 11994
rect 33982 11942 34034 11994
rect 34046 11942 34098 11994
rect 44737 11942 44789 11994
rect 44801 11942 44853 11994
rect 44865 11942 44917 11994
rect 44929 11942 44981 11994
rect 44993 11942 45045 11994
rect 4528 11772 4580 11824
rect 4252 11704 4304 11756
rect 5080 11772 5132 11824
rect 7380 11883 7432 11892
rect 7380 11849 7389 11883
rect 7389 11849 7423 11883
rect 7423 11849 7432 11883
rect 7380 11840 7432 11849
rect 7748 11840 7800 11892
rect 8208 11883 8260 11892
rect 8208 11849 8217 11883
rect 8217 11849 8251 11883
rect 8251 11849 8260 11883
rect 8208 11840 8260 11849
rect 13360 11840 13412 11892
rect 10784 11772 10836 11824
rect 10324 11747 10376 11756
rect 10324 11713 10333 11747
rect 10333 11713 10367 11747
rect 10367 11713 10376 11747
rect 10324 11704 10376 11713
rect 12900 11704 12952 11756
rect 13176 11747 13228 11756
rect 13176 11713 13185 11747
rect 13185 11713 13219 11747
rect 13219 11713 13228 11747
rect 13176 11704 13228 11713
rect 14648 11704 14700 11756
rect 16396 11704 16448 11756
rect 19984 11840 20036 11892
rect 22744 11840 22796 11892
rect 25872 11840 25924 11892
rect 29460 11840 29512 11892
rect 29736 11840 29788 11892
rect 33508 11883 33560 11892
rect 33508 11849 33517 11883
rect 33517 11849 33551 11883
rect 33551 11849 33560 11883
rect 33508 11840 33560 11849
rect 35440 11840 35492 11892
rect 36544 11840 36596 11892
rect 36636 11840 36688 11892
rect 37556 11840 37608 11892
rect 37648 11840 37700 11892
rect 38108 11883 38160 11892
rect 38108 11849 38117 11883
rect 38117 11849 38151 11883
rect 38151 11849 38160 11883
rect 38108 11840 38160 11849
rect 38568 11883 38620 11892
rect 38568 11849 38577 11883
rect 38577 11849 38611 11883
rect 38611 11849 38620 11883
rect 38568 11840 38620 11849
rect 38936 11883 38988 11892
rect 38936 11849 38945 11883
rect 38945 11849 38979 11883
rect 38979 11849 38988 11883
rect 38936 11840 38988 11849
rect 41420 11883 41472 11892
rect 41420 11849 41429 11883
rect 41429 11849 41463 11883
rect 41463 11849 41472 11883
rect 41420 11840 41472 11849
rect 21916 11772 21968 11824
rect 20996 11704 21048 11756
rect 21456 11747 21508 11756
rect 21456 11713 21465 11747
rect 21465 11713 21499 11747
rect 21499 11713 21508 11747
rect 21456 11704 21508 11713
rect 22100 11747 22152 11756
rect 22100 11713 22109 11747
rect 22109 11713 22143 11747
rect 22143 11713 22152 11747
rect 22100 11704 22152 11713
rect 22284 11704 22336 11756
rect 22836 11747 22888 11756
rect 22836 11713 22845 11747
rect 22845 11713 22879 11747
rect 22879 11713 22888 11747
rect 22836 11704 22888 11713
rect 25044 11772 25096 11824
rect 25136 11815 25188 11824
rect 25136 11781 25145 11815
rect 25145 11781 25179 11815
rect 25179 11781 25188 11815
rect 25136 11772 25188 11781
rect 26148 11704 26200 11756
rect 9680 11636 9732 11688
rect 10876 11636 10928 11688
rect 17040 11636 17092 11688
rect 17500 11679 17552 11688
rect 17500 11645 17509 11679
rect 17509 11645 17543 11679
rect 17543 11645 17552 11679
rect 17500 11636 17552 11645
rect 20260 11679 20312 11688
rect 20260 11645 20269 11679
rect 20269 11645 20303 11679
rect 20303 11645 20312 11679
rect 20260 11636 20312 11645
rect 20628 11636 20680 11688
rect 24860 11679 24912 11688
rect 24860 11645 24869 11679
rect 24869 11645 24903 11679
rect 24903 11645 24912 11679
rect 24860 11636 24912 11645
rect 4160 11568 4212 11620
rect 24768 11568 24820 11620
rect 29552 11747 29604 11756
rect 29552 11713 29561 11747
rect 29561 11713 29595 11747
rect 29595 11713 29604 11747
rect 29552 11704 29604 11713
rect 29644 11636 29696 11688
rect 30656 11772 30708 11824
rect 31208 11772 31260 11824
rect 32128 11772 32180 11824
rect 31852 11704 31904 11756
rect 31944 11704 31996 11756
rect 32772 11772 32824 11824
rect 35624 11772 35676 11824
rect 35716 11772 35768 11824
rect 35256 11704 35308 11756
rect 35808 11747 35860 11756
rect 35808 11713 35817 11747
rect 35817 11713 35851 11747
rect 35851 11713 35860 11747
rect 35808 11704 35860 11713
rect 36084 11704 36136 11756
rect 36636 11747 36688 11756
rect 36636 11713 36645 11747
rect 36645 11713 36679 11747
rect 36679 11713 36688 11747
rect 36636 11704 36688 11713
rect 37740 11815 37792 11824
rect 37740 11781 37749 11815
rect 37749 11781 37783 11815
rect 37783 11781 37792 11815
rect 37740 11772 37792 11781
rect 40868 11772 40920 11824
rect 41788 11815 41840 11824
rect 41788 11781 41797 11815
rect 41797 11781 41831 11815
rect 41831 11781 41840 11815
rect 41788 11772 41840 11781
rect 42248 11772 42300 11824
rect 42800 11772 42852 11824
rect 38384 11704 38436 11756
rect 38844 11747 38896 11756
rect 38844 11713 38853 11747
rect 38853 11713 38887 11747
rect 38887 11713 38896 11747
rect 38844 11704 38896 11713
rect 30288 11679 30340 11688
rect 30288 11645 30297 11679
rect 30297 11645 30331 11679
rect 30331 11645 30340 11679
rect 30288 11636 30340 11645
rect 31760 11636 31812 11688
rect 33508 11636 33560 11688
rect 33692 11636 33744 11688
rect 3976 11500 4028 11552
rect 4068 11500 4120 11552
rect 5632 11500 5684 11552
rect 7196 11500 7248 11552
rect 10232 11500 10284 11552
rect 16856 11543 16908 11552
rect 16856 11509 16865 11543
rect 16865 11509 16899 11543
rect 16899 11509 16908 11543
rect 16856 11500 16908 11509
rect 19708 11500 19760 11552
rect 20996 11543 21048 11552
rect 20996 11509 21005 11543
rect 21005 11509 21039 11543
rect 21039 11509 21048 11543
rect 20996 11500 21048 11509
rect 22652 11500 22704 11552
rect 29644 11500 29696 11552
rect 35992 11636 36044 11688
rect 36544 11568 36596 11620
rect 37556 11636 37608 11688
rect 38108 11636 38160 11688
rect 39212 11679 39264 11688
rect 39212 11645 39221 11679
rect 39221 11645 39255 11679
rect 39255 11645 39264 11679
rect 39212 11636 39264 11645
rect 41512 11704 41564 11756
rect 41604 11747 41656 11756
rect 41604 11713 41613 11747
rect 41613 11713 41647 11747
rect 41647 11713 41656 11747
rect 41604 11704 41656 11713
rect 41972 11704 42024 11756
rect 37648 11568 37700 11620
rect 38292 11568 38344 11620
rect 43168 11636 43220 11688
rect 40040 11568 40092 11620
rect 31760 11500 31812 11552
rect 32772 11500 32824 11552
rect 33324 11543 33376 11552
rect 33324 11509 33333 11543
rect 33333 11509 33367 11543
rect 33367 11509 33376 11543
rect 33324 11500 33376 11509
rect 35900 11543 35952 11552
rect 35900 11509 35909 11543
rect 35909 11509 35943 11543
rect 35943 11509 35952 11543
rect 35900 11500 35952 11509
rect 36728 11543 36780 11552
rect 36728 11509 36737 11543
rect 36737 11509 36771 11543
rect 36771 11509 36780 11543
rect 36728 11500 36780 11509
rect 37556 11500 37608 11552
rect 6423 11398 6475 11450
rect 6487 11398 6539 11450
rect 6551 11398 6603 11450
rect 6615 11398 6667 11450
rect 6679 11398 6731 11450
rect 17370 11398 17422 11450
rect 17434 11398 17486 11450
rect 17498 11398 17550 11450
rect 17562 11398 17614 11450
rect 17626 11398 17678 11450
rect 28317 11398 28369 11450
rect 28381 11398 28433 11450
rect 28445 11398 28497 11450
rect 28509 11398 28561 11450
rect 28573 11398 28625 11450
rect 39264 11398 39316 11450
rect 39328 11398 39380 11450
rect 39392 11398 39444 11450
rect 39456 11398 39508 11450
rect 39520 11398 39572 11450
rect 3424 11339 3476 11348
rect 3424 11305 3433 11339
rect 3433 11305 3467 11339
rect 3467 11305 3476 11339
rect 3424 11296 3476 11305
rect 5540 11339 5592 11348
rect 5540 11305 5549 11339
rect 5549 11305 5583 11339
rect 5583 11305 5592 11339
rect 5540 11296 5592 11305
rect 6000 11339 6052 11348
rect 6000 11305 6009 11339
rect 6009 11305 6043 11339
rect 6043 11305 6052 11339
rect 6000 11296 6052 11305
rect 3976 11160 4028 11212
rect 3148 11135 3200 11144
rect 3148 11101 3157 11135
rect 3157 11101 3191 11135
rect 3191 11101 3200 11135
rect 3148 11092 3200 11101
rect 3240 11135 3292 11144
rect 3240 11101 3249 11135
rect 3249 11101 3283 11135
rect 3283 11101 3292 11135
rect 3240 11092 3292 11101
rect 4160 11135 4212 11144
rect 4160 11101 4169 11135
rect 4169 11101 4203 11135
rect 4203 11101 4212 11135
rect 4160 11092 4212 11101
rect 7196 11203 7248 11212
rect 7196 11169 7205 11203
rect 7205 11169 7239 11203
rect 7239 11169 7248 11203
rect 7196 11160 7248 11169
rect 7564 11160 7616 11212
rect 9864 11160 9916 11212
rect 11428 11160 11480 11212
rect 7932 11135 7984 11144
rect 7932 11101 7941 11135
rect 7941 11101 7975 11135
rect 7975 11101 7984 11135
rect 7932 11092 7984 11101
rect 10232 11135 10284 11144
rect 10232 11101 10266 11135
rect 10266 11101 10284 11135
rect 10232 11092 10284 11101
rect 14648 11339 14700 11348
rect 14648 11305 14657 11339
rect 14657 11305 14691 11339
rect 14691 11305 14700 11339
rect 14648 11296 14700 11305
rect 17132 11339 17184 11348
rect 17132 11305 17141 11339
rect 17141 11305 17175 11339
rect 17175 11305 17184 11339
rect 17132 11296 17184 11305
rect 17868 11296 17920 11348
rect 21456 11296 21508 11348
rect 21824 11296 21876 11348
rect 25504 11339 25556 11348
rect 25504 11305 25513 11339
rect 25513 11305 25547 11339
rect 25547 11305 25556 11339
rect 25504 11296 25556 11305
rect 26148 11339 26200 11348
rect 26148 11305 26157 11339
rect 26157 11305 26191 11339
rect 26191 11305 26200 11339
rect 26148 11296 26200 11305
rect 29644 11296 29696 11348
rect 14372 11135 14424 11144
rect 14372 11101 14381 11135
rect 14381 11101 14415 11135
rect 14415 11101 14424 11135
rect 14372 11092 14424 11101
rect 19708 11203 19760 11212
rect 19708 11169 19717 11203
rect 19717 11169 19751 11203
rect 19751 11169 19760 11203
rect 19708 11160 19760 11169
rect 8300 11024 8352 11076
rect 10876 11024 10928 11076
rect 12348 11024 12400 11076
rect 12900 11024 12952 11076
rect 16764 11092 16816 11144
rect 18512 11092 18564 11144
rect 20812 11092 20864 11144
rect 15844 11024 15896 11076
rect 22836 11228 22888 11280
rect 22652 11135 22704 11144
rect 22652 11101 22661 11135
rect 22661 11101 22695 11135
rect 22695 11101 22704 11135
rect 22652 11092 22704 11101
rect 28908 11228 28960 11280
rect 31852 11296 31904 11348
rect 33232 11296 33284 11348
rect 35256 11339 35308 11348
rect 35256 11305 35265 11339
rect 35265 11305 35299 11339
rect 35299 11305 35308 11339
rect 35256 11296 35308 11305
rect 36728 11296 36780 11348
rect 36452 11228 36504 11280
rect 24768 11203 24820 11212
rect 24768 11169 24777 11203
rect 24777 11169 24811 11203
rect 24811 11169 24820 11203
rect 24768 11160 24820 11169
rect 25044 11160 25096 11212
rect 33140 11160 33192 11212
rect 24676 11135 24728 11144
rect 24676 11101 24685 11135
rect 24685 11101 24719 11135
rect 24719 11101 24728 11135
rect 24676 11092 24728 11101
rect 25320 11092 25372 11144
rect 25412 11135 25464 11144
rect 25412 11101 25421 11135
rect 25421 11101 25455 11135
rect 25455 11101 25464 11135
rect 25412 11092 25464 11101
rect 25504 11092 25556 11144
rect 26056 11135 26108 11144
rect 26056 11101 26065 11135
rect 26065 11101 26099 11135
rect 26099 11101 26108 11135
rect 26056 11092 26108 11101
rect 29184 11092 29236 11144
rect 29736 11092 29788 11144
rect 30288 11135 30340 11144
rect 30288 11101 30297 11135
rect 30297 11101 30331 11135
rect 30331 11101 30340 11135
rect 30288 11092 30340 11101
rect 30656 11135 30708 11144
rect 30656 11101 30665 11135
rect 30665 11101 30699 11135
rect 30699 11101 30708 11135
rect 30656 11092 30708 11101
rect 32496 11092 32548 11144
rect 32588 11135 32640 11144
rect 32588 11101 32597 11135
rect 32597 11101 32631 11135
rect 32631 11101 32640 11135
rect 32588 11092 32640 11101
rect 32680 11092 32732 11144
rect 34980 11092 35032 11144
rect 35900 11160 35952 11212
rect 38384 11228 38436 11280
rect 38476 11228 38528 11280
rect 39120 11228 39172 11280
rect 35164 11092 35216 11144
rect 35992 11092 36044 11144
rect 36544 11135 36596 11144
rect 36544 11101 36553 11135
rect 36553 11101 36587 11135
rect 36587 11101 36596 11135
rect 36544 11092 36596 11101
rect 37648 11092 37700 11144
rect 38016 11135 38068 11144
rect 38016 11101 38025 11135
rect 38025 11101 38059 11135
rect 38059 11101 38068 11135
rect 38016 11092 38068 11101
rect 38752 11160 38804 11212
rect 38936 11160 38988 11212
rect 38292 11135 38344 11144
rect 38292 11101 38301 11135
rect 38301 11101 38335 11135
rect 38335 11101 38344 11135
rect 38292 11092 38344 11101
rect 38476 11092 38528 11144
rect 38660 11092 38712 11144
rect 38844 11092 38896 11144
rect 26240 11024 26292 11076
rect 32404 11024 32456 11076
rect 36452 11024 36504 11076
rect 36636 11024 36688 11076
rect 9588 10956 9640 11008
rect 11336 10999 11388 11008
rect 11336 10965 11345 10999
rect 11345 10965 11379 10999
rect 11379 10965 11388 10999
rect 11336 10956 11388 10965
rect 17224 10956 17276 11008
rect 21088 10956 21140 11008
rect 23204 10956 23256 11008
rect 24952 10956 25004 11008
rect 25228 10956 25280 11008
rect 26056 10956 26108 11008
rect 30932 10956 30984 11008
rect 32680 10956 32732 11008
rect 36360 10999 36412 11008
rect 36360 10965 36369 10999
rect 36369 10965 36403 10999
rect 36403 10965 36412 10999
rect 36360 10956 36412 10965
rect 37924 11024 37976 11076
rect 39764 11092 39816 11144
rect 40592 11160 40644 11212
rect 41696 11135 41748 11144
rect 41696 11101 41730 11135
rect 41730 11101 41748 11135
rect 41696 11092 41748 11101
rect 45008 11092 45060 11144
rect 42892 11024 42944 11076
rect 42800 10999 42852 11008
rect 42800 10965 42809 10999
rect 42809 10965 42843 10999
rect 42843 10965 42852 10999
rect 42800 10956 42852 10965
rect 11896 10854 11948 10906
rect 11960 10854 12012 10906
rect 12024 10854 12076 10906
rect 12088 10854 12140 10906
rect 12152 10854 12204 10906
rect 22843 10854 22895 10906
rect 22907 10854 22959 10906
rect 22971 10854 23023 10906
rect 23035 10854 23087 10906
rect 23099 10854 23151 10906
rect 33790 10854 33842 10906
rect 33854 10854 33906 10906
rect 33918 10854 33970 10906
rect 33982 10854 34034 10906
rect 34046 10854 34098 10906
rect 44737 10854 44789 10906
rect 44801 10854 44853 10906
rect 44865 10854 44917 10906
rect 44929 10854 44981 10906
rect 44993 10854 45045 10906
rect 4620 10752 4672 10804
rect 8300 10795 8352 10804
rect 8300 10761 8309 10795
rect 8309 10761 8343 10795
rect 8343 10761 8352 10795
rect 8300 10752 8352 10761
rect 10784 10795 10836 10804
rect 10784 10761 10793 10795
rect 10793 10761 10827 10795
rect 10827 10761 10836 10795
rect 10784 10752 10836 10761
rect 15844 10752 15896 10804
rect 16580 10752 16632 10804
rect 17040 10752 17092 10804
rect 17132 10752 17184 10804
rect 18696 10752 18748 10804
rect 3148 10684 3200 10736
rect 6092 10684 6144 10736
rect 1952 10616 2004 10668
rect 4068 10616 4120 10668
rect 4252 10659 4304 10668
rect 4252 10625 4286 10659
rect 4286 10625 4304 10659
rect 4252 10616 4304 10625
rect 9864 10684 9916 10736
rect 11336 10684 11388 10736
rect 8392 10616 8444 10668
rect 10968 10616 11020 10668
rect 11428 10616 11480 10668
rect 13912 10659 13964 10668
rect 13912 10625 13921 10659
rect 13921 10625 13955 10659
rect 13955 10625 13964 10659
rect 13912 10616 13964 10625
rect 14004 10616 14056 10668
rect 16856 10684 16908 10736
rect 20260 10727 20312 10736
rect 20260 10693 20269 10727
rect 20269 10693 20303 10727
rect 20303 10693 20312 10727
rect 20260 10684 20312 10693
rect 16304 10659 16356 10668
rect 16304 10625 16313 10659
rect 16313 10625 16347 10659
rect 16347 10625 16356 10659
rect 16304 10616 16356 10625
rect 17224 10616 17276 10668
rect 3148 10412 3200 10464
rect 10324 10480 10376 10532
rect 10876 10591 10928 10600
rect 10876 10557 10885 10591
rect 10885 10557 10919 10591
rect 10919 10557 10928 10591
rect 10876 10548 10928 10557
rect 14096 10591 14148 10600
rect 14096 10557 14105 10591
rect 14105 10557 14139 10591
rect 14139 10557 14148 10591
rect 14096 10548 14148 10557
rect 19432 10616 19484 10668
rect 20168 10616 20220 10668
rect 20812 10795 20864 10804
rect 20812 10761 20821 10795
rect 20821 10761 20855 10795
rect 20855 10761 20864 10795
rect 20812 10752 20864 10761
rect 21088 10752 21140 10804
rect 22652 10752 22704 10804
rect 25228 10752 25280 10804
rect 25320 10752 25372 10804
rect 26148 10795 26200 10804
rect 26148 10761 26157 10795
rect 26157 10761 26191 10795
rect 26191 10761 26200 10795
rect 26148 10752 26200 10761
rect 27436 10752 27488 10804
rect 30656 10752 30708 10804
rect 30932 10752 30984 10804
rect 32404 10795 32456 10804
rect 32404 10761 32413 10795
rect 32413 10761 32447 10795
rect 32447 10761 32456 10795
rect 32404 10752 32456 10761
rect 36452 10752 36504 10804
rect 38844 10795 38896 10804
rect 38844 10761 38853 10795
rect 38853 10761 38887 10795
rect 38887 10761 38896 10795
rect 38844 10752 38896 10761
rect 39028 10752 39080 10804
rect 43168 10795 43220 10804
rect 43168 10761 43177 10795
rect 43177 10761 43211 10795
rect 43211 10761 43220 10795
rect 43168 10752 43220 10761
rect 23204 10684 23256 10736
rect 24676 10684 24728 10736
rect 24768 10684 24820 10736
rect 25780 10684 25832 10736
rect 26056 10659 26108 10668
rect 26056 10625 26065 10659
rect 26065 10625 26099 10659
rect 26099 10625 26108 10659
rect 26056 10616 26108 10625
rect 38660 10684 38712 10736
rect 44456 10684 44508 10736
rect 27252 10659 27304 10668
rect 27252 10625 27261 10659
rect 27261 10625 27295 10659
rect 27295 10625 27304 10659
rect 27252 10616 27304 10625
rect 27620 10616 27672 10668
rect 28724 10616 28776 10668
rect 11060 10480 11112 10532
rect 14188 10480 14240 10532
rect 21180 10548 21232 10600
rect 22560 10548 22612 10600
rect 24584 10548 24636 10600
rect 31300 10659 31352 10668
rect 31300 10625 31309 10659
rect 31309 10625 31343 10659
rect 31343 10625 31352 10659
rect 31300 10616 31352 10625
rect 4620 10412 4672 10464
rect 15200 10412 15252 10464
rect 18696 10455 18748 10464
rect 18696 10421 18705 10455
rect 18705 10421 18739 10455
rect 18739 10421 18748 10455
rect 18696 10412 18748 10421
rect 22192 10455 22244 10464
rect 22192 10421 22201 10455
rect 22201 10421 22235 10455
rect 22235 10421 22244 10455
rect 22192 10412 22244 10421
rect 25412 10480 25464 10532
rect 35992 10659 36044 10668
rect 35992 10625 36001 10659
rect 36001 10625 36035 10659
rect 36035 10625 36044 10659
rect 35992 10616 36044 10625
rect 36820 10616 36872 10668
rect 37556 10616 37608 10668
rect 42800 10659 42852 10668
rect 42800 10625 42809 10659
rect 42809 10625 42843 10659
rect 42843 10625 42852 10659
rect 42800 10616 42852 10625
rect 44272 10548 44324 10600
rect 32864 10480 32916 10532
rect 38476 10480 38528 10532
rect 25320 10412 25372 10464
rect 29736 10412 29788 10464
rect 33508 10412 33560 10464
rect 36268 10412 36320 10464
rect 36360 10455 36412 10464
rect 36360 10421 36369 10455
rect 36369 10421 36403 10455
rect 36403 10421 36412 10455
rect 36360 10412 36412 10421
rect 36912 10412 36964 10464
rect 6423 10310 6475 10362
rect 6487 10310 6539 10362
rect 6551 10310 6603 10362
rect 6615 10310 6667 10362
rect 6679 10310 6731 10362
rect 17370 10310 17422 10362
rect 17434 10310 17486 10362
rect 17498 10310 17550 10362
rect 17562 10310 17614 10362
rect 17626 10310 17678 10362
rect 28317 10310 28369 10362
rect 28381 10310 28433 10362
rect 28445 10310 28497 10362
rect 28509 10310 28561 10362
rect 28573 10310 28625 10362
rect 39264 10310 39316 10362
rect 39328 10310 39380 10362
rect 39392 10310 39444 10362
rect 39456 10310 39508 10362
rect 39520 10310 39572 10362
rect 940 10208 992 10260
rect 7932 10251 7984 10260
rect 7932 10217 7941 10251
rect 7941 10217 7975 10251
rect 7975 10217 7984 10251
rect 7932 10208 7984 10217
rect 8392 10251 8444 10260
rect 8392 10217 8401 10251
rect 8401 10217 8435 10251
rect 8435 10217 8444 10251
rect 8392 10208 8444 10217
rect 11428 10208 11480 10260
rect 8484 10140 8536 10192
rect 3148 10115 3200 10124
rect 3148 10081 3157 10115
rect 3157 10081 3191 10115
rect 3191 10081 3200 10115
rect 3148 10072 3200 10081
rect 3424 10072 3476 10124
rect 9588 10115 9640 10124
rect 9588 10081 9597 10115
rect 9597 10081 9631 10115
rect 9631 10081 9640 10115
rect 9588 10072 9640 10081
rect 10600 10140 10652 10192
rect 24584 10208 24636 10260
rect 24676 10251 24728 10260
rect 24676 10217 24685 10251
rect 24685 10217 24719 10251
rect 24719 10217 24728 10251
rect 24676 10208 24728 10217
rect 38016 10208 38068 10260
rect 38292 10208 38344 10260
rect 38752 10251 38804 10260
rect 38752 10217 38761 10251
rect 38761 10217 38795 10251
rect 38795 10217 38804 10251
rect 38752 10208 38804 10217
rect 42892 10251 42944 10260
rect 42892 10217 42901 10251
rect 42901 10217 42935 10251
rect 42935 10217 42944 10251
rect 42892 10208 42944 10217
rect 14004 10140 14056 10192
rect 16304 10140 16356 10192
rect 16764 10140 16816 10192
rect 2780 10004 2832 10056
rect 3332 10004 3384 10056
rect 4620 10004 4672 10056
rect 7196 10004 7248 10056
rect 8576 10047 8628 10056
rect 8576 10013 8585 10047
rect 8585 10013 8619 10047
rect 8619 10013 8628 10047
rect 8576 10004 8628 10013
rect 10416 9979 10468 9988
rect 10416 9945 10425 9979
rect 10425 9945 10459 9979
rect 10459 9945 10468 9979
rect 10416 9936 10468 9945
rect 2228 9868 2280 9920
rect 4344 9868 4396 9920
rect 5908 9911 5960 9920
rect 5908 9877 5917 9911
rect 5917 9877 5951 9911
rect 5951 9877 5960 9911
rect 5908 9868 5960 9877
rect 9312 9868 9364 9920
rect 10048 9868 10100 9920
rect 13636 10072 13688 10124
rect 14280 10004 14332 10056
rect 14648 10047 14700 10056
rect 14648 10013 14657 10047
rect 14657 10013 14691 10047
rect 14691 10013 14700 10047
rect 14648 10004 14700 10013
rect 18420 10072 18472 10124
rect 19156 10072 19208 10124
rect 22744 10140 22796 10192
rect 17960 10004 18012 10056
rect 24952 10140 25004 10192
rect 24860 10072 24912 10124
rect 31852 10115 31904 10124
rect 31852 10081 31861 10115
rect 31861 10081 31895 10115
rect 31895 10081 31904 10115
rect 31852 10072 31904 10081
rect 36268 10072 36320 10124
rect 36820 10115 36872 10124
rect 36820 10081 36829 10115
rect 36829 10081 36863 10115
rect 36863 10081 36872 10115
rect 36820 10072 36872 10081
rect 21180 10047 21232 10056
rect 15660 9979 15712 9988
rect 15660 9945 15669 9979
rect 15669 9945 15703 9979
rect 15703 9945 15712 9979
rect 15660 9936 15712 9945
rect 13820 9868 13872 9920
rect 14372 9868 14424 9920
rect 14648 9868 14700 9920
rect 18052 9911 18104 9920
rect 18052 9877 18061 9911
rect 18061 9877 18095 9911
rect 18095 9877 18104 9911
rect 18052 9868 18104 9877
rect 18420 9911 18472 9920
rect 18420 9877 18429 9911
rect 18429 9877 18463 9911
rect 18463 9877 18472 9911
rect 18420 9868 18472 9877
rect 19524 9911 19576 9920
rect 19524 9877 19533 9911
rect 19533 9877 19567 9911
rect 19567 9877 19576 9911
rect 19524 9868 19576 9877
rect 21180 10013 21189 10047
rect 21189 10013 21223 10047
rect 21223 10013 21232 10047
rect 21180 10004 21232 10013
rect 22192 9936 22244 9988
rect 25504 10004 25556 10056
rect 29000 10004 29052 10056
rect 29736 10047 29788 10056
rect 29736 10013 29745 10047
rect 29745 10013 29779 10047
rect 29779 10013 29788 10047
rect 29736 10004 29788 10013
rect 29828 10004 29880 10056
rect 30932 10004 30984 10056
rect 31760 10047 31812 10056
rect 31760 10013 31769 10047
rect 31769 10013 31803 10047
rect 31803 10013 31812 10047
rect 31760 10004 31812 10013
rect 32680 10047 32732 10056
rect 32680 10013 32689 10047
rect 32689 10013 32723 10047
rect 32723 10013 32732 10047
rect 32680 10004 32732 10013
rect 32772 10047 32824 10056
rect 32772 10013 32781 10047
rect 32781 10013 32815 10047
rect 32815 10013 32824 10047
rect 32772 10004 32824 10013
rect 38660 10047 38712 10056
rect 38660 10013 38669 10047
rect 38669 10013 38703 10047
rect 38703 10013 38712 10047
rect 38660 10004 38712 10013
rect 43444 10004 43496 10056
rect 26424 9936 26476 9988
rect 36728 9936 36780 9988
rect 23572 9868 23624 9920
rect 25320 9868 25372 9920
rect 30656 9868 30708 9920
rect 32496 9868 32548 9920
rect 11896 9766 11948 9818
rect 11960 9766 12012 9818
rect 12024 9766 12076 9818
rect 12088 9766 12140 9818
rect 12152 9766 12204 9818
rect 22843 9766 22895 9818
rect 22907 9766 22959 9818
rect 22971 9766 23023 9818
rect 23035 9766 23087 9818
rect 23099 9766 23151 9818
rect 33790 9766 33842 9818
rect 33854 9766 33906 9818
rect 33918 9766 33970 9818
rect 33982 9766 34034 9818
rect 34046 9766 34098 9818
rect 44737 9766 44789 9818
rect 44801 9766 44853 9818
rect 44865 9766 44917 9818
rect 44929 9766 44981 9818
rect 44993 9766 45045 9818
rect 4620 9664 4672 9716
rect 6092 9664 6144 9716
rect 13820 9664 13872 9716
rect 14280 9707 14332 9716
rect 14280 9673 14289 9707
rect 14289 9673 14323 9707
rect 14323 9673 14332 9707
rect 14280 9664 14332 9673
rect 22652 9664 22704 9716
rect 2228 9571 2280 9580
rect 2228 9537 2237 9571
rect 2237 9537 2271 9571
rect 2271 9537 2280 9571
rect 2228 9528 2280 9537
rect 3332 9571 3384 9580
rect 3332 9537 3341 9571
rect 3341 9537 3375 9571
rect 3375 9537 3384 9571
rect 3332 9528 3384 9537
rect 4528 9392 4580 9444
rect 5540 9639 5592 9648
rect 5540 9605 5549 9639
rect 5549 9605 5583 9639
rect 5583 9605 5592 9639
rect 5540 9596 5592 9605
rect 9128 9596 9180 9648
rect 15200 9639 15252 9648
rect 6276 9528 6328 9580
rect 7196 9571 7248 9580
rect 7196 9537 7205 9571
rect 7205 9537 7239 9571
rect 7239 9537 7248 9571
rect 7196 9528 7248 9537
rect 7932 9528 7984 9580
rect 9772 9528 9824 9580
rect 11612 9528 11664 9580
rect 5540 9460 5592 9512
rect 5816 9503 5868 9512
rect 5816 9469 5825 9503
rect 5825 9469 5859 9503
rect 5859 9469 5868 9503
rect 5816 9460 5868 9469
rect 10692 9460 10744 9512
rect 12900 9571 12952 9580
rect 12900 9537 12909 9571
rect 12909 9537 12943 9571
rect 12943 9537 12952 9571
rect 12900 9528 12952 9537
rect 13176 9571 13228 9580
rect 13176 9537 13210 9571
rect 13210 9537 13228 9571
rect 13176 9528 13228 9537
rect 15200 9605 15234 9639
rect 15234 9605 15252 9639
rect 15200 9596 15252 9605
rect 18052 9596 18104 9648
rect 19524 9596 19576 9648
rect 22744 9596 22796 9648
rect 23572 9596 23624 9648
rect 25136 9664 25188 9716
rect 26424 9707 26476 9716
rect 26424 9673 26433 9707
rect 26433 9673 26467 9707
rect 26467 9673 26476 9707
rect 26424 9664 26476 9673
rect 31300 9664 31352 9716
rect 36728 9707 36780 9716
rect 36728 9673 36737 9707
rect 36737 9673 36771 9707
rect 36771 9673 36780 9707
rect 36728 9664 36780 9673
rect 25320 9596 25372 9648
rect 17960 9528 18012 9580
rect 18696 9528 18748 9580
rect 22560 9571 22612 9580
rect 22560 9537 22569 9571
rect 22569 9537 22603 9571
rect 22603 9537 22612 9571
rect 22560 9528 22612 9537
rect 25596 9528 25648 9580
rect 25780 9528 25832 9580
rect 16764 9460 16816 9512
rect 6920 9392 6972 9444
rect 10968 9392 11020 9444
rect 16396 9392 16448 9444
rect 2044 9367 2096 9376
rect 2044 9333 2053 9367
rect 2053 9333 2087 9367
rect 2087 9333 2096 9367
rect 2044 9324 2096 9333
rect 4252 9324 4304 9376
rect 8300 9324 8352 9376
rect 10324 9324 10376 9376
rect 16948 9367 17000 9376
rect 16948 9333 16957 9367
rect 16957 9333 16991 9367
rect 16991 9333 17000 9367
rect 16948 9324 17000 9333
rect 17776 9324 17828 9376
rect 20720 9324 20772 9376
rect 25044 9324 25096 9376
rect 26240 9571 26292 9580
rect 26240 9537 26249 9571
rect 26249 9537 26283 9571
rect 26283 9537 26292 9571
rect 26240 9528 26292 9537
rect 29000 9596 29052 9648
rect 29184 9596 29236 9648
rect 30656 9639 30708 9648
rect 30656 9605 30665 9639
rect 30665 9605 30699 9639
rect 30699 9605 30708 9639
rect 30656 9596 30708 9605
rect 27620 9460 27672 9512
rect 32772 9596 32824 9648
rect 32496 9571 32548 9580
rect 32496 9537 32505 9571
rect 32505 9537 32539 9571
rect 32539 9537 32548 9571
rect 32496 9528 32548 9537
rect 33508 9596 33560 9648
rect 33692 9596 33744 9648
rect 44088 9596 44140 9648
rect 30932 9435 30984 9444
rect 30932 9401 30941 9435
rect 30941 9401 30975 9435
rect 30975 9401 30984 9435
rect 30932 9392 30984 9401
rect 36360 9528 36412 9580
rect 36912 9571 36964 9580
rect 36912 9537 36921 9571
rect 36921 9537 36955 9571
rect 36955 9537 36964 9571
rect 36912 9528 36964 9537
rect 37740 9571 37792 9580
rect 37740 9537 37749 9571
rect 37749 9537 37783 9571
rect 37783 9537 37792 9571
rect 37740 9528 37792 9537
rect 34980 9503 35032 9512
rect 34980 9469 34989 9503
rect 34989 9469 35023 9503
rect 35023 9469 35032 9503
rect 34980 9460 35032 9469
rect 29828 9324 29880 9376
rect 31668 9324 31720 9376
rect 32956 9324 33008 9376
rect 35716 9392 35768 9444
rect 34336 9324 34388 9376
rect 37556 9367 37608 9376
rect 37556 9333 37565 9367
rect 37565 9333 37599 9367
rect 37599 9333 37608 9367
rect 37556 9324 37608 9333
rect 6423 9222 6475 9274
rect 6487 9222 6539 9274
rect 6551 9222 6603 9274
rect 6615 9222 6667 9274
rect 6679 9222 6731 9274
rect 17370 9222 17422 9274
rect 17434 9222 17486 9274
rect 17498 9222 17550 9274
rect 17562 9222 17614 9274
rect 17626 9222 17678 9274
rect 28317 9222 28369 9274
rect 28381 9222 28433 9274
rect 28445 9222 28497 9274
rect 28509 9222 28561 9274
rect 28573 9222 28625 9274
rect 39264 9222 39316 9274
rect 39328 9222 39380 9274
rect 39392 9222 39444 9274
rect 39456 9222 39508 9274
rect 39520 9222 39572 9274
rect 10692 9120 10744 9172
rect 11612 9163 11664 9172
rect 11612 9129 11621 9163
rect 11621 9129 11655 9163
rect 11655 9129 11664 9163
rect 11612 9120 11664 9129
rect 13912 9120 13964 9172
rect 16120 9120 16172 9172
rect 17960 9120 18012 9172
rect 18420 9120 18472 9172
rect 19064 9120 19116 9172
rect 19432 9163 19484 9172
rect 19432 9129 19441 9163
rect 19441 9129 19475 9163
rect 19475 9129 19484 9163
rect 19432 9120 19484 9129
rect 3424 8984 3476 9036
rect 5816 8984 5868 9036
rect 8484 9027 8536 9036
rect 8484 8993 8493 9027
rect 8493 8993 8527 9027
rect 8527 8993 8536 9027
rect 8484 8984 8536 8993
rect 9772 9027 9824 9036
rect 9772 8993 9781 9027
rect 9781 8993 9815 9027
rect 9815 8993 9824 9027
rect 9772 8984 9824 8993
rect 5356 8916 5408 8968
rect 5632 8959 5684 8968
rect 5632 8925 5641 8959
rect 5641 8925 5675 8959
rect 5675 8925 5684 8959
rect 5632 8916 5684 8925
rect 8208 8916 8260 8968
rect 9312 8959 9364 8968
rect 9312 8925 9321 8959
rect 9321 8925 9355 8959
rect 9355 8925 9364 8959
rect 9312 8916 9364 8925
rect 10324 8916 10376 8968
rect 3240 8848 3292 8900
rect 13636 9052 13688 9104
rect 15476 8984 15528 9036
rect 16948 8984 17000 9036
rect 19156 8984 19208 9036
rect 11796 8959 11848 8968
rect 11796 8925 11805 8959
rect 11805 8925 11839 8959
rect 11839 8925 11848 8959
rect 11796 8916 11848 8925
rect 13176 8916 13228 8968
rect 16856 8916 16908 8968
rect 17132 8916 17184 8968
rect 2228 8780 2280 8832
rect 6828 8780 6880 8832
rect 8944 8780 8996 8832
rect 14740 8823 14792 8832
rect 14740 8789 14749 8823
rect 14749 8789 14783 8823
rect 14783 8789 14792 8823
rect 14740 8780 14792 8789
rect 16212 8823 16264 8832
rect 16212 8789 16221 8823
rect 16221 8789 16255 8823
rect 16255 8789 16264 8823
rect 16212 8780 16264 8789
rect 17776 8848 17828 8900
rect 20720 8848 20772 8900
rect 32956 9120 33008 9172
rect 33692 9120 33744 9172
rect 34152 9163 34204 9172
rect 34152 9129 34161 9163
rect 34161 9129 34195 9163
rect 34195 9129 34204 9163
rect 34152 9120 34204 9129
rect 20996 9052 21048 9104
rect 21916 9052 21968 9104
rect 27528 9052 27580 9104
rect 29184 9052 29236 9104
rect 29828 9095 29880 9104
rect 29828 9061 29837 9095
rect 29837 9061 29871 9095
rect 29871 9061 29880 9095
rect 29828 9052 29880 9061
rect 32680 9052 32732 9104
rect 35716 9120 35768 9172
rect 36360 9163 36412 9172
rect 36360 9129 36369 9163
rect 36369 9129 36403 9163
rect 36403 9129 36412 9163
rect 36360 9120 36412 9129
rect 25044 9027 25096 9036
rect 25044 8993 25053 9027
rect 25053 8993 25087 9027
rect 25087 8993 25096 9027
rect 25044 8984 25096 8993
rect 25780 8984 25832 9036
rect 21548 8916 21600 8968
rect 24584 8916 24636 8968
rect 26608 8984 26660 9036
rect 27344 8984 27396 9036
rect 29000 8959 29052 8968
rect 29000 8925 29009 8959
rect 29009 8925 29043 8959
rect 29043 8925 29052 8959
rect 29000 8916 29052 8925
rect 30656 8984 30708 9036
rect 21088 8848 21140 8900
rect 22744 8848 22796 8900
rect 25688 8848 25740 8900
rect 27712 8891 27764 8900
rect 27712 8857 27721 8891
rect 27721 8857 27755 8891
rect 27755 8857 27764 8891
rect 27712 8848 27764 8857
rect 28908 8848 28960 8900
rect 22652 8780 22704 8832
rect 24032 8823 24084 8832
rect 24032 8789 24041 8823
rect 24041 8789 24075 8823
rect 24075 8789 24084 8823
rect 24032 8780 24084 8789
rect 25964 8780 26016 8832
rect 27620 8823 27672 8832
rect 27620 8789 27629 8823
rect 27629 8789 27663 8823
rect 27663 8789 27672 8823
rect 27620 8780 27672 8789
rect 30196 8823 30248 8832
rect 30196 8789 30205 8823
rect 30205 8789 30239 8823
rect 30239 8789 30248 8823
rect 30196 8780 30248 8789
rect 30288 8823 30340 8832
rect 30288 8789 30297 8823
rect 30297 8789 30331 8823
rect 30331 8789 30340 8823
rect 30288 8780 30340 8789
rect 31576 8916 31628 8968
rect 34520 8984 34572 9036
rect 32956 8959 33008 8968
rect 32956 8925 32965 8959
rect 32965 8925 32999 8959
rect 32999 8925 33008 8959
rect 32956 8916 33008 8925
rect 34336 8959 34388 8968
rect 34336 8925 34345 8959
rect 34345 8925 34379 8959
rect 34379 8925 34388 8959
rect 34336 8916 34388 8925
rect 34612 8916 34664 8968
rect 37464 8959 37516 8968
rect 37464 8925 37473 8959
rect 37473 8925 37507 8959
rect 37507 8925 37516 8959
rect 37464 8916 37516 8925
rect 37556 8916 37608 8968
rect 44364 8959 44416 8968
rect 44364 8925 44373 8959
rect 44373 8925 44407 8959
rect 44407 8925 44416 8959
rect 44364 8916 44416 8925
rect 31484 8848 31536 8900
rect 34152 8848 34204 8900
rect 31944 8780 31996 8832
rect 34980 8780 35032 8832
rect 38936 8848 38988 8900
rect 37924 8780 37976 8832
rect 44180 8823 44232 8832
rect 44180 8789 44189 8823
rect 44189 8789 44223 8823
rect 44223 8789 44232 8823
rect 44180 8780 44232 8789
rect 11896 8678 11948 8730
rect 11960 8678 12012 8730
rect 12024 8678 12076 8730
rect 12088 8678 12140 8730
rect 12152 8678 12204 8730
rect 22843 8678 22895 8730
rect 22907 8678 22959 8730
rect 22971 8678 23023 8730
rect 23035 8678 23087 8730
rect 23099 8678 23151 8730
rect 33790 8678 33842 8730
rect 33854 8678 33906 8730
rect 33918 8678 33970 8730
rect 33982 8678 34034 8730
rect 34046 8678 34098 8730
rect 44737 8678 44789 8730
rect 44801 8678 44853 8730
rect 44865 8678 44917 8730
rect 44929 8678 44981 8730
rect 44993 8678 45045 8730
rect 2044 8576 2096 8628
rect 4344 8576 4396 8628
rect 2228 8440 2280 8492
rect 8208 8619 8260 8628
rect 8208 8585 8217 8619
rect 8217 8585 8251 8619
rect 8251 8585 8260 8619
rect 8208 8576 8260 8585
rect 9680 8576 9732 8628
rect 10048 8619 10100 8628
rect 10048 8585 10057 8619
rect 10057 8585 10091 8619
rect 10091 8585 10100 8619
rect 10048 8576 10100 8585
rect 15660 8576 15712 8628
rect 8944 8551 8996 8560
rect 8944 8517 8978 8551
rect 8978 8517 8996 8551
rect 8944 8508 8996 8517
rect 3976 8483 4028 8492
rect 3976 8449 3985 8483
rect 3985 8449 4019 8483
rect 4019 8449 4028 8483
rect 3976 8440 4028 8449
rect 9496 8440 9548 8492
rect 8300 8372 8352 8424
rect 8668 8415 8720 8424
rect 8668 8381 8677 8415
rect 8677 8381 8711 8415
rect 8711 8381 8720 8415
rect 8668 8372 8720 8381
rect 14372 8483 14424 8492
rect 14372 8449 14381 8483
rect 14381 8449 14415 8483
rect 14415 8449 14424 8483
rect 14372 8440 14424 8449
rect 16120 8483 16172 8492
rect 16120 8449 16129 8483
rect 16129 8449 16163 8483
rect 16163 8449 16172 8483
rect 16120 8440 16172 8449
rect 17132 8508 17184 8560
rect 17224 8508 17276 8560
rect 20260 8508 20312 8560
rect 21088 8508 21140 8560
rect 24032 8508 24084 8560
rect 25596 8619 25648 8628
rect 25596 8585 25605 8619
rect 25605 8585 25639 8619
rect 25639 8585 25648 8619
rect 25596 8576 25648 8585
rect 25964 8619 26016 8628
rect 25964 8585 25973 8619
rect 25973 8585 26007 8619
rect 26007 8585 26016 8619
rect 25964 8576 26016 8585
rect 30196 8576 30248 8628
rect 31484 8619 31536 8628
rect 31484 8585 31493 8619
rect 31493 8585 31527 8619
rect 31527 8585 31536 8619
rect 31484 8576 31536 8585
rect 28724 8508 28776 8560
rect 19064 8483 19116 8492
rect 19064 8449 19073 8483
rect 19073 8449 19107 8483
rect 19107 8449 19116 8483
rect 19064 8440 19116 8449
rect 19800 8440 19852 8492
rect 19892 8483 19944 8492
rect 19892 8449 19901 8483
rect 19901 8449 19935 8483
rect 19935 8449 19944 8483
rect 19892 8440 19944 8449
rect 20352 8440 20404 8492
rect 20720 8483 20772 8492
rect 20720 8449 20729 8483
rect 20729 8449 20763 8483
rect 20763 8449 20772 8483
rect 20720 8440 20772 8449
rect 22008 8483 22060 8492
rect 22008 8449 22017 8483
rect 22017 8449 22051 8483
rect 22051 8449 22060 8483
rect 22008 8440 22060 8449
rect 23388 8440 23440 8492
rect 27620 8440 27672 8492
rect 32496 8508 32548 8560
rect 34520 8576 34572 8628
rect 37740 8576 37792 8628
rect 37832 8576 37884 8628
rect 29736 8440 29788 8492
rect 30196 8440 30248 8492
rect 31576 8440 31628 8492
rect 31668 8483 31720 8492
rect 31668 8449 31677 8483
rect 31677 8449 31711 8483
rect 31711 8449 31720 8483
rect 31668 8440 31720 8449
rect 34520 8440 34572 8492
rect 34612 8483 34664 8492
rect 34612 8449 34621 8483
rect 34621 8449 34655 8483
rect 34655 8449 34664 8483
rect 34612 8440 34664 8449
rect 37924 8440 37976 8492
rect 42616 8440 42668 8492
rect 14924 8372 14976 8424
rect 16212 8372 16264 8424
rect 26148 8415 26200 8424
rect 26148 8381 26157 8415
rect 26157 8381 26191 8415
rect 26191 8381 26200 8415
rect 26148 8372 26200 8381
rect 3240 8304 3292 8356
rect 6920 8347 6972 8356
rect 6920 8313 6929 8347
rect 6929 8313 6963 8347
rect 6963 8313 6972 8347
rect 6920 8304 6972 8313
rect 14648 8236 14700 8288
rect 18604 8347 18656 8356
rect 18604 8313 18613 8347
rect 18613 8313 18647 8347
rect 18647 8313 18656 8347
rect 18604 8304 18656 8313
rect 17224 8236 17276 8288
rect 20076 8236 20128 8288
rect 22192 8236 22244 8288
rect 28172 8236 28224 8288
rect 28908 8372 28960 8424
rect 35716 8372 35768 8424
rect 35624 8304 35676 8356
rect 41420 8304 41472 8356
rect 29184 8279 29236 8288
rect 29184 8245 29193 8279
rect 29193 8245 29227 8279
rect 29227 8245 29236 8279
rect 29184 8236 29236 8245
rect 6423 8134 6475 8186
rect 6487 8134 6539 8186
rect 6551 8134 6603 8186
rect 6615 8134 6667 8186
rect 6679 8134 6731 8186
rect 17370 8134 17422 8186
rect 17434 8134 17486 8186
rect 17498 8134 17550 8186
rect 17562 8134 17614 8186
rect 17626 8134 17678 8186
rect 28317 8134 28369 8186
rect 28381 8134 28433 8186
rect 28445 8134 28497 8186
rect 28509 8134 28561 8186
rect 28573 8134 28625 8186
rect 39264 8134 39316 8186
rect 39328 8134 39380 8186
rect 39392 8134 39444 8186
rect 39456 8134 39508 8186
rect 39520 8134 39572 8186
rect 5356 8075 5408 8084
rect 5356 8041 5365 8075
rect 5365 8041 5399 8075
rect 5399 8041 5408 8075
rect 5356 8032 5408 8041
rect 6276 8032 6328 8084
rect 8576 8032 8628 8084
rect 11796 8032 11848 8084
rect 14924 8032 14976 8084
rect 3332 7896 3384 7948
rect 3884 7896 3936 7948
rect 5908 7939 5960 7948
rect 5908 7905 5917 7939
rect 5917 7905 5951 7939
rect 5951 7905 5960 7939
rect 5908 7896 5960 7905
rect 9128 7939 9180 7948
rect 9128 7905 9137 7939
rect 9137 7905 9171 7939
rect 9171 7905 9180 7939
rect 9128 7896 9180 7905
rect 2320 7803 2372 7812
rect 2320 7769 2354 7803
rect 2354 7769 2372 7803
rect 2320 7760 2372 7769
rect 8024 7871 8076 7880
rect 8024 7837 8033 7871
rect 8033 7837 8067 7871
rect 8067 7837 8076 7871
rect 8024 7828 8076 7837
rect 8576 7828 8628 7880
rect 10508 7828 10560 7880
rect 14096 7896 14148 7948
rect 4436 7760 4488 7812
rect 7932 7760 7984 7812
rect 8300 7760 8352 7812
rect 9772 7760 9824 7812
rect 11152 7760 11204 7812
rect 13360 7871 13412 7880
rect 13360 7837 13369 7871
rect 13369 7837 13403 7871
rect 13403 7837 13412 7871
rect 13360 7828 13412 7837
rect 14464 7828 14516 7880
rect 15292 7828 15344 7880
rect 18144 7896 18196 7948
rect 16120 7828 16172 7880
rect 17132 7871 17184 7880
rect 17132 7837 17141 7871
rect 17141 7837 17175 7871
rect 17175 7837 17184 7871
rect 17132 7828 17184 7837
rect 25688 8075 25740 8084
rect 25688 8041 25697 8075
rect 25697 8041 25731 8075
rect 25731 8041 25740 8075
rect 25688 8032 25740 8041
rect 29736 8075 29788 8084
rect 29736 8041 29745 8075
rect 29745 8041 29779 8075
rect 29779 8041 29788 8075
rect 29736 8032 29788 8041
rect 34520 8032 34572 8084
rect 23940 7964 23992 8016
rect 29000 7964 29052 8016
rect 30196 7964 30248 8016
rect 19800 7896 19852 7948
rect 20352 7896 20404 7948
rect 13728 7760 13780 7812
rect 15016 7760 15068 7812
rect 5632 7692 5684 7744
rect 10508 7735 10560 7744
rect 10508 7701 10517 7735
rect 10517 7701 10551 7735
rect 10551 7701 10560 7735
rect 10508 7692 10560 7701
rect 11612 7735 11664 7744
rect 11612 7701 11621 7735
rect 11621 7701 11655 7735
rect 11655 7701 11664 7735
rect 11612 7692 11664 7701
rect 12992 7692 13044 7744
rect 14372 7692 14424 7744
rect 15108 7692 15160 7744
rect 15200 7735 15252 7744
rect 15200 7701 15209 7735
rect 15209 7701 15243 7735
rect 15243 7701 15252 7735
rect 15200 7692 15252 7701
rect 19892 7871 19944 7880
rect 19892 7837 19901 7871
rect 19901 7837 19935 7871
rect 19935 7837 19944 7871
rect 19892 7828 19944 7837
rect 20260 7871 20312 7880
rect 20260 7837 20269 7871
rect 20269 7837 20303 7871
rect 20303 7837 20312 7871
rect 20260 7828 20312 7837
rect 21548 7939 21600 7948
rect 21548 7905 21557 7939
rect 21557 7905 21591 7939
rect 21591 7905 21600 7939
rect 21548 7896 21600 7905
rect 24032 7896 24084 7948
rect 21088 7871 21140 7880
rect 21088 7837 21097 7871
rect 21097 7837 21131 7871
rect 21131 7837 21140 7871
rect 21088 7828 21140 7837
rect 22376 7828 22428 7880
rect 25964 7896 26016 7948
rect 27620 7896 27672 7948
rect 32956 7896 33008 7948
rect 34704 7896 34756 7948
rect 35716 7896 35768 7948
rect 37924 7896 37976 7948
rect 40500 8032 40552 8084
rect 25504 7828 25556 7880
rect 29184 7828 29236 7880
rect 19340 7692 19392 7744
rect 19984 7692 20036 7744
rect 20720 7692 20772 7744
rect 20996 7735 21048 7744
rect 20996 7701 21005 7735
rect 21005 7701 21039 7735
rect 21039 7701 21048 7735
rect 20996 7692 21048 7701
rect 22008 7692 22060 7744
rect 31024 7828 31076 7880
rect 32588 7871 32640 7880
rect 32588 7837 32597 7871
rect 32597 7837 32631 7871
rect 32631 7837 32640 7871
rect 32588 7828 32640 7837
rect 35624 7828 35676 7880
rect 39120 7828 39172 7880
rect 38936 7760 38988 7812
rect 39304 7871 39356 7880
rect 39304 7837 39313 7871
rect 39313 7837 39347 7871
rect 39347 7837 39356 7871
rect 39304 7828 39356 7837
rect 40040 7871 40092 7880
rect 40040 7837 40049 7871
rect 40049 7837 40083 7871
rect 40083 7837 40092 7871
rect 40040 7828 40092 7837
rect 41420 7828 41472 7880
rect 39856 7760 39908 7812
rect 40316 7803 40368 7812
rect 40316 7769 40325 7803
rect 40325 7769 40359 7803
rect 40359 7769 40368 7803
rect 40316 7760 40368 7769
rect 42524 7803 42576 7812
rect 42524 7769 42533 7803
rect 42533 7769 42567 7803
rect 42567 7769 42576 7803
rect 42524 7760 42576 7769
rect 42984 7760 43036 7812
rect 32404 7735 32456 7744
rect 32404 7701 32413 7735
rect 32413 7701 32447 7735
rect 32447 7701 32456 7735
rect 32404 7692 32456 7701
rect 35532 7692 35584 7744
rect 38752 7692 38804 7744
rect 40224 7692 40276 7744
rect 40408 7692 40460 7744
rect 43996 7735 44048 7744
rect 43996 7701 44005 7735
rect 44005 7701 44039 7735
rect 44039 7701 44048 7735
rect 43996 7692 44048 7701
rect 11896 7590 11948 7642
rect 11960 7590 12012 7642
rect 12024 7590 12076 7642
rect 12088 7590 12140 7642
rect 12152 7590 12204 7642
rect 22843 7590 22895 7642
rect 22907 7590 22959 7642
rect 22971 7590 23023 7642
rect 23035 7590 23087 7642
rect 23099 7590 23151 7642
rect 33790 7590 33842 7642
rect 33854 7590 33906 7642
rect 33918 7590 33970 7642
rect 33982 7590 34034 7642
rect 34046 7590 34098 7642
rect 44737 7590 44789 7642
rect 44801 7590 44853 7642
rect 44865 7590 44917 7642
rect 44929 7590 44981 7642
rect 44993 7590 45045 7642
rect 3884 7531 3936 7540
rect 3884 7497 3893 7531
rect 3893 7497 3927 7531
rect 3927 7497 3936 7531
rect 3884 7488 3936 7497
rect 5632 7531 5684 7540
rect 5632 7497 5641 7531
rect 5641 7497 5675 7531
rect 5675 7497 5684 7531
rect 5632 7488 5684 7497
rect 5724 7488 5776 7540
rect 9128 7531 9180 7540
rect 9128 7497 9137 7531
rect 9137 7497 9171 7531
rect 9171 7497 9180 7531
rect 9128 7488 9180 7497
rect 9496 7488 9548 7540
rect 11612 7488 11664 7540
rect 14464 7531 14516 7540
rect 14464 7497 14473 7531
rect 14473 7497 14507 7531
rect 14507 7497 14516 7531
rect 14464 7488 14516 7497
rect 16856 7531 16908 7540
rect 16856 7497 16865 7531
rect 16865 7497 16899 7531
rect 16899 7497 16908 7531
rect 16856 7488 16908 7497
rect 17868 7488 17920 7540
rect 18144 7531 18196 7540
rect 18144 7497 18153 7531
rect 18153 7497 18187 7531
rect 18187 7497 18196 7531
rect 18144 7488 18196 7497
rect 19340 7488 19392 7540
rect 20168 7488 20220 7540
rect 20996 7488 21048 7540
rect 22376 7531 22428 7540
rect 22376 7497 22385 7531
rect 22385 7497 22419 7531
rect 22419 7497 22428 7531
rect 22376 7488 22428 7497
rect 22744 7488 22796 7540
rect 30748 7531 30800 7540
rect 30748 7497 30757 7531
rect 30757 7497 30791 7531
rect 30791 7497 30800 7531
rect 30748 7488 30800 7497
rect 6828 7420 6880 7472
rect 7932 7420 7984 7472
rect 940 7352 992 7404
rect 5540 7395 5592 7404
rect 5540 7361 5549 7395
rect 5549 7361 5583 7395
rect 5583 7361 5592 7395
rect 5540 7352 5592 7361
rect 5356 7284 5408 7336
rect 9312 7352 9364 7404
rect 12624 7395 12676 7404
rect 12624 7361 12633 7395
rect 12633 7361 12667 7395
rect 12667 7361 12676 7395
rect 12624 7352 12676 7361
rect 15200 7420 15252 7472
rect 17224 7463 17276 7472
rect 17224 7429 17233 7463
rect 17233 7429 17267 7463
rect 17267 7429 17276 7463
rect 17224 7420 17276 7429
rect 18604 7420 18656 7472
rect 5816 7327 5868 7336
rect 5816 7293 5825 7327
rect 5825 7293 5859 7327
rect 5859 7293 5868 7327
rect 5816 7284 5868 7293
rect 8024 7284 8076 7336
rect 9772 7284 9824 7336
rect 10600 7327 10652 7336
rect 10600 7293 10609 7327
rect 10609 7293 10643 7327
rect 10643 7293 10652 7327
rect 10600 7284 10652 7293
rect 12256 7284 12308 7336
rect 14924 7395 14976 7404
rect 14924 7361 14933 7395
rect 14933 7361 14967 7395
rect 14967 7361 14976 7395
rect 14924 7352 14976 7361
rect 15108 7395 15160 7404
rect 15108 7361 15117 7395
rect 15117 7361 15151 7395
rect 15151 7361 15160 7395
rect 15108 7352 15160 7361
rect 18328 7284 18380 7336
rect 18880 7352 18932 7404
rect 20076 7395 20128 7404
rect 20076 7361 20085 7395
rect 20085 7361 20119 7395
rect 20119 7361 20128 7395
rect 20076 7352 20128 7361
rect 20720 7395 20772 7404
rect 20720 7361 20729 7395
rect 20729 7361 20763 7395
rect 20763 7361 20772 7395
rect 20720 7352 20772 7361
rect 21916 7420 21968 7472
rect 32404 7420 32456 7472
rect 32680 7420 32732 7472
rect 22652 7352 22704 7404
rect 23756 7395 23808 7404
rect 23756 7361 23765 7395
rect 23765 7361 23799 7395
rect 23799 7361 23808 7395
rect 23756 7352 23808 7361
rect 25504 7352 25556 7404
rect 28816 7395 28868 7404
rect 28816 7361 28850 7395
rect 28850 7361 28868 7395
rect 28816 7352 28868 7361
rect 38752 7463 38804 7472
rect 38752 7429 38761 7463
rect 38761 7429 38795 7463
rect 38795 7429 38804 7463
rect 38752 7420 38804 7429
rect 38936 7463 38988 7472
rect 38936 7429 38945 7463
rect 38945 7429 38979 7463
rect 38979 7429 38988 7463
rect 38936 7420 38988 7429
rect 19156 7284 19208 7336
rect 20996 7327 21048 7336
rect 20996 7293 21005 7327
rect 21005 7293 21039 7327
rect 21039 7293 21048 7327
rect 20996 7284 21048 7293
rect 23940 7327 23992 7336
rect 23940 7293 23949 7327
rect 23949 7293 23983 7327
rect 23983 7293 23992 7327
rect 23940 7284 23992 7293
rect 28172 7284 28224 7336
rect 30472 7284 30524 7336
rect 35532 7395 35584 7404
rect 35532 7361 35541 7395
rect 35541 7361 35575 7395
rect 35575 7361 35584 7395
rect 35532 7352 35584 7361
rect 35624 7352 35676 7404
rect 36084 7395 36136 7404
rect 36084 7361 36093 7395
rect 36093 7361 36127 7395
rect 36127 7361 36136 7395
rect 36084 7352 36136 7361
rect 39304 7488 39356 7540
rect 42524 7488 42576 7540
rect 42984 7488 43036 7540
rect 44272 7488 44324 7540
rect 31208 7284 31260 7336
rect 5172 7191 5224 7200
rect 5172 7157 5181 7191
rect 5181 7157 5215 7191
rect 5215 7157 5224 7191
rect 5172 7148 5224 7157
rect 12440 7191 12492 7200
rect 12440 7157 12449 7191
rect 12449 7157 12483 7191
rect 12483 7157 12492 7191
rect 12440 7148 12492 7157
rect 14740 7148 14792 7200
rect 14924 7191 14976 7200
rect 14924 7157 14933 7191
rect 14933 7157 14967 7191
rect 14967 7157 14976 7191
rect 14924 7148 14976 7157
rect 15016 7148 15068 7200
rect 19892 7148 19944 7200
rect 20720 7148 20772 7200
rect 20812 7191 20864 7200
rect 20812 7157 20821 7191
rect 20821 7157 20855 7191
rect 20855 7157 20864 7191
rect 20812 7148 20864 7157
rect 22192 7191 22244 7200
rect 22192 7157 22201 7191
rect 22201 7157 22235 7191
rect 22235 7157 22244 7191
rect 22192 7148 22244 7157
rect 25596 7148 25648 7200
rect 30012 7148 30064 7200
rect 33508 7148 33560 7200
rect 35440 7284 35492 7336
rect 35900 7327 35952 7336
rect 35900 7293 35909 7327
rect 35909 7293 35943 7327
rect 35943 7293 35952 7327
rect 35900 7284 35952 7293
rect 36360 7284 36412 7336
rect 39856 7395 39908 7404
rect 39856 7361 39865 7395
rect 39865 7361 39899 7395
rect 39899 7361 39908 7395
rect 39856 7352 39908 7361
rect 40224 7420 40276 7472
rect 40500 7420 40552 7472
rect 40224 7284 40276 7336
rect 40316 7216 40368 7268
rect 42616 7395 42668 7404
rect 42616 7361 42625 7395
rect 42625 7361 42659 7395
rect 42659 7361 42668 7395
rect 42616 7352 42668 7361
rect 44364 7395 44416 7404
rect 44364 7361 44373 7395
rect 44373 7361 44407 7395
rect 44407 7361 44416 7395
rect 44364 7352 44416 7361
rect 35256 7148 35308 7200
rect 36268 7191 36320 7200
rect 36268 7157 36277 7191
rect 36277 7157 36311 7191
rect 36311 7157 36320 7191
rect 36268 7148 36320 7157
rect 39948 7148 40000 7200
rect 41236 7148 41288 7200
rect 6423 7046 6475 7098
rect 6487 7046 6539 7098
rect 6551 7046 6603 7098
rect 6615 7046 6667 7098
rect 6679 7046 6731 7098
rect 17370 7046 17422 7098
rect 17434 7046 17486 7098
rect 17498 7046 17550 7098
rect 17562 7046 17614 7098
rect 17626 7046 17678 7098
rect 28317 7046 28369 7098
rect 28381 7046 28433 7098
rect 28445 7046 28497 7098
rect 28509 7046 28561 7098
rect 28573 7046 28625 7098
rect 39264 7046 39316 7098
rect 39328 7046 39380 7098
rect 39392 7046 39444 7098
rect 39456 7046 39508 7098
rect 39520 7046 39572 7098
rect 8576 6987 8628 6996
rect 8576 6953 8585 6987
rect 8585 6953 8619 6987
rect 8619 6953 8628 6987
rect 8576 6944 8628 6953
rect 12532 6944 12584 6996
rect 13728 6987 13780 6996
rect 13728 6953 13737 6987
rect 13737 6953 13771 6987
rect 13771 6953 13780 6987
rect 13728 6944 13780 6953
rect 14648 6987 14700 6996
rect 14648 6953 14657 6987
rect 14657 6953 14691 6987
rect 14691 6953 14700 6987
rect 14648 6944 14700 6953
rect 3424 6808 3476 6860
rect 3976 6851 4028 6860
rect 3976 6817 3985 6851
rect 3985 6817 4019 6851
rect 4019 6817 4028 6851
rect 3976 6808 4028 6817
rect 11612 6808 11664 6860
rect 7932 6740 7984 6792
rect 8668 6740 8720 6792
rect 9128 6740 9180 6792
rect 9772 6783 9824 6792
rect 9772 6749 9781 6783
rect 9781 6749 9815 6783
rect 9815 6749 9824 6783
rect 9772 6740 9824 6749
rect 11796 6740 11848 6792
rect 2136 6647 2188 6656
rect 2136 6613 2145 6647
rect 2145 6613 2179 6647
rect 2179 6613 2188 6647
rect 2136 6604 2188 6613
rect 2872 6604 2924 6656
rect 3240 6672 3292 6724
rect 14832 6808 14884 6860
rect 12256 6740 12308 6792
rect 12440 6740 12492 6792
rect 14280 6783 14332 6792
rect 14280 6749 14289 6783
rect 14289 6749 14323 6783
rect 14323 6749 14332 6783
rect 14280 6740 14332 6749
rect 14924 6740 14976 6792
rect 19340 6944 19392 6996
rect 18420 6876 18472 6928
rect 28816 6944 28868 6996
rect 32588 6944 32640 6996
rect 39120 6987 39172 6996
rect 39120 6953 39129 6987
rect 39129 6953 39163 6987
rect 39163 6953 39172 6987
rect 39120 6944 39172 6953
rect 39488 6944 39540 6996
rect 17224 6783 17276 6792
rect 17224 6749 17230 6783
rect 17230 6749 17264 6783
rect 17264 6749 17276 6783
rect 17224 6740 17276 6749
rect 18788 6808 18840 6860
rect 18880 6851 18932 6860
rect 18880 6817 18889 6851
rect 18889 6817 18923 6851
rect 18923 6817 18932 6851
rect 18880 6808 18932 6817
rect 5264 6604 5316 6656
rect 5540 6604 5592 6656
rect 6000 6604 6052 6656
rect 9404 6604 9456 6656
rect 9680 6647 9732 6656
rect 9680 6613 9689 6647
rect 9689 6613 9723 6647
rect 9723 6613 9732 6647
rect 9680 6604 9732 6613
rect 14464 6672 14516 6724
rect 15108 6672 15160 6724
rect 18420 6783 18472 6792
rect 18420 6749 18429 6783
rect 18429 6749 18463 6783
rect 18463 6749 18472 6783
rect 18420 6740 18472 6749
rect 18512 6783 18564 6792
rect 18512 6749 18521 6783
rect 18521 6749 18555 6783
rect 18555 6749 18564 6783
rect 18512 6740 18564 6749
rect 18604 6740 18656 6792
rect 19616 6783 19668 6792
rect 19616 6749 19625 6783
rect 19625 6749 19659 6783
rect 19659 6749 19668 6783
rect 19616 6740 19668 6749
rect 19892 6740 19944 6792
rect 12808 6604 12860 6656
rect 13636 6604 13688 6656
rect 14648 6647 14700 6656
rect 14648 6613 14657 6647
rect 14657 6613 14691 6647
rect 14691 6613 14700 6647
rect 14648 6604 14700 6613
rect 15292 6604 15344 6656
rect 20720 6672 20772 6724
rect 21640 6672 21692 6724
rect 18512 6604 18564 6656
rect 20996 6604 21048 6656
rect 21456 6647 21508 6656
rect 21456 6613 21465 6647
rect 21465 6613 21499 6647
rect 21499 6613 21508 6647
rect 21456 6604 21508 6613
rect 21824 6783 21876 6792
rect 21824 6749 21833 6783
rect 21833 6749 21867 6783
rect 21867 6749 21876 6783
rect 21824 6740 21876 6749
rect 32680 6808 32732 6860
rect 33048 6808 33100 6860
rect 22008 6740 22060 6792
rect 22652 6783 22704 6792
rect 22652 6749 22661 6783
rect 22661 6749 22695 6783
rect 22695 6749 22704 6783
rect 22652 6740 22704 6749
rect 24032 6783 24084 6792
rect 24032 6749 24041 6783
rect 24041 6749 24075 6783
rect 24075 6749 24084 6783
rect 24032 6740 24084 6749
rect 24584 6783 24636 6792
rect 24584 6749 24593 6783
rect 24593 6749 24627 6783
rect 24627 6749 24636 6783
rect 24584 6740 24636 6749
rect 25596 6672 25648 6724
rect 30012 6740 30064 6792
rect 30748 6740 30800 6792
rect 33508 6740 33560 6792
rect 34428 6808 34480 6860
rect 33692 6740 33744 6792
rect 35256 6783 35308 6792
rect 35256 6749 35265 6783
rect 35265 6749 35299 6783
rect 35299 6749 35308 6783
rect 35256 6740 35308 6749
rect 35440 6783 35492 6792
rect 35440 6749 35447 6783
rect 35447 6749 35492 6783
rect 35440 6740 35492 6749
rect 35624 6808 35676 6860
rect 37464 6808 37516 6860
rect 40040 6944 40092 6996
rect 40224 6987 40276 6996
rect 40224 6953 40233 6987
rect 40233 6953 40267 6987
rect 40267 6953 40276 6987
rect 40224 6944 40276 6953
rect 43996 6944 44048 6996
rect 39856 6876 39908 6928
rect 40500 6876 40552 6928
rect 35900 6740 35952 6792
rect 29736 6672 29788 6724
rect 32588 6672 32640 6724
rect 33140 6672 33192 6724
rect 25228 6604 25280 6656
rect 27988 6647 28040 6656
rect 27988 6613 27997 6647
rect 27997 6613 28031 6647
rect 28031 6613 28040 6647
rect 27988 6604 28040 6613
rect 32772 6604 32824 6656
rect 33692 6604 33744 6656
rect 36084 6672 36136 6724
rect 38476 6783 38528 6792
rect 38476 6749 38485 6783
rect 38485 6749 38519 6783
rect 38519 6749 38528 6783
rect 38476 6740 38528 6749
rect 39948 6740 40000 6792
rect 38936 6715 38988 6724
rect 38936 6681 38945 6715
rect 38945 6681 38979 6715
rect 38979 6681 38988 6715
rect 38936 6672 38988 6681
rect 40132 6808 40184 6860
rect 40776 6808 40828 6860
rect 41236 6808 41288 6860
rect 40868 6783 40920 6792
rect 40868 6749 40877 6783
rect 40877 6749 40911 6783
rect 40911 6749 40920 6783
rect 40868 6740 40920 6749
rect 34152 6647 34204 6656
rect 34152 6613 34161 6647
rect 34161 6613 34195 6647
rect 34195 6613 34204 6647
rect 34152 6604 34204 6613
rect 34980 6604 35032 6656
rect 39672 6604 39724 6656
rect 40316 6672 40368 6724
rect 42616 6740 42668 6792
rect 40132 6604 40184 6656
rect 40408 6647 40460 6656
rect 40408 6613 40417 6647
rect 40417 6613 40451 6647
rect 40451 6613 40460 6647
rect 40408 6604 40460 6613
rect 40684 6604 40736 6656
rect 42248 6604 42300 6656
rect 11896 6502 11948 6554
rect 11960 6502 12012 6554
rect 12024 6502 12076 6554
rect 12088 6502 12140 6554
rect 12152 6502 12204 6554
rect 22843 6502 22895 6554
rect 22907 6502 22959 6554
rect 22971 6502 23023 6554
rect 23035 6502 23087 6554
rect 23099 6502 23151 6554
rect 33790 6502 33842 6554
rect 33854 6502 33906 6554
rect 33918 6502 33970 6554
rect 33982 6502 34034 6554
rect 34046 6502 34098 6554
rect 44737 6502 44789 6554
rect 44801 6502 44853 6554
rect 44865 6502 44917 6554
rect 44929 6502 44981 6554
rect 44993 6502 45045 6554
rect 2872 6443 2924 6452
rect 2872 6409 2881 6443
rect 2881 6409 2915 6443
rect 2915 6409 2924 6443
rect 2872 6400 2924 6409
rect 940 6264 992 6316
rect 2320 6307 2372 6316
rect 2320 6273 2329 6307
rect 2329 6273 2363 6307
rect 2363 6273 2372 6307
rect 2320 6264 2372 6273
rect 3332 6307 3384 6316
rect 3332 6273 3341 6307
rect 3341 6273 3375 6307
rect 3375 6273 3384 6307
rect 3332 6264 3384 6273
rect 6920 6332 6972 6384
rect 9312 6443 9364 6452
rect 9312 6409 9321 6443
rect 9321 6409 9355 6443
rect 9355 6409 9364 6443
rect 9312 6400 9364 6409
rect 11152 6443 11204 6452
rect 11152 6409 11161 6443
rect 11161 6409 11195 6443
rect 11195 6409 11204 6443
rect 11152 6400 11204 6409
rect 10508 6332 10560 6384
rect 12532 6400 12584 6452
rect 12624 6400 12676 6452
rect 13728 6400 13780 6452
rect 13176 6332 13228 6384
rect 7932 6307 7984 6316
rect 7932 6273 7941 6307
rect 7941 6273 7975 6307
rect 7975 6273 7984 6307
rect 7932 6264 7984 6273
rect 8668 6264 8720 6316
rect 9588 6264 9640 6316
rect 12072 6264 12124 6316
rect 13452 6332 13504 6384
rect 14280 6332 14332 6384
rect 14832 6375 14884 6384
rect 14832 6341 14841 6375
rect 14841 6341 14875 6375
rect 14875 6341 14884 6375
rect 14832 6332 14884 6341
rect 14924 6332 14976 6384
rect 19892 6400 19944 6452
rect 20812 6400 20864 6452
rect 20996 6400 21048 6452
rect 21916 6400 21968 6452
rect 22652 6400 22704 6452
rect 24032 6400 24084 6452
rect 25228 6443 25280 6452
rect 25228 6409 25237 6443
rect 25237 6409 25271 6443
rect 25271 6409 25280 6443
rect 25228 6400 25280 6409
rect 32864 6400 32916 6452
rect 34336 6400 34388 6452
rect 35440 6400 35492 6452
rect 38476 6400 38528 6452
rect 39488 6400 39540 6452
rect 40868 6400 40920 6452
rect 18420 6332 18472 6384
rect 18604 6332 18656 6384
rect 14096 6264 14148 6316
rect 18788 6264 18840 6316
rect 13360 6196 13412 6248
rect 17776 6239 17828 6248
rect 17776 6205 17785 6239
rect 17785 6205 17819 6239
rect 17819 6205 17828 6239
rect 17776 6196 17828 6205
rect 18328 6196 18380 6248
rect 18972 6239 19024 6248
rect 18972 6205 18981 6239
rect 18981 6205 19015 6239
rect 19015 6205 19024 6239
rect 18972 6196 19024 6205
rect 19156 6239 19208 6248
rect 19156 6205 19165 6239
rect 19165 6205 19199 6239
rect 19199 6205 19208 6239
rect 19156 6196 19208 6205
rect 19708 6307 19760 6316
rect 19708 6273 19717 6307
rect 19717 6273 19751 6307
rect 19751 6273 19760 6307
rect 19708 6264 19760 6273
rect 19892 6307 19944 6316
rect 19892 6273 19901 6307
rect 19901 6273 19935 6307
rect 19935 6273 19944 6307
rect 19892 6264 19944 6273
rect 19984 6307 20036 6316
rect 19984 6273 19993 6307
rect 19993 6273 20027 6307
rect 20027 6273 20036 6307
rect 19984 6264 20036 6273
rect 21456 6332 21508 6384
rect 21548 6264 21600 6316
rect 27988 6332 28040 6384
rect 27896 6264 27948 6316
rect 20352 6196 20404 6248
rect 21180 6196 21232 6248
rect 25320 6239 25372 6248
rect 25320 6205 25329 6239
rect 25329 6205 25363 6239
rect 25363 6205 25372 6239
rect 25320 6196 25372 6205
rect 11704 6128 11756 6180
rect 12532 6171 12584 6180
rect 12532 6137 12541 6171
rect 12541 6137 12575 6171
rect 12575 6137 12584 6171
rect 12532 6128 12584 6137
rect 12992 6171 13044 6180
rect 12992 6137 13001 6171
rect 13001 6137 13035 6171
rect 13035 6137 13044 6171
rect 12992 6128 13044 6137
rect 13176 6060 13228 6112
rect 14648 6128 14700 6180
rect 20812 6128 20864 6180
rect 20904 6128 20956 6180
rect 14096 6060 14148 6112
rect 14924 6060 14976 6112
rect 15292 6060 15344 6112
rect 16028 6060 16080 6112
rect 19248 6060 19300 6112
rect 19708 6060 19760 6112
rect 24400 6128 24452 6180
rect 26148 6196 26200 6248
rect 27988 6196 28040 6248
rect 26792 6128 26844 6180
rect 28172 6128 28224 6180
rect 31944 6196 31996 6248
rect 32220 6264 32272 6316
rect 33048 6307 33100 6316
rect 33048 6273 33057 6307
rect 33057 6273 33091 6307
rect 33091 6273 33100 6307
rect 33048 6264 33100 6273
rect 33140 6307 33192 6316
rect 33140 6273 33149 6307
rect 33149 6273 33183 6307
rect 33183 6273 33192 6307
rect 33140 6264 33192 6273
rect 33416 6307 33468 6316
rect 33416 6273 33425 6307
rect 33425 6273 33459 6307
rect 33459 6273 33468 6307
rect 33416 6264 33468 6273
rect 34060 6307 34112 6316
rect 34060 6273 34069 6307
rect 34069 6273 34103 6307
rect 34103 6273 34112 6307
rect 34060 6264 34112 6273
rect 32864 6128 32916 6180
rect 33968 6196 34020 6248
rect 34244 6264 34296 6316
rect 34336 6239 34388 6248
rect 34336 6205 34345 6239
rect 34345 6205 34379 6239
rect 34379 6205 34388 6239
rect 34336 6196 34388 6205
rect 34980 6307 35032 6316
rect 34980 6273 34989 6307
rect 34989 6273 35023 6307
rect 35023 6273 35032 6307
rect 34980 6264 35032 6273
rect 36268 6332 36320 6384
rect 38936 6332 38988 6384
rect 35900 6307 35952 6316
rect 35900 6273 35909 6307
rect 35909 6273 35943 6307
rect 35943 6273 35952 6307
rect 35900 6264 35952 6273
rect 36084 6307 36136 6316
rect 36084 6273 36093 6307
rect 36093 6273 36127 6307
rect 36127 6273 36136 6307
rect 36084 6264 36136 6273
rect 38936 6196 38988 6248
rect 39488 6307 39540 6316
rect 39488 6273 39497 6307
rect 39497 6273 39531 6307
rect 39531 6273 39540 6307
rect 39488 6264 39540 6273
rect 40224 6332 40276 6384
rect 40500 6332 40552 6384
rect 40040 6264 40092 6316
rect 42616 6307 42668 6316
rect 42616 6273 42625 6307
rect 42625 6273 42659 6307
rect 42659 6273 42668 6307
rect 42616 6264 42668 6273
rect 33324 6128 33376 6180
rect 26332 6060 26384 6112
rect 30104 6060 30156 6112
rect 32036 6060 32088 6112
rect 32680 6060 32732 6112
rect 35348 6103 35400 6112
rect 35348 6069 35357 6103
rect 35357 6069 35391 6103
rect 35391 6069 35400 6103
rect 35348 6060 35400 6069
rect 35992 6103 36044 6112
rect 35992 6069 36001 6103
rect 36001 6069 36035 6103
rect 36035 6069 36044 6103
rect 35992 6060 36044 6069
rect 39120 6103 39172 6112
rect 39120 6069 39129 6103
rect 39129 6069 39163 6103
rect 39163 6069 39172 6103
rect 39120 6060 39172 6069
rect 40592 6239 40644 6248
rect 40592 6205 40601 6239
rect 40601 6205 40635 6239
rect 40635 6205 40644 6239
rect 40592 6196 40644 6205
rect 40132 6060 40184 6112
rect 40224 6060 40276 6112
rect 6423 5958 6475 6010
rect 6487 5958 6539 6010
rect 6551 5958 6603 6010
rect 6615 5958 6667 6010
rect 6679 5958 6731 6010
rect 17370 5958 17422 6010
rect 17434 5958 17486 6010
rect 17498 5958 17550 6010
rect 17562 5958 17614 6010
rect 17626 5958 17678 6010
rect 28317 5958 28369 6010
rect 28381 5958 28433 6010
rect 28445 5958 28497 6010
rect 28509 5958 28561 6010
rect 28573 5958 28625 6010
rect 39264 5958 39316 6010
rect 39328 5958 39380 6010
rect 39392 5958 39444 6010
rect 39456 5958 39508 6010
rect 39520 5958 39572 6010
rect 3240 5899 3292 5908
rect 3240 5865 3249 5899
rect 3249 5865 3283 5899
rect 3283 5865 3292 5899
rect 3240 5856 3292 5865
rect 5264 5856 5316 5908
rect 9588 5856 9640 5908
rect 12256 5856 12308 5908
rect 12992 5856 13044 5908
rect 13728 5856 13780 5908
rect 14464 5899 14516 5908
rect 14464 5865 14473 5899
rect 14473 5865 14507 5899
rect 14507 5865 14516 5899
rect 14464 5856 14516 5865
rect 15292 5856 15344 5908
rect 12532 5788 12584 5840
rect 14188 5788 14240 5840
rect 3976 5763 4028 5772
rect 3976 5729 3985 5763
rect 3985 5729 4019 5763
rect 4019 5729 4028 5763
rect 3976 5720 4028 5729
rect 5816 5763 5868 5772
rect 5816 5729 5825 5763
rect 5825 5729 5859 5763
rect 5859 5729 5868 5763
rect 5816 5720 5868 5729
rect 13360 5720 13412 5772
rect 14648 5720 14700 5772
rect 17132 5720 17184 5772
rect 18420 5856 18472 5908
rect 20904 5856 20956 5908
rect 18328 5788 18380 5840
rect 19156 5788 19208 5840
rect 2136 5652 2188 5704
rect 5172 5652 5224 5704
rect 6000 5695 6052 5704
rect 6000 5661 6009 5695
rect 6009 5661 6043 5695
rect 6043 5661 6052 5695
rect 6000 5652 6052 5661
rect 9588 5695 9640 5704
rect 9588 5661 9597 5695
rect 9597 5661 9631 5695
rect 9631 5661 9640 5695
rect 9588 5652 9640 5661
rect 10048 5652 10100 5704
rect 10416 5695 10468 5704
rect 10416 5661 10425 5695
rect 10425 5661 10459 5695
rect 10459 5661 10468 5695
rect 10416 5652 10468 5661
rect 13176 5652 13228 5704
rect 14832 5652 14884 5704
rect 16028 5695 16080 5704
rect 16028 5661 16037 5695
rect 16037 5661 16071 5695
rect 16071 5661 16080 5695
rect 16028 5652 16080 5661
rect 18696 5695 18748 5704
rect 18696 5661 18705 5695
rect 18705 5661 18739 5695
rect 18739 5661 18748 5695
rect 18696 5652 18748 5661
rect 20352 5720 20404 5772
rect 21548 5856 21600 5908
rect 21916 5856 21968 5908
rect 24400 5856 24452 5908
rect 29736 5899 29788 5908
rect 29736 5865 29745 5899
rect 29745 5865 29779 5899
rect 29779 5865 29788 5899
rect 29736 5856 29788 5865
rect 31944 5856 31996 5908
rect 32496 5856 32548 5908
rect 33416 5856 33468 5908
rect 34152 5856 34204 5908
rect 34428 5856 34480 5908
rect 35900 5856 35952 5908
rect 27896 5788 27948 5840
rect 16764 5627 16816 5636
rect 16764 5593 16773 5627
rect 16773 5593 16807 5627
rect 16807 5593 16816 5627
rect 16764 5584 16816 5593
rect 20536 5695 20588 5704
rect 20536 5661 20545 5695
rect 20545 5661 20579 5695
rect 20579 5661 20588 5695
rect 20536 5652 20588 5661
rect 20628 5695 20680 5704
rect 20628 5661 20637 5695
rect 20637 5661 20671 5695
rect 20671 5661 20680 5695
rect 20628 5652 20680 5661
rect 20996 5652 21048 5704
rect 24584 5720 24636 5772
rect 26792 5763 26844 5772
rect 26792 5729 26801 5763
rect 26801 5729 26835 5763
rect 26835 5729 26844 5763
rect 26792 5720 26844 5729
rect 27988 5720 28040 5772
rect 30472 5720 30524 5772
rect 33600 5788 33652 5840
rect 33692 5788 33744 5840
rect 21916 5652 21968 5704
rect 26332 5695 26384 5704
rect 26332 5661 26341 5695
rect 26341 5661 26375 5695
rect 26375 5661 26384 5695
rect 26332 5652 26384 5661
rect 27436 5652 27488 5704
rect 30104 5695 30156 5704
rect 30104 5661 30113 5695
rect 30113 5661 30147 5695
rect 30147 5661 30156 5695
rect 30104 5652 30156 5661
rect 31944 5652 31996 5704
rect 32036 5695 32088 5704
rect 32036 5661 32045 5695
rect 32045 5661 32079 5695
rect 32079 5661 32088 5695
rect 32036 5652 32088 5661
rect 32220 5695 32272 5704
rect 32220 5661 32229 5695
rect 32229 5661 32263 5695
rect 32263 5661 32272 5695
rect 32220 5652 32272 5661
rect 32956 5652 33008 5704
rect 7748 5516 7800 5568
rect 9956 5559 10008 5568
rect 9956 5525 9965 5559
rect 9965 5525 9999 5559
rect 9999 5525 10008 5559
rect 9956 5516 10008 5525
rect 16580 5516 16632 5568
rect 20444 5516 20496 5568
rect 20996 5516 21048 5568
rect 21180 5516 21232 5568
rect 30196 5627 30248 5636
rect 30196 5593 30205 5627
rect 30205 5593 30239 5627
rect 30239 5593 30248 5627
rect 30196 5584 30248 5593
rect 35348 5720 35400 5772
rect 33692 5652 33744 5704
rect 28264 5516 28316 5568
rect 32128 5559 32180 5568
rect 32128 5525 32137 5559
rect 32137 5525 32171 5559
rect 32171 5525 32180 5559
rect 32128 5516 32180 5525
rect 32772 5516 32824 5568
rect 34060 5584 34112 5636
rect 34152 5584 34204 5636
rect 33968 5516 34020 5568
rect 39672 5856 39724 5908
rect 40132 5899 40184 5908
rect 40132 5865 40141 5899
rect 40141 5865 40175 5899
rect 40175 5865 40184 5899
rect 40132 5856 40184 5865
rect 40408 5856 40460 5908
rect 40500 5856 40552 5908
rect 40868 5856 40920 5908
rect 39028 5788 39080 5840
rect 40040 5788 40092 5840
rect 37464 5720 37516 5772
rect 40224 5720 40276 5772
rect 40316 5763 40368 5772
rect 40316 5729 40325 5763
rect 40325 5729 40359 5763
rect 40359 5729 40368 5763
rect 40316 5720 40368 5729
rect 40132 5652 40184 5704
rect 42248 5652 42300 5704
rect 44088 5695 44140 5704
rect 44088 5661 44097 5695
rect 44097 5661 44131 5695
rect 44131 5661 44140 5695
rect 44088 5652 44140 5661
rect 36084 5516 36136 5568
rect 37188 5584 37240 5636
rect 38016 5627 38068 5636
rect 38016 5593 38025 5627
rect 38025 5593 38059 5627
rect 38059 5593 38068 5627
rect 38016 5584 38068 5593
rect 38660 5584 38712 5636
rect 41144 5627 41196 5636
rect 41144 5593 41153 5627
rect 41153 5593 41187 5627
rect 41187 5593 41196 5627
rect 41144 5584 41196 5593
rect 36912 5559 36964 5568
rect 36912 5525 36921 5559
rect 36921 5525 36955 5559
rect 36955 5525 36964 5559
rect 36912 5516 36964 5525
rect 41052 5516 41104 5568
rect 45008 5516 45060 5568
rect 11896 5414 11948 5466
rect 11960 5414 12012 5466
rect 12024 5414 12076 5466
rect 12088 5414 12140 5466
rect 12152 5414 12204 5466
rect 22843 5414 22895 5466
rect 22907 5414 22959 5466
rect 22971 5414 23023 5466
rect 23035 5414 23087 5466
rect 23099 5414 23151 5466
rect 33790 5414 33842 5466
rect 33854 5414 33906 5466
rect 33918 5414 33970 5466
rect 33982 5414 34034 5466
rect 34046 5414 34098 5466
rect 44737 5414 44789 5466
rect 44801 5414 44853 5466
rect 44865 5414 44917 5466
rect 44929 5414 44981 5466
rect 44993 5414 45045 5466
rect 5356 5355 5408 5364
rect 5356 5321 5365 5355
rect 5365 5321 5399 5355
rect 5399 5321 5408 5355
rect 5356 5312 5408 5321
rect 14096 5312 14148 5364
rect 15476 5312 15528 5364
rect 3976 5219 4028 5228
rect 3976 5185 3985 5219
rect 3985 5185 4019 5219
rect 4019 5185 4028 5219
rect 3976 5176 4028 5185
rect 4252 5219 4304 5228
rect 940 5108 992 5160
rect 4252 5185 4286 5219
rect 4286 5185 4304 5219
rect 4252 5176 4304 5185
rect 9588 5244 9640 5296
rect 9312 5176 9364 5228
rect 12256 5219 12308 5228
rect 12256 5185 12265 5219
rect 12265 5185 12299 5219
rect 12299 5185 12308 5219
rect 12256 5176 12308 5185
rect 13084 5176 13136 5228
rect 14096 5219 14148 5228
rect 14096 5185 14105 5219
rect 14105 5185 14139 5219
rect 14139 5185 14148 5219
rect 14096 5176 14148 5185
rect 14740 5176 14792 5228
rect 17132 5244 17184 5296
rect 18420 5244 18472 5296
rect 18604 5355 18656 5364
rect 18604 5321 18613 5355
rect 18613 5321 18647 5355
rect 18647 5321 18656 5355
rect 18604 5312 18656 5321
rect 21824 5312 21876 5364
rect 24400 5355 24452 5364
rect 24400 5321 24409 5355
rect 24409 5321 24443 5355
rect 24443 5321 24452 5355
rect 24400 5312 24452 5321
rect 28172 5312 28224 5364
rect 31208 5312 31260 5364
rect 32864 5312 32916 5364
rect 34152 5312 34204 5364
rect 34612 5312 34664 5364
rect 35440 5312 35492 5364
rect 36912 5312 36964 5364
rect 39120 5312 39172 5364
rect 40500 5355 40552 5364
rect 40500 5321 40509 5355
rect 40509 5321 40543 5355
rect 40543 5321 40552 5355
rect 40500 5312 40552 5321
rect 40592 5312 40644 5364
rect 19248 5219 19300 5228
rect 19248 5185 19257 5219
rect 19257 5185 19291 5219
rect 19291 5185 19300 5219
rect 19248 5176 19300 5185
rect 20996 5219 21048 5228
rect 20996 5185 21005 5219
rect 21005 5185 21039 5219
rect 21039 5185 21048 5219
rect 20996 5176 21048 5185
rect 21180 5219 21232 5228
rect 21180 5185 21189 5219
rect 21189 5185 21223 5219
rect 21223 5185 21232 5219
rect 21180 5176 21232 5185
rect 14188 5151 14240 5160
rect 14188 5117 14197 5151
rect 14197 5117 14231 5151
rect 14231 5117 14240 5151
rect 14188 5108 14240 5117
rect 14648 5108 14700 5160
rect 13544 4972 13596 5024
rect 14280 5015 14332 5024
rect 14280 4981 14289 5015
rect 14289 4981 14323 5015
rect 14323 4981 14332 5015
rect 14280 4972 14332 4981
rect 15200 4972 15252 5024
rect 24584 5244 24636 5296
rect 28724 5244 28776 5296
rect 23296 5219 23348 5228
rect 23296 5185 23330 5219
rect 23330 5185 23348 5219
rect 23296 5176 23348 5185
rect 32128 5176 32180 5228
rect 32220 5108 32272 5160
rect 32680 5219 32732 5228
rect 32680 5185 32689 5219
rect 32689 5185 32723 5219
rect 32723 5185 32732 5219
rect 32680 5176 32732 5185
rect 32496 5040 32548 5092
rect 32864 5219 32916 5228
rect 32864 5185 32873 5219
rect 32873 5185 32907 5219
rect 32907 5185 32916 5219
rect 32864 5176 32916 5185
rect 33324 5176 33376 5228
rect 40132 5244 40184 5296
rect 40684 5244 40736 5296
rect 36268 5176 36320 5228
rect 37372 5176 37424 5228
rect 38660 5176 38712 5228
rect 39672 5176 39724 5228
rect 40776 5176 40828 5228
rect 41052 5219 41104 5228
rect 41052 5185 41061 5219
rect 41061 5185 41095 5219
rect 41095 5185 41104 5219
rect 41052 5176 41104 5185
rect 42984 5219 43036 5228
rect 42984 5185 42993 5219
rect 42993 5185 43027 5219
rect 43027 5185 43036 5219
rect 42984 5176 43036 5185
rect 35900 5040 35952 5092
rect 27344 4972 27396 5024
rect 31484 4972 31536 5024
rect 35992 4972 36044 5024
rect 41144 5040 41196 5092
rect 38844 5015 38896 5024
rect 38844 4981 38853 5015
rect 38853 4981 38887 5015
rect 38887 4981 38896 5015
rect 38844 4972 38896 4981
rect 44088 4972 44140 5024
rect 6423 4870 6475 4922
rect 6487 4870 6539 4922
rect 6551 4870 6603 4922
rect 6615 4870 6667 4922
rect 6679 4870 6731 4922
rect 17370 4870 17422 4922
rect 17434 4870 17486 4922
rect 17498 4870 17550 4922
rect 17562 4870 17614 4922
rect 17626 4870 17678 4922
rect 28317 4870 28369 4922
rect 28381 4870 28433 4922
rect 28445 4870 28497 4922
rect 28509 4870 28561 4922
rect 28573 4870 28625 4922
rect 39264 4870 39316 4922
rect 39328 4870 39380 4922
rect 39392 4870 39444 4922
rect 39456 4870 39508 4922
rect 39520 4870 39572 4922
rect 4252 4768 4304 4820
rect 13176 4811 13228 4820
rect 13176 4777 13185 4811
rect 13185 4777 13219 4811
rect 13219 4777 13228 4811
rect 13176 4768 13228 4777
rect 18420 4811 18472 4820
rect 18420 4777 18429 4811
rect 18429 4777 18463 4811
rect 18463 4777 18472 4811
rect 18420 4768 18472 4777
rect 18972 4700 19024 4752
rect 5816 4632 5868 4684
rect 20536 4675 20588 4684
rect 20536 4641 20545 4675
rect 20545 4641 20579 4675
rect 20579 4641 20588 4675
rect 20536 4632 20588 4641
rect 20812 4675 20864 4684
rect 20812 4641 20821 4675
rect 20821 4641 20855 4675
rect 20855 4641 20864 4675
rect 20812 4632 20864 4641
rect 5264 4564 5316 4616
rect 15200 4607 15252 4616
rect 15200 4573 15209 4607
rect 15209 4573 15243 4607
rect 15243 4573 15252 4607
rect 15200 4564 15252 4573
rect 15660 4607 15712 4616
rect 15660 4573 15669 4607
rect 15669 4573 15703 4607
rect 15703 4573 15712 4607
rect 15660 4564 15712 4573
rect 17960 4564 18012 4616
rect 18696 4564 18748 4616
rect 11612 4496 11664 4548
rect 12256 4496 12308 4548
rect 17132 4496 17184 4548
rect 17868 4496 17920 4548
rect 20720 4496 20772 4548
rect 22100 4496 22152 4548
rect 27804 4768 27856 4820
rect 33692 4768 33744 4820
rect 37188 4811 37240 4820
rect 37188 4777 37197 4811
rect 37197 4777 37231 4811
rect 37231 4777 37240 4811
rect 37188 4768 37240 4777
rect 38016 4768 38068 4820
rect 33140 4700 33192 4752
rect 33324 4700 33376 4752
rect 26792 4632 26844 4684
rect 31208 4675 31260 4684
rect 31208 4641 31217 4675
rect 31217 4641 31251 4675
rect 31251 4641 31260 4675
rect 31208 4632 31260 4641
rect 31484 4675 31536 4684
rect 31484 4641 31493 4675
rect 31493 4641 31527 4675
rect 31527 4641 31536 4675
rect 31484 4632 31536 4641
rect 35440 4675 35492 4684
rect 35440 4641 35449 4675
rect 35449 4641 35483 4675
rect 35483 4641 35492 4675
rect 35440 4632 35492 4641
rect 28172 4564 28224 4616
rect 32864 4564 32916 4616
rect 33876 4607 33928 4616
rect 33876 4573 33885 4607
rect 33885 4573 33919 4607
rect 33919 4573 33928 4607
rect 33876 4564 33928 4573
rect 37372 4564 37424 4616
rect 38844 4564 38896 4616
rect 44088 4607 44140 4616
rect 44088 4573 44097 4607
rect 44097 4573 44131 4607
rect 44131 4573 44140 4607
rect 44088 4564 44140 4573
rect 27896 4496 27948 4548
rect 33508 4496 33560 4548
rect 35072 4496 35124 4548
rect 5908 4428 5960 4480
rect 14832 4428 14884 4480
rect 19432 4428 19484 4480
rect 23204 4471 23256 4480
rect 23204 4437 23213 4471
rect 23213 4437 23247 4471
rect 23247 4437 23256 4471
rect 23204 4428 23256 4437
rect 33140 4428 33192 4480
rect 44272 4471 44324 4480
rect 44272 4437 44281 4471
rect 44281 4437 44315 4471
rect 44315 4437 44324 4471
rect 44272 4428 44324 4437
rect 11896 4326 11948 4378
rect 11960 4326 12012 4378
rect 12024 4326 12076 4378
rect 12088 4326 12140 4378
rect 12152 4326 12204 4378
rect 22843 4326 22895 4378
rect 22907 4326 22959 4378
rect 22971 4326 23023 4378
rect 23035 4326 23087 4378
rect 23099 4326 23151 4378
rect 33790 4326 33842 4378
rect 33854 4326 33906 4378
rect 33918 4326 33970 4378
rect 33982 4326 34034 4378
rect 34046 4326 34098 4378
rect 44737 4326 44789 4378
rect 44801 4326 44853 4378
rect 44865 4326 44917 4378
rect 44929 4326 44981 4378
rect 44993 4326 45045 4378
rect 13084 4267 13136 4276
rect 13084 4233 13093 4267
rect 13093 4233 13127 4267
rect 13127 4233 13136 4267
rect 13084 4224 13136 4233
rect 13544 4224 13596 4276
rect 42984 4224 43036 4276
rect 14832 4199 14884 4208
rect 14832 4165 14841 4199
rect 14841 4165 14875 4199
rect 14875 4165 14884 4199
rect 14832 4156 14884 4165
rect 17592 4156 17644 4208
rect 19432 4156 19484 4208
rect 20720 4156 20772 4208
rect 14280 4020 14332 4072
rect 16764 4088 16816 4140
rect 17960 4088 18012 4140
rect 23940 4156 23992 4208
rect 27804 4199 27856 4208
rect 27804 4165 27813 4199
rect 27813 4165 27847 4199
rect 27847 4165 27856 4199
rect 27804 4156 27856 4165
rect 22100 4131 22152 4140
rect 22100 4097 22109 4131
rect 22109 4097 22143 4131
rect 22143 4097 22152 4131
rect 22100 4088 22152 4097
rect 23204 4088 23256 4140
rect 27896 4131 27948 4140
rect 27896 4097 27905 4131
rect 27905 4097 27939 4131
rect 27939 4097 27948 4131
rect 27896 4088 27948 4097
rect 14556 4063 14608 4072
rect 14556 4029 14565 4063
rect 14565 4029 14599 4063
rect 14599 4029 14608 4063
rect 14556 4020 14608 4029
rect 15292 4020 15344 4072
rect 17868 4020 17920 4072
rect 20812 4020 20864 4072
rect 27988 4063 28040 4072
rect 27988 4029 27997 4063
rect 27997 4029 28031 4063
rect 28031 4029 28040 4063
rect 27988 4020 28040 4029
rect 23296 3952 23348 4004
rect 27436 3995 27488 4004
rect 27436 3961 27445 3995
rect 27445 3961 27479 3995
rect 27479 3961 27488 3995
rect 27436 3952 27488 3961
rect 15844 3884 15896 3936
rect 17592 3927 17644 3936
rect 17592 3893 17601 3927
rect 17601 3893 17635 3927
rect 17635 3893 17644 3927
rect 17592 3884 17644 3893
rect 23756 3884 23808 3936
rect 31024 3884 31076 3936
rect 33140 4088 33192 4140
rect 38200 4156 38252 4208
rect 32128 4020 32180 4072
rect 33508 4131 33560 4140
rect 33508 4097 33517 4131
rect 33517 4097 33551 4131
rect 33551 4097 33560 4131
rect 33508 4088 33560 4097
rect 35900 4088 35952 4140
rect 36360 4131 36412 4140
rect 36360 4097 36369 4131
rect 36369 4097 36403 4131
rect 36403 4097 36412 4131
rect 36360 4088 36412 4097
rect 31944 3952 31996 4004
rect 32864 3952 32916 4004
rect 35072 3995 35124 4004
rect 35072 3961 35081 3995
rect 35081 3961 35115 3995
rect 35115 3961 35124 3995
rect 35072 3952 35124 3961
rect 36268 4063 36320 4072
rect 36268 4029 36277 4063
rect 36277 4029 36311 4063
rect 36311 4029 36320 4063
rect 36268 4020 36320 4029
rect 37372 4088 37424 4140
rect 37464 4131 37516 4140
rect 37464 4097 37473 4131
rect 37473 4097 37507 4131
rect 37507 4097 37516 4131
rect 37464 4088 37516 4097
rect 31668 3927 31720 3936
rect 31668 3893 31677 3927
rect 31677 3893 31711 3927
rect 31711 3893 31720 3927
rect 31668 3884 31720 3893
rect 32036 3884 32088 3936
rect 36360 3884 36412 3936
rect 44088 3884 44140 3936
rect 6423 3782 6475 3834
rect 6487 3782 6539 3834
rect 6551 3782 6603 3834
rect 6615 3782 6667 3834
rect 6679 3782 6731 3834
rect 17370 3782 17422 3834
rect 17434 3782 17486 3834
rect 17498 3782 17550 3834
rect 17562 3782 17614 3834
rect 17626 3782 17678 3834
rect 28317 3782 28369 3834
rect 28381 3782 28433 3834
rect 28445 3782 28497 3834
rect 28509 3782 28561 3834
rect 28573 3782 28625 3834
rect 39264 3782 39316 3834
rect 39328 3782 39380 3834
rect 39392 3782 39444 3834
rect 39456 3782 39508 3834
rect 39520 3782 39572 3834
rect 9956 3680 10008 3732
rect 26884 3680 26936 3732
rect 32036 3680 32088 3732
rect 32864 3723 32916 3732
rect 32864 3689 32873 3723
rect 32873 3689 32907 3723
rect 32907 3689 32916 3723
rect 32864 3680 32916 3689
rect 38200 3680 38252 3732
rect 23756 3612 23808 3664
rect 23388 3544 23440 3596
rect 33508 3544 33560 3596
rect 940 3476 992 3528
rect 5908 3519 5960 3528
rect 5908 3485 5917 3519
rect 5917 3485 5951 3519
rect 5951 3485 5960 3519
rect 5908 3476 5960 3485
rect 14556 3519 14608 3528
rect 14556 3485 14565 3519
rect 14565 3485 14599 3519
rect 14599 3485 14608 3519
rect 14556 3476 14608 3485
rect 14832 3476 14884 3528
rect 16948 3476 17000 3528
rect 17040 3519 17092 3528
rect 17040 3485 17049 3519
rect 17049 3485 17083 3519
rect 17083 3485 17092 3519
rect 17040 3476 17092 3485
rect 17868 3476 17920 3528
rect 20536 3476 20588 3528
rect 31116 3519 31168 3528
rect 31116 3485 31125 3519
rect 31125 3485 31159 3519
rect 31159 3485 31168 3519
rect 31116 3476 31168 3485
rect 37372 3476 37424 3528
rect 44640 3476 44692 3528
rect 16580 3408 16632 3460
rect 5724 3383 5776 3392
rect 5724 3349 5733 3383
rect 5733 3349 5767 3383
rect 5767 3349 5776 3383
rect 5724 3340 5776 3349
rect 14464 3340 14516 3392
rect 17040 3340 17092 3392
rect 18880 3408 18932 3460
rect 22100 3451 22152 3460
rect 22100 3417 22109 3451
rect 22109 3417 22143 3451
rect 22143 3417 22152 3451
rect 22100 3408 22152 3417
rect 31668 3408 31720 3460
rect 18604 3340 18656 3392
rect 30288 3340 30340 3392
rect 36360 3408 36412 3460
rect 11896 3238 11948 3290
rect 11960 3238 12012 3290
rect 12024 3238 12076 3290
rect 12088 3238 12140 3290
rect 12152 3238 12204 3290
rect 22843 3238 22895 3290
rect 22907 3238 22959 3290
rect 22971 3238 23023 3290
rect 23035 3238 23087 3290
rect 23099 3238 23151 3290
rect 33790 3238 33842 3290
rect 33854 3238 33906 3290
rect 33918 3238 33970 3290
rect 33982 3238 34034 3290
rect 34046 3238 34098 3290
rect 44737 3238 44789 3290
rect 44801 3238 44853 3290
rect 44865 3238 44917 3290
rect 44929 3238 44981 3290
rect 44993 3238 45045 3290
rect 7748 3043 7800 3052
rect 7748 3009 7757 3043
rect 7757 3009 7791 3043
rect 7791 3009 7800 3043
rect 7748 3000 7800 3009
rect 9404 3000 9456 3052
rect 16856 3136 16908 3188
rect 16948 3179 17000 3188
rect 16948 3145 16957 3179
rect 16957 3145 16991 3179
rect 16991 3145 17000 3179
rect 16948 3136 17000 3145
rect 15844 3068 15896 3120
rect 16580 3068 16632 3120
rect 14464 3043 14516 3052
rect 14464 3009 14473 3043
rect 14473 3009 14507 3043
rect 14507 3009 14516 3043
rect 14464 3000 14516 3009
rect 14832 3043 14884 3052
rect 14832 3009 14841 3043
rect 14841 3009 14875 3043
rect 14875 3009 14884 3043
rect 14832 3000 14884 3009
rect 17868 3068 17920 3120
rect 22100 3136 22152 3188
rect 26884 3136 26936 3188
rect 16764 2932 16816 2984
rect 18604 3000 18656 3052
rect 18880 3043 18932 3052
rect 18880 3009 18889 3043
rect 18889 3009 18923 3043
rect 18923 3009 18932 3043
rect 18880 3000 18932 3009
rect 22468 3043 22520 3052
rect 22468 3009 22477 3043
rect 22477 3009 22511 3043
rect 22511 3009 22520 3043
rect 22468 3000 22520 3009
rect 44456 3136 44508 3188
rect 45100 3000 45152 3052
rect 940 2796 992 2848
rect 9588 2796 9640 2848
rect 14188 2796 14240 2848
rect 22652 2796 22704 2848
rect 35532 2796 35584 2848
rect 6423 2694 6475 2746
rect 6487 2694 6539 2746
rect 6551 2694 6603 2746
rect 6615 2694 6667 2746
rect 6679 2694 6731 2746
rect 17370 2694 17422 2746
rect 17434 2694 17486 2746
rect 17498 2694 17550 2746
rect 17562 2694 17614 2746
rect 17626 2694 17678 2746
rect 28317 2694 28369 2746
rect 28381 2694 28433 2746
rect 28445 2694 28497 2746
rect 28509 2694 28561 2746
rect 28573 2694 28625 2746
rect 39264 2694 39316 2746
rect 39328 2694 39380 2746
rect 39392 2694 39444 2746
rect 39456 2694 39508 2746
rect 39520 2694 39572 2746
rect 17132 2592 17184 2644
rect 27344 2635 27396 2644
rect 27344 2601 27353 2635
rect 27353 2601 27387 2635
rect 27387 2601 27396 2635
rect 27344 2592 27396 2601
rect 38108 2592 38160 2644
rect 43444 2635 43496 2644
rect 43444 2601 43453 2635
rect 43453 2601 43487 2635
rect 43487 2601 43496 2635
rect 43444 2592 43496 2601
rect 30196 2524 30248 2576
rect 20 2456 72 2508
rect 12808 2456 12860 2508
rect 1308 2388 1360 2440
rect 4160 2431 4212 2440
rect 4160 2397 4169 2431
rect 4169 2397 4203 2431
rect 4203 2397 4212 2431
rect 4160 2388 4212 2397
rect 4528 2388 4580 2440
rect 5724 2388 5776 2440
rect 7748 2388 7800 2440
rect 9588 2388 9640 2440
rect 11060 2388 11112 2440
rect 12900 2431 12952 2440
rect 12900 2397 12909 2431
rect 12909 2397 12943 2431
rect 12943 2397 12952 2431
rect 12900 2388 12952 2397
rect 16120 2388 16172 2440
rect 16764 2388 16816 2440
rect 32588 2499 32640 2508
rect 32588 2465 32597 2499
rect 32597 2465 32631 2499
rect 32631 2465 32640 2499
rect 32588 2456 32640 2465
rect 17408 2388 17460 2440
rect 19340 2388 19392 2440
rect 20720 2388 20772 2440
rect 22652 2431 22704 2440
rect 22652 2397 22661 2431
rect 22661 2397 22695 2431
rect 22695 2397 22704 2431
rect 22652 2388 22704 2397
rect 23848 2388 23900 2440
rect 25780 2388 25832 2440
rect 27068 2388 27120 2440
rect 29000 2388 29052 2440
rect 30380 2388 30432 2440
rect 32220 2388 32272 2440
rect 35532 2431 35584 2440
rect 35532 2397 35541 2431
rect 35541 2397 35575 2431
rect 35575 2397 35584 2431
rect 35532 2388 35584 2397
rect 37648 2431 37700 2440
rect 37648 2397 37657 2431
rect 37657 2397 37691 2431
rect 37691 2397 37700 2431
rect 37648 2388 37700 2397
rect 38660 2388 38712 2440
rect 40040 2388 40092 2440
rect 43812 2388 43864 2440
rect 44088 2431 44140 2440
rect 44088 2397 44097 2431
rect 44097 2397 44131 2431
rect 44131 2397 44140 2431
rect 44088 2388 44140 2397
rect 41880 2320 41932 2372
rect 6460 2252 6512 2304
rect 9680 2252 9732 2304
rect 22560 2252 22612 2304
rect 31852 2252 31904 2304
rect 35440 2252 35492 2304
rect 44272 2295 44324 2304
rect 44272 2261 44281 2295
rect 44281 2261 44315 2295
rect 44315 2261 44324 2295
rect 44272 2252 44324 2261
rect 11896 2150 11948 2202
rect 11960 2150 12012 2202
rect 12024 2150 12076 2202
rect 12088 2150 12140 2202
rect 12152 2150 12204 2202
rect 22843 2150 22895 2202
rect 22907 2150 22959 2202
rect 22971 2150 23023 2202
rect 23035 2150 23087 2202
rect 23099 2150 23151 2202
rect 33790 2150 33842 2202
rect 33854 2150 33906 2202
rect 33918 2150 33970 2202
rect 33982 2150 34034 2202
rect 34046 2150 34098 2202
rect 44737 2150 44789 2202
rect 44801 2150 44853 2202
rect 44865 2150 44917 2202
rect 44929 2150 44981 2202
rect 44993 2150 45045 2202
rect 3240 892 3292 944
rect 4160 892 4212 944
rect 36728 892 36780 944
rect 37648 892 37700 944
<< metal2 >>
rect -10 19200 102 20000
rect 1278 19200 1390 20000
rect 3210 19200 3322 20000
rect 4498 19200 4610 20000
rect 6430 19200 6542 20000
rect 7718 19200 7830 20000
rect 9650 19200 9762 20000
rect 10938 19200 11050 20000
rect 12870 19200 12982 20000
rect 14158 19200 14270 20000
rect 16090 19200 16202 20000
rect 17378 19200 17490 20000
rect 19310 19200 19422 20000
rect 20598 19200 20710 20000
rect 22530 19200 22642 20000
rect 23818 19200 23930 20000
rect 25750 19200 25862 20000
rect 27682 19200 27794 20000
rect 28970 19200 29082 20000
rect 30902 19200 31014 20000
rect 32190 19200 32302 20000
rect 34122 19200 34234 20000
rect 35410 19200 35522 20000
rect 37342 19200 37454 20000
rect 38630 19200 38742 20000
rect 40562 19200 40674 20000
rect 41850 19200 41962 20000
rect 43782 19200 43894 20000
rect 45070 19200 45182 20000
rect 32 16590 60 19200
rect 1030 18456 1086 18465
rect 1030 18391 1086 18400
rect 940 17196 992 17202
rect 940 17138 992 17144
rect 952 17105 980 17138
rect 938 17096 994 17105
rect 938 17031 994 17040
rect 20 16584 72 16590
rect 20 16526 72 16532
rect 1044 16114 1072 18391
rect 1320 17270 1348 19200
rect 3252 17270 3280 19200
rect 4540 17270 4568 19200
rect 1308 17264 1360 17270
rect 1308 17206 1360 17212
rect 3240 17264 3292 17270
rect 3240 17206 3292 17212
rect 4528 17264 4580 17270
rect 4528 17206 4580 17212
rect 6472 17202 6500 19200
rect 7760 17202 7788 19200
rect 9692 17202 9720 19200
rect 10980 19122 11008 19200
rect 10980 19094 11100 19122
rect 11072 17270 11100 19094
rect 11896 17436 12204 17445
rect 11896 17434 11902 17436
rect 11958 17434 11982 17436
rect 12038 17434 12062 17436
rect 12118 17434 12142 17436
rect 12198 17434 12204 17436
rect 11958 17382 11960 17434
rect 12140 17382 12142 17434
rect 11896 17380 11902 17382
rect 11958 17380 11982 17382
rect 12038 17380 12062 17382
rect 12118 17380 12142 17382
rect 12198 17380 12204 17382
rect 11896 17371 12204 17380
rect 11060 17264 11112 17270
rect 11060 17206 11112 17212
rect 12912 17202 12940 19200
rect 14200 17202 14228 19200
rect 16132 17270 16160 19200
rect 17420 17338 17448 19200
rect 17408 17332 17460 17338
rect 17408 17274 17460 17280
rect 16120 17264 16172 17270
rect 16120 17206 16172 17212
rect 19352 17202 19380 19200
rect 20640 19122 20668 19200
rect 20640 19094 20760 19122
rect 20732 17338 20760 19094
rect 20720 17332 20772 17338
rect 20720 17274 20772 17280
rect 22572 17202 22600 19200
rect 22843 17436 23151 17445
rect 22843 17434 22849 17436
rect 22905 17434 22929 17436
rect 22985 17434 23009 17436
rect 23065 17434 23089 17436
rect 23145 17434 23151 17436
rect 22905 17382 22907 17434
rect 23087 17382 23089 17434
rect 22843 17380 22849 17382
rect 22905 17380 22929 17382
rect 22985 17380 23009 17382
rect 23065 17380 23089 17382
rect 23145 17380 23151 17382
rect 22843 17371 23151 17380
rect 23860 17202 23888 19200
rect 25792 17202 25820 19200
rect 27724 17202 27752 19200
rect 29012 17202 29040 19200
rect 30944 17202 30972 19200
rect 32232 17270 32260 19200
rect 34164 19106 34192 19200
rect 34152 19100 34204 19106
rect 34152 19042 34204 19048
rect 35072 19100 35124 19106
rect 35072 19042 35124 19048
rect 33790 17436 34098 17445
rect 33790 17434 33796 17436
rect 33852 17434 33876 17436
rect 33932 17434 33956 17436
rect 34012 17434 34036 17436
rect 34092 17434 34098 17436
rect 33852 17382 33854 17434
rect 34034 17382 34036 17434
rect 33790 17380 33796 17382
rect 33852 17380 33876 17382
rect 33932 17380 33956 17382
rect 34012 17380 34036 17382
rect 34092 17380 34098 17382
rect 33790 17371 34098 17380
rect 32220 17264 32272 17270
rect 32220 17206 32272 17212
rect 35084 17202 35112 19042
rect 35452 17202 35480 19200
rect 37384 17202 37412 19200
rect 38672 17270 38700 19200
rect 40604 17338 40632 19200
rect 41892 19106 41920 19200
rect 41880 19100 41932 19106
rect 41880 19042 41932 19048
rect 42800 19100 42852 19106
rect 42800 19042 42852 19048
rect 40592 17332 40644 17338
rect 40592 17274 40644 17280
rect 38660 17264 38712 17270
rect 38660 17206 38712 17212
rect 42812 17202 42840 19042
rect 43720 18012 43772 18018
rect 43720 17954 43772 17960
rect 6460 17196 6512 17202
rect 6460 17138 6512 17144
rect 7748 17196 7800 17202
rect 7748 17138 7800 17144
rect 9680 17196 9732 17202
rect 9680 17138 9732 17144
rect 12900 17196 12952 17202
rect 12900 17138 12952 17144
rect 14188 17196 14240 17202
rect 14188 17138 14240 17144
rect 16580 17196 16632 17202
rect 16580 17138 16632 17144
rect 19340 17196 19392 17202
rect 19340 17138 19392 17144
rect 20720 17196 20772 17202
rect 20720 17138 20772 17144
rect 22560 17196 22612 17202
rect 22560 17138 22612 17144
rect 23848 17196 23900 17202
rect 23848 17138 23900 17144
rect 25780 17196 25832 17202
rect 25780 17138 25832 17144
rect 27712 17196 27764 17202
rect 27712 17138 27764 17144
rect 29000 17196 29052 17202
rect 29000 17138 29052 17144
rect 30932 17196 30984 17202
rect 30932 17138 30984 17144
rect 35072 17196 35124 17202
rect 35072 17138 35124 17144
rect 35440 17196 35492 17202
rect 35440 17138 35492 17144
rect 37372 17196 37424 17202
rect 37372 17138 37424 17144
rect 40684 17196 40736 17202
rect 40684 17138 40736 17144
rect 42800 17196 42852 17202
rect 42800 17138 42852 17144
rect 1860 17060 1912 17066
rect 1860 17002 1912 17008
rect 4068 17060 4120 17066
rect 4068 17002 4120 17008
rect 13084 17060 13136 17066
rect 13084 17002 13136 17008
rect 16304 17060 16356 17066
rect 16304 17002 16356 17008
rect 1032 16108 1084 16114
rect 1032 16050 1084 16056
rect 940 15360 992 15366
rect 940 15302 992 15308
rect 952 15065 980 15302
rect 938 15056 994 15065
rect 938 14991 994 15000
rect 940 13864 992 13870
rect 940 13806 992 13812
rect 952 13705 980 13806
rect 1872 13802 1900 17002
rect 2504 16992 2556 16998
rect 2504 16934 2556 16940
rect 2516 16794 2544 16934
rect 2504 16788 2556 16794
rect 2504 16730 2556 16736
rect 1952 16652 2004 16658
rect 1952 16594 2004 16600
rect 1964 14618 1992 16594
rect 2964 15496 3016 15502
rect 2964 15438 3016 15444
rect 1952 14612 2004 14618
rect 1952 14554 2004 14560
rect 1860 13796 1912 13802
rect 1860 13738 1912 13744
rect 938 13696 994 13705
rect 938 13631 994 13640
rect 1964 10674 1992 14554
rect 2780 12640 2832 12646
rect 2780 12582 2832 12588
rect 1952 10668 2004 10674
rect 1952 10610 2004 10616
rect 938 10296 994 10305
rect 938 10231 940 10240
rect 992 10231 994 10240
rect 940 10202 992 10208
rect 2792 10062 2820 12582
rect 2976 12442 3004 15438
rect 3146 12880 3202 12889
rect 3146 12815 3148 12824
rect 3200 12815 3202 12824
rect 3976 12844 4028 12850
rect 3148 12786 3200 12792
rect 3976 12786 4028 12792
rect 2964 12436 3016 12442
rect 2964 12378 3016 12384
rect 3424 12232 3476 12238
rect 3424 12174 3476 12180
rect 3436 11354 3464 12174
rect 3988 11778 4016 12786
rect 4080 11937 4108 17002
rect 4804 16992 4856 16998
rect 4804 16934 4856 16940
rect 9956 16992 10008 16998
rect 9956 16934 10008 16940
rect 4816 12850 4844 16934
rect 6423 16892 6731 16901
rect 6423 16890 6429 16892
rect 6485 16890 6509 16892
rect 6565 16890 6589 16892
rect 6645 16890 6669 16892
rect 6725 16890 6731 16892
rect 6485 16838 6487 16890
rect 6667 16838 6669 16890
rect 6423 16836 6429 16838
rect 6485 16836 6509 16838
rect 6565 16836 6589 16838
rect 6645 16836 6669 16838
rect 6725 16836 6731 16838
rect 6423 16827 6731 16836
rect 6828 15904 6880 15910
rect 6828 15846 6880 15852
rect 6423 15804 6731 15813
rect 6423 15802 6429 15804
rect 6485 15802 6509 15804
rect 6565 15802 6589 15804
rect 6645 15802 6669 15804
rect 6725 15802 6731 15804
rect 6485 15750 6487 15802
rect 6667 15750 6669 15802
rect 6423 15748 6429 15750
rect 6485 15748 6509 15750
rect 6565 15748 6589 15750
rect 6645 15748 6669 15750
rect 6725 15748 6731 15750
rect 6423 15739 6731 15748
rect 6423 14716 6731 14725
rect 6423 14714 6429 14716
rect 6485 14714 6509 14716
rect 6565 14714 6589 14716
rect 6645 14714 6669 14716
rect 6725 14714 6731 14716
rect 6485 14662 6487 14714
rect 6667 14662 6669 14714
rect 6423 14660 6429 14662
rect 6485 14660 6509 14662
rect 6565 14660 6589 14662
rect 6645 14660 6669 14662
rect 6725 14660 6731 14662
rect 6423 14651 6731 14660
rect 6840 14074 6868 15846
rect 9968 14414 9996 16934
rect 11896 16348 12204 16357
rect 11896 16346 11902 16348
rect 11958 16346 11982 16348
rect 12038 16346 12062 16348
rect 12118 16346 12142 16348
rect 12198 16346 12204 16348
rect 11958 16294 11960 16346
rect 12140 16294 12142 16346
rect 11896 16292 11902 16294
rect 11958 16292 11982 16294
rect 12038 16292 12062 16294
rect 12118 16292 12142 16294
rect 12198 16292 12204 16294
rect 11896 16283 12204 16292
rect 11896 15260 12204 15269
rect 11896 15258 11902 15260
rect 11958 15258 11982 15260
rect 12038 15258 12062 15260
rect 12118 15258 12142 15260
rect 12198 15258 12204 15260
rect 11958 15206 11960 15258
rect 12140 15206 12142 15258
rect 11896 15204 11902 15206
rect 11958 15204 11982 15206
rect 12038 15204 12062 15206
rect 12118 15204 12142 15206
rect 12198 15204 12204 15206
rect 11896 15195 12204 15204
rect 9864 14408 9916 14414
rect 9864 14350 9916 14356
rect 9956 14408 10008 14414
rect 9956 14350 10008 14356
rect 6828 14068 6880 14074
rect 6828 14010 6880 14016
rect 5540 14000 5592 14006
rect 5540 13942 5592 13948
rect 5356 13932 5408 13938
rect 5356 13874 5408 13880
rect 5080 13320 5132 13326
rect 5080 13262 5132 13268
rect 4344 12844 4396 12850
rect 4344 12786 4396 12792
rect 4804 12844 4856 12850
rect 4804 12786 4856 12792
rect 4356 12434 4384 12786
rect 5092 12782 5120 13262
rect 5368 12986 5396 13874
rect 5356 12980 5408 12986
rect 5356 12922 5408 12928
rect 5080 12776 5132 12782
rect 5080 12718 5132 12724
rect 4356 12406 4476 12434
rect 4252 12096 4304 12102
rect 4252 12038 4304 12044
rect 4066 11928 4122 11937
rect 4066 11863 4122 11872
rect 3988 11750 4200 11778
rect 4264 11762 4292 12038
rect 4066 11656 4122 11665
rect 4172 11626 4200 11750
rect 4252 11756 4304 11762
rect 4252 11698 4304 11704
rect 4066 11591 4122 11600
rect 4160 11620 4212 11626
rect 4080 11558 4108 11591
rect 4160 11562 4212 11568
rect 3976 11552 4028 11558
rect 3976 11494 4028 11500
rect 4068 11552 4120 11558
rect 4068 11494 4120 11500
rect 3424 11348 3476 11354
rect 3424 11290 3476 11296
rect 3988 11218 4016 11494
rect 3976 11212 4028 11218
rect 3976 11154 4028 11160
rect 4172 11150 4200 11562
rect 3148 11144 3200 11150
rect 3148 11086 3200 11092
rect 3240 11144 3292 11150
rect 4160 11144 4212 11150
rect 3240 11086 3292 11092
rect 4080 11092 4160 11098
rect 4080 11086 4212 11092
rect 3160 10742 3188 11086
rect 3148 10736 3200 10742
rect 3148 10678 3200 10684
rect 3148 10464 3200 10470
rect 3148 10406 3200 10412
rect 3160 10130 3188 10406
rect 3148 10124 3200 10130
rect 3148 10066 3200 10072
rect 2780 10056 2832 10062
rect 2780 9998 2832 10004
rect 2228 9920 2280 9926
rect 2228 9862 2280 9868
rect 2240 9586 2268 9862
rect 2228 9580 2280 9586
rect 2228 9522 2280 9528
rect 2044 9376 2096 9382
rect 2044 9318 2096 9324
rect 2056 8634 2084 9318
rect 3252 8906 3280 11086
rect 4080 11070 4200 11086
rect 4080 10674 4108 11070
rect 4068 10668 4120 10674
rect 4068 10610 4120 10616
rect 4252 10668 4304 10674
rect 4252 10610 4304 10616
rect 3424 10124 3476 10130
rect 3424 10066 3476 10072
rect 3332 10056 3384 10062
rect 3332 9998 3384 10004
rect 3344 9586 3372 9998
rect 3332 9580 3384 9586
rect 3332 9522 3384 9528
rect 3240 8900 3292 8906
rect 3240 8842 3292 8848
rect 2228 8832 2280 8838
rect 2228 8774 2280 8780
rect 2044 8628 2096 8634
rect 2044 8570 2096 8576
rect 2240 8498 2268 8774
rect 2228 8492 2280 8498
rect 2228 8434 2280 8440
rect 3252 8362 3280 8842
rect 3240 8356 3292 8362
rect 3240 8298 3292 8304
rect 938 8256 994 8265
rect 938 8191 994 8200
rect 952 7410 980 8191
rect 3344 7954 3372 9522
rect 3436 9042 3464 10066
rect 4264 9382 4292 10610
rect 4344 9920 4396 9926
rect 4344 9862 4396 9868
rect 4252 9376 4304 9382
rect 4252 9318 4304 9324
rect 3424 9036 3476 9042
rect 3424 8978 3476 8984
rect 3332 7948 3384 7954
rect 3332 7890 3384 7896
rect 2320 7812 2372 7818
rect 2320 7754 2372 7760
rect 940 7404 992 7410
rect 940 7346 992 7352
rect 938 6896 994 6905
rect 938 6831 994 6840
rect 952 6322 980 6831
rect 2136 6656 2188 6662
rect 2136 6598 2188 6604
rect 940 6316 992 6322
rect 940 6258 992 6264
rect 2148 5710 2176 6598
rect 2332 6322 2360 7754
rect 3240 6724 3292 6730
rect 3240 6666 3292 6672
rect 2872 6656 2924 6662
rect 2872 6598 2924 6604
rect 2884 6458 2912 6598
rect 2872 6452 2924 6458
rect 2872 6394 2924 6400
rect 2320 6316 2372 6322
rect 2320 6258 2372 6264
rect 3252 5914 3280 6666
rect 3344 6322 3372 7890
rect 3436 6866 3464 8978
rect 4356 8634 4384 9862
rect 4344 8628 4396 8634
rect 4344 8570 4396 8576
rect 3976 8492 4028 8498
rect 3976 8434 4028 8440
rect 3884 7948 3936 7954
rect 3884 7890 3936 7896
rect 3896 7546 3924 7890
rect 3884 7540 3936 7546
rect 3884 7482 3936 7488
rect 3988 6866 4016 8434
rect 4448 7818 4476 12406
rect 5092 12238 5120 12718
rect 5080 12232 5132 12238
rect 5080 12174 5132 12180
rect 4620 12096 4672 12102
rect 4620 12038 4672 12044
rect 4528 11824 4580 11830
rect 4528 11766 4580 11772
rect 4540 9450 4568 11766
rect 4632 10810 4660 12038
rect 5092 11830 5120 12174
rect 5080 11824 5132 11830
rect 5080 11766 5132 11772
rect 5552 11354 5580 13942
rect 6920 13932 6972 13938
rect 6920 13874 6972 13880
rect 5632 13728 5684 13734
rect 5632 13670 5684 13676
rect 5644 13326 5672 13670
rect 6423 13628 6731 13637
rect 6423 13626 6429 13628
rect 6485 13626 6509 13628
rect 6565 13626 6589 13628
rect 6645 13626 6669 13628
rect 6725 13626 6731 13628
rect 6485 13574 6487 13626
rect 6667 13574 6669 13626
rect 6423 13572 6429 13574
rect 6485 13572 6509 13574
rect 6565 13572 6589 13574
rect 6645 13572 6669 13574
rect 6725 13572 6731 13574
rect 6423 13563 6731 13572
rect 5632 13320 5684 13326
rect 5632 13262 5684 13268
rect 6423 12540 6731 12549
rect 6423 12538 6429 12540
rect 6485 12538 6509 12540
rect 6565 12538 6589 12540
rect 6645 12538 6669 12540
rect 6725 12538 6731 12540
rect 6485 12486 6487 12538
rect 6667 12486 6669 12538
rect 6423 12484 6429 12486
rect 6485 12484 6509 12486
rect 6565 12484 6589 12486
rect 6645 12484 6669 12486
rect 6725 12484 6731 12486
rect 6423 12475 6731 12484
rect 6000 12164 6052 12170
rect 6000 12106 6052 12112
rect 5632 11552 5684 11558
rect 5632 11494 5684 11500
rect 5540 11348 5592 11354
rect 5540 11290 5592 11296
rect 4620 10804 4672 10810
rect 4620 10746 4672 10752
rect 4620 10464 4672 10470
rect 4620 10406 4672 10412
rect 4632 10062 4660 10406
rect 4620 10056 4672 10062
rect 4620 9998 4672 10004
rect 4632 9722 4660 9998
rect 4620 9716 4672 9722
rect 4620 9658 4672 9664
rect 5552 9654 5580 11290
rect 5540 9648 5592 9654
rect 5540 9590 5592 9596
rect 5540 9512 5592 9518
rect 5540 9454 5592 9460
rect 4528 9444 4580 9450
rect 4528 9386 4580 9392
rect 5356 8968 5408 8974
rect 5356 8910 5408 8916
rect 5368 8090 5396 8910
rect 5356 8084 5408 8090
rect 5356 8026 5408 8032
rect 5552 7834 5580 9454
rect 5644 8974 5672 11494
rect 6012 11354 6040 12106
rect 6423 11452 6731 11461
rect 6423 11450 6429 11452
rect 6485 11450 6509 11452
rect 6565 11450 6589 11452
rect 6645 11450 6669 11452
rect 6725 11450 6731 11452
rect 6485 11398 6487 11450
rect 6667 11398 6669 11450
rect 6423 11396 6429 11398
rect 6485 11396 6509 11398
rect 6565 11396 6589 11398
rect 6645 11396 6669 11398
rect 6725 11396 6731 11398
rect 6423 11387 6731 11396
rect 6000 11348 6052 11354
rect 6000 11290 6052 11296
rect 6092 10736 6144 10742
rect 6092 10678 6144 10684
rect 5908 9920 5960 9926
rect 5908 9862 5960 9868
rect 5816 9512 5868 9518
rect 5816 9454 5868 9460
rect 5828 9042 5856 9454
rect 5816 9036 5868 9042
rect 5816 8978 5868 8984
rect 5632 8968 5684 8974
rect 5632 8910 5684 8916
rect 4436 7812 4488 7818
rect 5552 7806 5764 7834
rect 4436 7754 4488 7760
rect 5632 7744 5684 7750
rect 5632 7686 5684 7692
rect 5644 7546 5672 7686
rect 5736 7546 5764 7806
rect 5632 7540 5684 7546
rect 5632 7482 5684 7488
rect 5724 7540 5776 7546
rect 5724 7482 5776 7488
rect 5540 7404 5592 7410
rect 5540 7346 5592 7352
rect 5356 7336 5408 7342
rect 5356 7278 5408 7284
rect 5172 7200 5224 7206
rect 5172 7142 5224 7148
rect 3424 6860 3476 6866
rect 3424 6802 3476 6808
rect 3976 6860 4028 6866
rect 3976 6802 4028 6808
rect 3332 6316 3384 6322
rect 3332 6258 3384 6264
rect 3240 5908 3292 5914
rect 3240 5850 3292 5856
rect 3988 5778 4016 6802
rect 3976 5772 4028 5778
rect 3976 5714 4028 5720
rect 2136 5704 2188 5710
rect 2136 5646 2188 5652
rect 3988 5234 4016 5714
rect 5184 5710 5212 7142
rect 5264 6656 5316 6662
rect 5264 6598 5316 6604
rect 5276 5914 5304 6598
rect 5264 5908 5316 5914
rect 5264 5850 5316 5856
rect 5172 5704 5224 5710
rect 5172 5646 5224 5652
rect 3976 5228 4028 5234
rect 3976 5170 4028 5176
rect 4252 5228 4304 5234
rect 4252 5170 4304 5176
rect 940 5160 992 5166
rect 940 5102 992 5108
rect 952 4865 980 5102
rect 938 4856 994 4865
rect 4264 4826 4292 5170
rect 938 4791 994 4800
rect 4252 4820 4304 4826
rect 4252 4762 4304 4768
rect 5276 4622 5304 5850
rect 5368 5370 5396 7278
rect 5552 6662 5580 7346
rect 5828 7342 5856 8978
rect 5920 7954 5948 9862
rect 6104 9722 6132 10678
rect 6423 10364 6731 10373
rect 6423 10362 6429 10364
rect 6485 10362 6509 10364
rect 6565 10362 6589 10364
rect 6645 10362 6669 10364
rect 6725 10362 6731 10364
rect 6485 10310 6487 10362
rect 6667 10310 6669 10362
rect 6423 10308 6429 10310
rect 6485 10308 6509 10310
rect 6565 10308 6589 10310
rect 6645 10308 6669 10310
rect 6725 10308 6731 10310
rect 6423 10299 6731 10308
rect 6092 9716 6144 9722
rect 6092 9658 6144 9664
rect 6276 9580 6328 9586
rect 6276 9522 6328 9528
rect 6288 8090 6316 9522
rect 6932 9450 6960 13874
rect 8576 13456 8628 13462
rect 8576 13398 8628 13404
rect 7564 13388 7616 13394
rect 7564 13330 7616 13336
rect 7380 13184 7432 13190
rect 7380 13126 7432 13132
rect 7392 12442 7420 13126
rect 7380 12436 7432 12442
rect 7380 12378 7432 12384
rect 7576 12238 7604 13330
rect 8588 12850 8616 13398
rect 9876 12918 9904 14350
rect 11244 14272 11296 14278
rect 11244 14214 11296 14220
rect 11336 14272 11388 14278
rect 11336 14214 11388 14220
rect 11060 13388 11112 13394
rect 11060 13330 11112 13336
rect 10324 13184 10376 13190
rect 10324 13126 10376 13132
rect 9864 12912 9916 12918
rect 9864 12854 9916 12860
rect 8576 12844 8628 12850
rect 8576 12786 8628 12792
rect 7748 12640 7800 12646
rect 7748 12582 7800 12588
rect 7760 12238 7788 12582
rect 9680 12300 9732 12306
rect 9680 12242 9732 12248
rect 7564 12232 7616 12238
rect 7564 12174 7616 12180
rect 7748 12232 7800 12238
rect 7748 12174 7800 12180
rect 7380 12096 7432 12102
rect 7380 12038 7432 12044
rect 7392 11898 7420 12038
rect 7380 11892 7432 11898
rect 7380 11834 7432 11840
rect 7196 11552 7248 11558
rect 7196 11494 7248 11500
rect 7208 11218 7236 11494
rect 7576 11218 7604 12174
rect 7760 11898 7788 12174
rect 8208 12164 8260 12170
rect 8208 12106 8260 12112
rect 8220 11898 8248 12106
rect 7748 11892 7800 11898
rect 7748 11834 7800 11840
rect 8208 11892 8260 11898
rect 8208 11834 8260 11840
rect 9692 11694 9720 12242
rect 9680 11688 9732 11694
rect 9680 11630 9732 11636
rect 9876 11218 9904 12854
rect 10048 12844 10100 12850
rect 10048 12786 10100 12792
rect 10060 12442 10088 12786
rect 10048 12436 10100 12442
rect 10048 12378 10100 12384
rect 10336 12238 10364 13126
rect 11072 12442 11100 13330
rect 11256 13326 11284 14214
rect 11348 13870 11376 14214
rect 11896 14172 12204 14181
rect 11896 14170 11902 14172
rect 11958 14170 11982 14172
rect 12038 14170 12062 14172
rect 12118 14170 12142 14172
rect 12198 14170 12204 14172
rect 11958 14118 11960 14170
rect 12140 14118 12142 14170
rect 11896 14116 11902 14118
rect 11958 14116 11982 14118
rect 12038 14116 12062 14118
rect 12118 14116 12142 14118
rect 12198 14116 12204 14118
rect 11896 14107 12204 14116
rect 11336 13864 11388 13870
rect 11336 13806 11388 13812
rect 11428 13864 11480 13870
rect 11428 13806 11480 13812
rect 11440 13394 11468 13806
rect 12440 13728 12492 13734
rect 12440 13670 12492 13676
rect 11428 13388 11480 13394
rect 11428 13330 11480 13336
rect 11244 13320 11296 13326
rect 11244 13262 11296 13268
rect 11440 12918 11468 13330
rect 11796 13252 11848 13258
rect 11796 13194 11848 13200
rect 11704 13184 11756 13190
rect 11704 13126 11756 13132
rect 11716 12986 11744 13126
rect 11704 12980 11756 12986
rect 11704 12922 11756 12928
rect 11428 12912 11480 12918
rect 11428 12854 11480 12860
rect 11152 12844 11204 12850
rect 11152 12786 11204 12792
rect 11164 12646 11192 12786
rect 11152 12640 11204 12646
rect 11152 12582 11204 12588
rect 11060 12436 11112 12442
rect 11060 12378 11112 12384
rect 10324 12232 10376 12238
rect 10324 12174 10376 12180
rect 10784 11824 10836 11830
rect 10784 11766 10836 11772
rect 10324 11756 10376 11762
rect 10324 11698 10376 11704
rect 10232 11552 10284 11558
rect 10232 11494 10284 11500
rect 7196 11212 7248 11218
rect 7196 11154 7248 11160
rect 7564 11212 7616 11218
rect 7564 11154 7616 11160
rect 9864 11212 9916 11218
rect 9864 11154 9916 11160
rect 7932 11144 7984 11150
rect 7932 11086 7984 11092
rect 7944 10266 7972 11086
rect 8300 11076 8352 11082
rect 8300 11018 8352 11024
rect 8312 10810 8340 11018
rect 9588 11008 9640 11014
rect 9588 10950 9640 10956
rect 8300 10804 8352 10810
rect 8300 10746 8352 10752
rect 8392 10668 8444 10674
rect 8392 10610 8444 10616
rect 8404 10266 8432 10610
rect 7932 10260 7984 10266
rect 7932 10202 7984 10208
rect 8392 10260 8444 10266
rect 8392 10202 8444 10208
rect 7196 10056 7248 10062
rect 7196 9998 7248 10004
rect 7208 9586 7236 9998
rect 7944 9586 7972 10202
rect 8484 10192 8536 10198
rect 8484 10134 8536 10140
rect 7196 9580 7248 9586
rect 7196 9522 7248 9528
rect 7932 9580 7984 9586
rect 7932 9522 7984 9528
rect 6920 9444 6972 9450
rect 6920 9386 6972 9392
rect 8300 9376 8352 9382
rect 8300 9318 8352 9324
rect 6423 9276 6731 9285
rect 6423 9274 6429 9276
rect 6485 9274 6509 9276
rect 6565 9274 6589 9276
rect 6645 9274 6669 9276
rect 6725 9274 6731 9276
rect 6485 9222 6487 9274
rect 6667 9222 6669 9274
rect 6423 9220 6429 9222
rect 6485 9220 6509 9222
rect 6565 9220 6589 9222
rect 6645 9220 6669 9222
rect 6725 9220 6731 9222
rect 6423 9211 6731 9220
rect 8208 8968 8260 8974
rect 8208 8910 8260 8916
rect 6828 8832 6880 8838
rect 6828 8774 6880 8780
rect 6423 8188 6731 8197
rect 6423 8186 6429 8188
rect 6485 8186 6509 8188
rect 6565 8186 6589 8188
rect 6645 8186 6669 8188
rect 6725 8186 6731 8188
rect 6485 8134 6487 8186
rect 6667 8134 6669 8186
rect 6423 8132 6429 8134
rect 6485 8132 6509 8134
rect 6565 8132 6589 8134
rect 6645 8132 6669 8134
rect 6725 8132 6731 8134
rect 6423 8123 6731 8132
rect 6276 8084 6328 8090
rect 6276 8026 6328 8032
rect 5908 7948 5960 7954
rect 5908 7890 5960 7896
rect 6840 7478 6868 8774
rect 8220 8634 8248 8910
rect 8208 8628 8260 8634
rect 8208 8570 8260 8576
rect 8312 8430 8340 9318
rect 8496 9042 8524 10134
rect 9600 10130 9628 10950
rect 9876 10742 9904 11154
rect 10244 11150 10272 11494
rect 10232 11144 10284 11150
rect 10232 11086 10284 11092
rect 9864 10736 9916 10742
rect 9864 10678 9916 10684
rect 9588 10124 9640 10130
rect 9588 10066 9640 10072
rect 8576 10056 8628 10062
rect 8576 9998 8628 10004
rect 8484 9036 8536 9042
rect 8484 8978 8536 8984
rect 8300 8424 8352 8430
rect 8300 8366 8352 8372
rect 6920 8356 6972 8362
rect 6920 8298 6972 8304
rect 6828 7472 6880 7478
rect 6828 7414 6880 7420
rect 5816 7336 5868 7342
rect 5816 7278 5868 7284
rect 6423 7100 6731 7109
rect 6423 7098 6429 7100
rect 6485 7098 6509 7100
rect 6565 7098 6589 7100
rect 6645 7098 6669 7100
rect 6725 7098 6731 7100
rect 6485 7046 6487 7098
rect 6667 7046 6669 7098
rect 6423 7044 6429 7046
rect 6485 7044 6509 7046
rect 6565 7044 6589 7046
rect 6645 7044 6669 7046
rect 6725 7044 6731 7046
rect 6423 7035 6731 7044
rect 5540 6656 5592 6662
rect 5540 6598 5592 6604
rect 6000 6656 6052 6662
rect 6000 6598 6052 6604
rect 5816 5772 5868 5778
rect 5816 5714 5868 5720
rect 5356 5364 5408 5370
rect 5356 5306 5408 5312
rect 5828 4690 5856 5714
rect 6012 5710 6040 6598
rect 6932 6390 6960 8298
rect 8024 7880 8076 7886
rect 8024 7822 8076 7828
rect 7932 7812 7984 7818
rect 7932 7754 7984 7760
rect 7944 7478 7972 7754
rect 7932 7472 7984 7478
rect 7932 7414 7984 7420
rect 8036 7342 8064 7822
rect 8312 7818 8340 8366
rect 8588 8090 8616 9998
rect 9312 9920 9364 9926
rect 9312 9862 9364 9868
rect 9128 9648 9180 9654
rect 9128 9590 9180 9596
rect 8944 8832 8996 8838
rect 8944 8774 8996 8780
rect 8956 8566 8984 8774
rect 8944 8560 8996 8566
rect 8944 8502 8996 8508
rect 8668 8424 8720 8430
rect 8668 8366 8720 8372
rect 8576 8084 8628 8090
rect 8576 8026 8628 8032
rect 8576 7880 8628 7886
rect 8576 7822 8628 7828
rect 8300 7812 8352 7818
rect 8300 7754 8352 7760
rect 8024 7336 8076 7342
rect 8024 7278 8076 7284
rect 8588 7002 8616 7822
rect 8576 6996 8628 7002
rect 8576 6938 8628 6944
rect 8680 6798 8708 8366
rect 9140 7954 9168 9590
rect 9324 8974 9352 9862
rect 9876 9602 9904 10678
rect 10336 10538 10364 11698
rect 10796 10810 10824 11766
rect 10876 11688 10928 11694
rect 10876 11630 10928 11636
rect 10888 11082 10916 11630
rect 10876 11076 10928 11082
rect 10876 11018 10928 11024
rect 10784 10804 10836 10810
rect 10784 10746 10836 10752
rect 10888 10606 10916 11018
rect 10968 10668 11020 10674
rect 10968 10610 11020 10616
rect 10876 10600 10928 10606
rect 10876 10542 10928 10548
rect 10324 10532 10376 10538
rect 10324 10474 10376 10480
rect 10600 10192 10652 10198
rect 10600 10134 10652 10140
rect 10416 9988 10468 9994
rect 10416 9930 10468 9936
rect 10048 9920 10100 9926
rect 10048 9862 10100 9868
rect 9784 9586 9904 9602
rect 9772 9580 9904 9586
rect 9824 9574 9904 9580
rect 9772 9522 9824 9528
rect 9784 9042 9812 9522
rect 9772 9036 9824 9042
rect 9772 8978 9824 8984
rect 9312 8968 9364 8974
rect 9312 8910 9364 8916
rect 10060 8634 10088 9862
rect 10324 9376 10376 9382
rect 10324 9318 10376 9324
rect 10336 8974 10364 9318
rect 10324 8968 10376 8974
rect 10324 8910 10376 8916
rect 9680 8628 9732 8634
rect 9680 8570 9732 8576
rect 10048 8628 10100 8634
rect 10048 8570 10100 8576
rect 9496 8492 9548 8498
rect 9496 8434 9548 8440
rect 9128 7948 9180 7954
rect 9128 7890 9180 7896
rect 9140 7546 9168 7890
rect 9508 7546 9536 8434
rect 9128 7540 9180 7546
rect 9128 7482 9180 7488
rect 9496 7540 9548 7546
rect 9496 7482 9548 7488
rect 9140 6798 9168 7482
rect 9312 7404 9364 7410
rect 9312 7346 9364 7352
rect 7932 6792 7984 6798
rect 7932 6734 7984 6740
rect 8668 6792 8720 6798
rect 8668 6734 8720 6740
rect 9128 6792 9180 6798
rect 9128 6734 9180 6740
rect 6920 6384 6972 6390
rect 6920 6326 6972 6332
rect 7944 6322 7972 6734
rect 8680 6322 8708 6734
rect 9324 6458 9352 7346
rect 9692 6662 9720 8570
rect 9772 7812 9824 7818
rect 9772 7754 9824 7760
rect 9784 7342 9812 7754
rect 9772 7336 9824 7342
rect 9772 7278 9824 7284
rect 9784 6798 9812 7278
rect 9772 6792 9824 6798
rect 9772 6734 9824 6740
rect 9404 6656 9456 6662
rect 9404 6598 9456 6604
rect 9680 6656 9732 6662
rect 9680 6598 9732 6604
rect 9312 6452 9364 6458
rect 9312 6394 9364 6400
rect 7932 6316 7984 6322
rect 7932 6258 7984 6264
rect 8668 6316 8720 6322
rect 8668 6258 8720 6264
rect 6423 6012 6731 6021
rect 6423 6010 6429 6012
rect 6485 6010 6509 6012
rect 6565 6010 6589 6012
rect 6645 6010 6669 6012
rect 6725 6010 6731 6012
rect 6485 5958 6487 6010
rect 6667 5958 6669 6010
rect 6423 5956 6429 5958
rect 6485 5956 6509 5958
rect 6565 5956 6589 5958
rect 6645 5956 6669 5958
rect 6725 5956 6731 5958
rect 6423 5947 6731 5956
rect 6000 5704 6052 5710
rect 6000 5646 6052 5652
rect 7748 5568 7800 5574
rect 7748 5510 7800 5516
rect 6423 4924 6731 4933
rect 6423 4922 6429 4924
rect 6485 4922 6509 4924
rect 6565 4922 6589 4924
rect 6645 4922 6669 4924
rect 6725 4922 6731 4924
rect 6485 4870 6487 4922
rect 6667 4870 6669 4922
rect 6423 4868 6429 4870
rect 6485 4868 6509 4870
rect 6565 4868 6589 4870
rect 6645 4868 6669 4870
rect 6725 4868 6731 4870
rect 6423 4859 6731 4868
rect 5816 4684 5868 4690
rect 5816 4626 5868 4632
rect 5264 4616 5316 4622
rect 5264 4558 5316 4564
rect 5908 4480 5960 4486
rect 5908 4422 5960 4428
rect 5920 3534 5948 4422
rect 6423 3836 6731 3845
rect 6423 3834 6429 3836
rect 6485 3834 6509 3836
rect 6565 3834 6589 3836
rect 6645 3834 6669 3836
rect 6725 3834 6731 3836
rect 6485 3782 6487 3834
rect 6667 3782 6669 3834
rect 6423 3780 6429 3782
rect 6485 3780 6509 3782
rect 6565 3780 6589 3782
rect 6645 3780 6669 3782
rect 6725 3780 6731 3782
rect 6423 3771 6731 3780
rect 940 3528 992 3534
rect 938 3496 940 3505
rect 5908 3528 5960 3534
rect 992 3496 994 3505
rect 5908 3470 5960 3476
rect 938 3431 994 3440
rect 5724 3392 5776 3398
rect 5724 3334 5776 3340
rect 940 2848 992 2854
rect 940 2790 992 2796
rect 20 2508 72 2514
rect 20 2450 72 2456
rect 32 800 60 2450
rect 952 1465 980 2790
rect 5736 2446 5764 3334
rect 7760 3058 7788 5510
rect 9324 5234 9352 6394
rect 9312 5228 9364 5234
rect 9312 5170 9364 5176
rect 9416 3058 9444 6598
rect 9588 6316 9640 6322
rect 9588 6258 9640 6264
rect 9600 5914 9628 6258
rect 9588 5908 9640 5914
rect 9588 5850 9640 5856
rect 10060 5710 10088 8570
rect 10428 5710 10456 9930
rect 10508 7880 10560 7886
rect 10508 7822 10560 7828
rect 10520 7750 10548 7822
rect 10508 7744 10560 7750
rect 10508 7686 10560 7692
rect 10520 6390 10548 7686
rect 10612 7342 10640 10134
rect 10692 9512 10744 9518
rect 10692 9454 10744 9460
rect 10704 9178 10732 9454
rect 10980 9450 11008 10610
rect 11072 10538 11100 12378
rect 11164 12102 11192 12582
rect 11440 12238 11468 12854
rect 11808 12442 11836 13194
rect 11896 13084 12204 13093
rect 11896 13082 11902 13084
rect 11958 13082 11982 13084
rect 12038 13082 12062 13084
rect 12118 13082 12142 13084
rect 12198 13082 12204 13084
rect 11958 13030 11960 13082
rect 12140 13030 12142 13082
rect 11896 13028 11902 13030
rect 11958 13028 11982 13030
rect 12038 13028 12062 13030
rect 12118 13028 12142 13030
rect 12198 13028 12204 13030
rect 11896 13019 12204 13028
rect 12348 12776 12400 12782
rect 12348 12718 12400 12724
rect 11796 12436 11848 12442
rect 11796 12378 11848 12384
rect 12360 12374 12388 12718
rect 12348 12368 12400 12374
rect 12348 12310 12400 12316
rect 11428 12232 11480 12238
rect 11428 12174 11480 12180
rect 11152 12096 11204 12102
rect 11152 12038 11204 12044
rect 11440 11218 11468 12174
rect 11896 11996 12204 12005
rect 11896 11994 11902 11996
rect 11958 11994 11982 11996
rect 12038 11994 12062 11996
rect 12118 11994 12142 11996
rect 12198 11994 12204 11996
rect 11958 11942 11960 11994
rect 12140 11942 12142 11994
rect 11896 11940 11902 11942
rect 11958 11940 11982 11942
rect 12038 11940 12062 11942
rect 12118 11940 12142 11942
rect 12198 11940 12204 11942
rect 11896 11931 12204 11940
rect 11428 11212 11480 11218
rect 11428 11154 11480 11160
rect 11336 11008 11388 11014
rect 11336 10950 11388 10956
rect 11348 10742 11376 10950
rect 11336 10736 11388 10742
rect 11336 10678 11388 10684
rect 11440 10674 11468 11154
rect 12360 11082 12388 12310
rect 12452 12170 12480 13670
rect 12808 13184 12860 13190
rect 12808 13126 12860 13132
rect 12440 12164 12492 12170
rect 12440 12106 12492 12112
rect 12348 11076 12400 11082
rect 12348 11018 12400 11024
rect 11896 10908 12204 10917
rect 11896 10906 11902 10908
rect 11958 10906 11982 10908
rect 12038 10906 12062 10908
rect 12118 10906 12142 10908
rect 12198 10906 12204 10908
rect 11958 10854 11960 10906
rect 12140 10854 12142 10906
rect 11896 10852 11902 10854
rect 11958 10852 11982 10854
rect 12038 10852 12062 10854
rect 12118 10852 12142 10854
rect 12198 10852 12204 10854
rect 11896 10843 12204 10852
rect 11428 10668 11480 10674
rect 11428 10610 11480 10616
rect 11060 10532 11112 10538
rect 11060 10474 11112 10480
rect 11440 10266 11468 10610
rect 11428 10260 11480 10266
rect 11428 10202 11480 10208
rect 12820 10033 12848 13126
rect 12900 11756 12952 11762
rect 12900 11698 12952 11704
rect 12912 11082 12940 11698
rect 12900 11076 12952 11082
rect 12900 11018 12952 11024
rect 12806 10024 12862 10033
rect 12806 9959 12862 9968
rect 11896 9820 12204 9829
rect 11896 9818 11902 9820
rect 11958 9818 11982 9820
rect 12038 9818 12062 9820
rect 12118 9818 12142 9820
rect 12198 9818 12204 9820
rect 11958 9766 11960 9818
rect 12140 9766 12142 9818
rect 11896 9764 11902 9766
rect 11958 9764 11982 9766
rect 12038 9764 12062 9766
rect 12118 9764 12142 9766
rect 12198 9764 12204 9766
rect 11896 9755 12204 9764
rect 12912 9586 12940 11018
rect 13096 9602 13124 17002
rect 14188 16584 14240 16590
rect 14188 16526 14240 16532
rect 13360 14340 13412 14346
rect 13360 14282 13412 14288
rect 13372 13938 13400 14282
rect 13360 13932 13412 13938
rect 13360 13874 13412 13880
rect 13820 12844 13872 12850
rect 13820 12786 13872 12792
rect 13176 12776 13228 12782
rect 13176 12718 13228 12724
rect 13188 11762 13216 12718
rect 13832 12442 13860 12786
rect 14096 12640 14148 12646
rect 14096 12582 14148 12588
rect 13820 12436 13872 12442
rect 13820 12378 13872 12384
rect 13360 12096 13412 12102
rect 13360 12038 13412 12044
rect 13372 11898 13400 12038
rect 13360 11892 13412 11898
rect 13360 11834 13412 11840
rect 13176 11756 13228 11762
rect 13176 11698 13228 11704
rect 13912 10668 13964 10674
rect 13912 10610 13964 10616
rect 14004 10668 14056 10674
rect 14004 10610 14056 10616
rect 13636 10124 13688 10130
rect 13636 10066 13688 10072
rect 13096 9586 13216 9602
rect 11612 9580 11664 9586
rect 11612 9522 11664 9528
rect 12900 9580 12952 9586
rect 13096 9580 13228 9586
rect 13096 9574 13176 9580
rect 12900 9522 12952 9528
rect 13176 9522 13228 9528
rect 10968 9444 11020 9450
rect 10968 9386 11020 9392
rect 11624 9178 11652 9522
rect 10692 9172 10744 9178
rect 10692 9114 10744 9120
rect 11612 9172 11664 9178
rect 11612 9114 11664 9120
rect 13188 8974 13216 9522
rect 13648 9110 13676 10066
rect 13820 9920 13872 9926
rect 13820 9862 13872 9868
rect 13832 9722 13860 9862
rect 13820 9716 13872 9722
rect 13820 9658 13872 9664
rect 13924 9178 13952 10610
rect 14016 10198 14044 10610
rect 14108 10606 14136 12582
rect 14096 10600 14148 10606
rect 14096 10542 14148 10548
rect 14004 10192 14056 10198
rect 14004 10134 14056 10140
rect 13912 9172 13964 9178
rect 13912 9114 13964 9120
rect 13636 9104 13688 9110
rect 13636 9046 13688 9052
rect 11796 8968 11848 8974
rect 11796 8910 11848 8916
rect 13176 8968 13228 8974
rect 13176 8910 13228 8916
rect 11808 8090 11836 8910
rect 11896 8732 12204 8741
rect 11896 8730 11902 8732
rect 11958 8730 11982 8732
rect 12038 8730 12062 8732
rect 12118 8730 12142 8732
rect 12198 8730 12204 8732
rect 11958 8678 11960 8730
rect 12140 8678 12142 8730
rect 11896 8676 11902 8678
rect 11958 8676 11982 8678
rect 12038 8676 12062 8678
rect 12118 8676 12142 8678
rect 12198 8676 12204 8678
rect 11896 8667 12204 8676
rect 11796 8084 11848 8090
rect 11796 8026 11848 8032
rect 14108 7954 14136 10542
rect 14200 10538 14228 16526
rect 16316 14521 16344 17002
rect 16302 14512 16358 14521
rect 16302 14447 16358 14456
rect 14372 14272 14424 14278
rect 14372 14214 14424 14220
rect 14384 13326 14412 14214
rect 16316 14074 16344 14447
rect 16304 14068 16356 14074
rect 16304 14010 16356 14016
rect 14648 14000 14700 14006
rect 14648 13942 14700 13948
rect 14464 13728 14516 13734
rect 14464 13670 14516 13676
rect 14476 13326 14504 13670
rect 14660 13530 14688 13942
rect 14648 13524 14700 13530
rect 14648 13466 14700 13472
rect 14372 13320 14424 13326
rect 14372 13262 14424 13268
rect 14464 13320 14516 13326
rect 14464 13262 14516 13268
rect 14384 12646 14412 13262
rect 14556 12980 14608 12986
rect 14556 12922 14608 12928
rect 14372 12640 14424 12646
rect 14372 12582 14424 12588
rect 14568 12238 14596 12922
rect 14556 12232 14608 12238
rect 14556 12174 14608 12180
rect 14648 11756 14700 11762
rect 14648 11698 14700 11704
rect 16396 11756 16448 11762
rect 16396 11698 16448 11704
rect 14660 11354 14688 11698
rect 14648 11348 14700 11354
rect 14648 11290 14700 11296
rect 14372 11144 14424 11150
rect 14372 11086 14424 11092
rect 14188 10532 14240 10538
rect 14188 10474 14240 10480
rect 14280 10056 14332 10062
rect 14280 9998 14332 10004
rect 14292 9722 14320 9998
rect 14384 9926 14412 11086
rect 15844 11076 15896 11082
rect 15844 11018 15896 11024
rect 15856 10810 15884 11018
rect 15844 10804 15896 10810
rect 15844 10746 15896 10752
rect 16304 10668 16356 10674
rect 16304 10610 16356 10616
rect 15200 10464 15252 10470
rect 15200 10406 15252 10412
rect 14648 10056 14700 10062
rect 14648 9998 14700 10004
rect 14660 9926 14688 9998
rect 14372 9920 14424 9926
rect 14372 9862 14424 9868
rect 14648 9920 14700 9926
rect 14648 9862 14700 9868
rect 14280 9716 14332 9722
rect 14280 9658 14332 9664
rect 14660 8922 14688 9862
rect 15212 9654 15240 10406
rect 16316 10198 16344 10610
rect 16304 10192 16356 10198
rect 16304 10134 16356 10140
rect 15660 9988 15712 9994
rect 15660 9930 15712 9936
rect 15200 9648 15252 9654
rect 15200 9590 15252 9596
rect 15476 9036 15528 9042
rect 15476 8978 15528 8984
rect 14660 8894 14872 8922
rect 14740 8832 14792 8838
rect 14740 8774 14792 8780
rect 14372 8492 14424 8498
rect 14372 8434 14424 8440
rect 14096 7948 14148 7954
rect 14096 7890 14148 7896
rect 13360 7880 13412 7886
rect 13360 7822 13412 7828
rect 11152 7812 11204 7818
rect 11152 7754 11204 7760
rect 10600 7336 10652 7342
rect 10600 7278 10652 7284
rect 11164 6458 11192 7754
rect 11612 7744 11664 7750
rect 11612 7686 11664 7692
rect 12992 7744 13044 7750
rect 12992 7686 13044 7692
rect 11624 7546 11652 7686
rect 11896 7644 12204 7653
rect 11896 7642 11902 7644
rect 11958 7642 11982 7644
rect 12038 7642 12062 7644
rect 12118 7642 12142 7644
rect 12198 7642 12204 7644
rect 11958 7590 11960 7642
rect 12140 7590 12142 7642
rect 11896 7588 11902 7590
rect 11958 7588 11982 7590
rect 12038 7588 12062 7590
rect 12118 7588 12142 7590
rect 12198 7588 12204 7590
rect 11896 7579 12204 7588
rect 11612 7540 11664 7546
rect 11612 7482 11664 7488
rect 12624 7404 12676 7410
rect 12624 7346 12676 7352
rect 12256 7336 12308 7342
rect 12256 7278 12308 7284
rect 11612 6860 11664 6866
rect 11612 6802 11664 6808
rect 11152 6452 11204 6458
rect 11152 6394 11204 6400
rect 10508 6384 10560 6390
rect 10508 6326 10560 6332
rect 9588 5704 9640 5710
rect 9588 5646 9640 5652
rect 10048 5704 10100 5710
rect 10048 5646 10100 5652
rect 10416 5704 10468 5710
rect 10416 5646 10468 5652
rect 9600 5302 9628 5646
rect 9956 5568 10008 5574
rect 9956 5510 10008 5516
rect 9588 5296 9640 5302
rect 9588 5238 9640 5244
rect 9968 3738 9996 5510
rect 11624 4554 11652 6802
rect 12268 6798 12296 7278
rect 12440 7200 12492 7206
rect 12440 7142 12492 7148
rect 12452 6798 12480 7142
rect 12532 6996 12584 7002
rect 12532 6938 12584 6944
rect 11796 6792 11848 6798
rect 11716 6752 11796 6780
rect 11716 6186 11744 6752
rect 11796 6734 11848 6740
rect 12256 6792 12308 6798
rect 12256 6734 12308 6740
rect 12440 6792 12492 6798
rect 12440 6734 12492 6740
rect 11896 6556 12204 6565
rect 11896 6554 11902 6556
rect 11958 6554 11982 6556
rect 12038 6554 12062 6556
rect 12118 6554 12142 6556
rect 12198 6554 12204 6556
rect 11958 6502 11960 6554
rect 12140 6502 12142 6554
rect 11896 6500 11902 6502
rect 11958 6500 11982 6502
rect 12038 6500 12062 6502
rect 12118 6500 12142 6502
rect 12198 6500 12204 6502
rect 11896 6491 12204 6500
rect 12070 6352 12126 6361
rect 12070 6287 12072 6296
rect 12124 6287 12126 6296
rect 12072 6258 12124 6264
rect 11704 6180 11756 6186
rect 11704 6122 11756 6128
rect 12268 5914 12296 6734
rect 12544 6458 12572 6938
rect 12636 6458 12664 7346
rect 12808 6656 12860 6662
rect 12808 6598 12860 6604
rect 12532 6452 12584 6458
rect 12532 6394 12584 6400
rect 12624 6452 12676 6458
rect 12624 6394 12676 6400
rect 12532 6180 12584 6186
rect 12532 6122 12584 6128
rect 12256 5908 12308 5914
rect 12256 5850 12308 5856
rect 11896 5468 12204 5477
rect 11896 5466 11902 5468
rect 11958 5466 11982 5468
rect 12038 5466 12062 5468
rect 12118 5466 12142 5468
rect 12198 5466 12204 5468
rect 11958 5414 11960 5466
rect 12140 5414 12142 5466
rect 11896 5412 11902 5414
rect 11958 5412 11982 5414
rect 12038 5412 12062 5414
rect 12118 5412 12142 5414
rect 12198 5412 12204 5414
rect 11896 5403 12204 5412
rect 12268 5234 12296 5850
rect 12544 5846 12572 6122
rect 12532 5840 12584 5846
rect 12532 5782 12584 5788
rect 12256 5228 12308 5234
rect 12256 5170 12308 5176
rect 12268 4554 12296 5170
rect 11612 4548 11664 4554
rect 11612 4490 11664 4496
rect 12256 4548 12308 4554
rect 12256 4490 12308 4496
rect 11896 4380 12204 4389
rect 11896 4378 11902 4380
rect 11958 4378 11982 4380
rect 12038 4378 12062 4380
rect 12118 4378 12142 4380
rect 12198 4378 12204 4380
rect 11958 4326 11960 4378
rect 12140 4326 12142 4378
rect 11896 4324 11902 4326
rect 11958 4324 11982 4326
rect 12038 4324 12062 4326
rect 12118 4324 12142 4326
rect 12198 4324 12204 4326
rect 11896 4315 12204 4324
rect 9956 3732 10008 3738
rect 9956 3674 10008 3680
rect 11896 3292 12204 3301
rect 11896 3290 11902 3292
rect 11958 3290 11982 3292
rect 12038 3290 12062 3292
rect 12118 3290 12142 3292
rect 12198 3290 12204 3292
rect 11958 3238 11960 3290
rect 12140 3238 12142 3290
rect 11896 3236 11902 3238
rect 11958 3236 11982 3238
rect 12038 3236 12062 3238
rect 12118 3236 12142 3238
rect 12198 3236 12204 3238
rect 11896 3227 12204 3236
rect 7748 3052 7800 3058
rect 7748 2994 7800 3000
rect 9404 3052 9456 3058
rect 9404 2994 9456 3000
rect 9588 2848 9640 2854
rect 9588 2790 9640 2796
rect 6423 2748 6731 2757
rect 6423 2746 6429 2748
rect 6485 2746 6509 2748
rect 6565 2746 6589 2748
rect 6645 2746 6669 2748
rect 6725 2746 6731 2748
rect 6485 2694 6487 2746
rect 6667 2694 6669 2746
rect 6423 2692 6429 2694
rect 6485 2692 6509 2694
rect 6565 2692 6589 2694
rect 6645 2692 6669 2694
rect 6725 2692 6731 2694
rect 6423 2683 6731 2692
rect 9600 2446 9628 2790
rect 12820 2514 12848 6598
rect 13004 6186 13032 7686
rect 13176 6384 13228 6390
rect 13372 6372 13400 7822
rect 13728 7812 13780 7818
rect 13728 7754 13780 7760
rect 13740 7002 13768 7754
rect 14384 7750 14412 8434
rect 14648 8288 14700 8294
rect 14648 8230 14700 8236
rect 14464 7880 14516 7886
rect 14464 7822 14516 7828
rect 14372 7744 14424 7750
rect 14372 7686 14424 7692
rect 14476 7546 14504 7822
rect 14464 7540 14516 7546
rect 14464 7482 14516 7488
rect 14660 7002 14688 8230
rect 14752 7206 14780 8774
rect 14844 7993 14872 8894
rect 14924 8424 14976 8430
rect 14924 8366 14976 8372
rect 14936 8090 14964 8366
rect 14924 8084 14976 8090
rect 14924 8026 14976 8032
rect 14830 7984 14886 7993
rect 14830 7919 14886 7928
rect 14740 7200 14792 7206
rect 14740 7142 14792 7148
rect 14844 7018 14872 7919
rect 14936 7410 14964 8026
rect 15292 7880 15344 7886
rect 15292 7822 15344 7828
rect 15016 7812 15068 7818
rect 15016 7754 15068 7760
rect 14924 7404 14976 7410
rect 14924 7346 14976 7352
rect 15028 7206 15056 7754
rect 15108 7744 15160 7750
rect 15108 7686 15160 7692
rect 15200 7744 15252 7750
rect 15200 7686 15252 7692
rect 15120 7410 15148 7686
rect 15212 7478 15240 7686
rect 15200 7472 15252 7478
rect 15200 7414 15252 7420
rect 15108 7404 15160 7410
rect 15108 7346 15160 7352
rect 14924 7200 14976 7206
rect 14924 7142 14976 7148
rect 15016 7200 15068 7206
rect 15016 7142 15068 7148
rect 13728 6996 13780 7002
rect 13728 6938 13780 6944
rect 14648 6996 14700 7002
rect 14648 6938 14700 6944
rect 14752 6990 14872 7018
rect 13636 6656 13688 6662
rect 13636 6598 13688 6604
rect 13740 6610 13768 6938
rect 14280 6792 14332 6798
rect 14280 6734 14332 6740
rect 13452 6384 13504 6390
rect 13228 6344 13452 6372
rect 13176 6326 13228 6332
rect 13452 6326 13504 6332
rect 13360 6248 13412 6254
rect 13648 6225 13676 6598
rect 13740 6582 13952 6610
rect 13728 6452 13780 6458
rect 13728 6394 13780 6400
rect 13360 6190 13412 6196
rect 13634 6216 13690 6225
rect 12992 6180 13044 6186
rect 12992 6122 13044 6128
rect 13004 5914 13032 6122
rect 13176 6112 13228 6118
rect 13176 6054 13228 6060
rect 12992 5908 13044 5914
rect 12992 5850 13044 5856
rect 13188 5710 13216 6054
rect 13372 5778 13400 6190
rect 13634 6151 13690 6160
rect 13740 5914 13768 6394
rect 13924 6338 13952 6582
rect 14292 6390 14320 6734
rect 14464 6724 14516 6730
rect 14464 6666 14516 6672
rect 14280 6384 14332 6390
rect 13924 6322 14136 6338
rect 14280 6326 14332 6332
rect 13924 6316 14148 6322
rect 13924 6310 14096 6316
rect 14096 6258 14148 6264
rect 14096 6112 14148 6118
rect 14096 6054 14148 6060
rect 13728 5908 13780 5914
rect 13728 5850 13780 5856
rect 13360 5772 13412 5778
rect 13360 5714 13412 5720
rect 13176 5704 13228 5710
rect 13176 5646 13228 5652
rect 13084 5228 13136 5234
rect 13084 5170 13136 5176
rect 13096 4282 13124 5170
rect 13188 4826 13216 5646
rect 14108 5370 14136 6054
rect 14476 5914 14504 6666
rect 14648 6656 14700 6662
rect 14648 6598 14700 6604
rect 14660 6186 14688 6598
rect 14648 6180 14700 6186
rect 14648 6122 14700 6128
rect 14464 5908 14516 5914
rect 14464 5850 14516 5856
rect 14188 5840 14240 5846
rect 14188 5782 14240 5788
rect 14096 5364 14148 5370
rect 14096 5306 14148 5312
rect 14108 5234 14136 5306
rect 14096 5228 14148 5234
rect 14096 5170 14148 5176
rect 14200 5166 14228 5782
rect 14660 5778 14688 6122
rect 14648 5772 14700 5778
rect 14648 5714 14700 5720
rect 14660 5166 14688 5714
rect 14752 5234 14780 6990
rect 14832 6860 14884 6866
rect 14832 6802 14884 6808
rect 14844 6390 14872 6802
rect 14936 6798 14964 7142
rect 14924 6792 14976 6798
rect 14924 6734 14976 6740
rect 15120 6730 15148 7346
rect 15108 6724 15160 6730
rect 15108 6666 15160 6672
rect 15304 6662 15332 7822
rect 15292 6656 15344 6662
rect 15292 6598 15344 6604
rect 14832 6384 14884 6390
rect 14832 6326 14884 6332
rect 14924 6384 14976 6390
rect 14924 6326 14976 6332
rect 14844 5710 14872 6326
rect 14936 6118 14964 6326
rect 14924 6112 14976 6118
rect 14924 6054 14976 6060
rect 15292 6112 15344 6118
rect 15292 6054 15344 6060
rect 15304 5914 15332 6054
rect 15292 5908 15344 5914
rect 15292 5850 15344 5856
rect 14832 5704 14884 5710
rect 14832 5646 14884 5652
rect 14740 5228 14792 5234
rect 14740 5170 14792 5176
rect 14188 5160 14240 5166
rect 14188 5102 14240 5108
rect 14648 5160 14700 5166
rect 14648 5102 14700 5108
rect 13544 5024 13596 5030
rect 13544 4966 13596 4972
rect 14280 5024 14332 5030
rect 14280 4966 14332 4972
rect 15200 5024 15252 5030
rect 15200 4966 15252 4972
rect 13176 4820 13228 4826
rect 13176 4762 13228 4768
rect 13556 4282 13584 4966
rect 13084 4276 13136 4282
rect 13084 4218 13136 4224
rect 13544 4276 13596 4282
rect 13544 4218 13596 4224
rect 14292 4078 14320 4966
rect 15212 4622 15240 4966
rect 15200 4616 15252 4622
rect 15200 4558 15252 4564
rect 14832 4480 14884 4486
rect 14832 4422 14884 4428
rect 14844 4214 14872 4422
rect 14832 4208 14884 4214
rect 14832 4150 14884 4156
rect 15304 4078 15332 5850
rect 15488 5370 15516 8978
rect 15672 8634 15700 9930
rect 16408 9450 16436 11698
rect 16592 10810 16620 17138
rect 17370 16892 17678 16901
rect 17370 16890 17376 16892
rect 17432 16890 17456 16892
rect 17512 16890 17536 16892
rect 17592 16890 17616 16892
rect 17672 16890 17678 16892
rect 17432 16838 17434 16890
rect 17614 16838 17616 16890
rect 17370 16836 17376 16838
rect 17432 16836 17456 16838
rect 17512 16836 17536 16838
rect 17592 16836 17616 16838
rect 17672 16836 17678 16838
rect 17370 16827 17678 16836
rect 20732 16454 20760 17138
rect 23296 16992 23348 16998
rect 23296 16934 23348 16940
rect 30932 16992 30984 16998
rect 30932 16934 30984 16940
rect 32220 16992 32272 16998
rect 32220 16934 32272 16940
rect 34888 16992 34940 16998
rect 34888 16934 34940 16940
rect 38936 16992 38988 16998
rect 38936 16934 38988 16940
rect 20720 16448 20772 16454
rect 20720 16390 20772 16396
rect 22843 16348 23151 16357
rect 22843 16346 22849 16348
rect 22905 16346 22929 16348
rect 22985 16346 23009 16348
rect 23065 16346 23089 16348
rect 23145 16346 23151 16348
rect 22905 16294 22907 16346
rect 23087 16294 23089 16346
rect 22843 16292 22849 16294
rect 22905 16292 22929 16294
rect 22985 16292 23009 16294
rect 23065 16292 23089 16294
rect 23145 16292 23151 16294
rect 22843 16283 23151 16292
rect 17370 15804 17678 15813
rect 17370 15802 17376 15804
rect 17432 15802 17456 15804
rect 17512 15802 17536 15804
rect 17592 15802 17616 15804
rect 17672 15802 17678 15804
rect 17432 15750 17434 15802
rect 17614 15750 17616 15802
rect 17370 15748 17376 15750
rect 17432 15748 17456 15750
rect 17512 15748 17536 15750
rect 17592 15748 17616 15750
rect 17672 15748 17678 15750
rect 17370 15739 17678 15748
rect 22843 15260 23151 15269
rect 22843 15258 22849 15260
rect 22905 15258 22929 15260
rect 22985 15258 23009 15260
rect 23065 15258 23089 15260
rect 23145 15258 23151 15260
rect 22905 15206 22907 15258
rect 23087 15206 23089 15258
rect 22843 15204 22849 15206
rect 22905 15204 22929 15206
rect 22985 15204 23009 15206
rect 23065 15204 23089 15206
rect 23145 15204 23151 15206
rect 22843 15195 23151 15204
rect 23308 15162 23336 16934
rect 28317 16892 28625 16901
rect 28317 16890 28323 16892
rect 28379 16890 28403 16892
rect 28459 16890 28483 16892
rect 28539 16890 28563 16892
rect 28619 16890 28625 16892
rect 28379 16838 28381 16890
rect 28561 16838 28563 16890
rect 28317 16836 28323 16838
rect 28379 16836 28403 16838
rect 28459 16836 28483 16838
rect 28539 16836 28563 16838
rect 28619 16836 28625 16838
rect 28317 16827 28625 16836
rect 27620 16584 27672 16590
rect 27620 16526 27672 16532
rect 23296 15156 23348 15162
rect 23296 15098 23348 15104
rect 18880 15088 18932 15094
rect 18880 15030 18932 15036
rect 26240 15088 26292 15094
rect 26240 15030 26292 15036
rect 18144 14952 18196 14958
rect 18144 14894 18196 14900
rect 17370 14716 17678 14725
rect 17370 14714 17376 14716
rect 17432 14714 17456 14716
rect 17512 14714 17536 14716
rect 17592 14714 17616 14716
rect 17672 14714 17678 14716
rect 17432 14662 17434 14714
rect 17614 14662 17616 14714
rect 17370 14660 17376 14662
rect 17432 14660 17456 14662
rect 17512 14660 17536 14662
rect 17592 14660 17616 14662
rect 17672 14660 17678 14662
rect 17370 14651 17678 14660
rect 18156 14482 18184 14894
rect 18420 14816 18472 14822
rect 18420 14758 18472 14764
rect 18144 14476 18196 14482
rect 18144 14418 18196 14424
rect 18052 14272 18104 14278
rect 18052 14214 18104 14220
rect 17960 14068 18012 14074
rect 17960 14010 18012 14016
rect 17224 13932 17276 13938
rect 17224 13874 17276 13880
rect 17236 12850 17264 13874
rect 17370 13628 17678 13637
rect 17370 13626 17376 13628
rect 17432 13626 17456 13628
rect 17512 13626 17536 13628
rect 17592 13626 17616 13628
rect 17672 13626 17678 13628
rect 17432 13574 17434 13626
rect 17614 13574 17616 13626
rect 17370 13572 17376 13574
rect 17432 13572 17456 13574
rect 17512 13572 17536 13574
rect 17592 13572 17616 13574
rect 17672 13572 17678 13574
rect 17370 13563 17678 13572
rect 17972 13258 18000 14010
rect 17960 13252 18012 13258
rect 17960 13194 18012 13200
rect 18064 13190 18092 14214
rect 18156 14006 18184 14418
rect 18432 14278 18460 14758
rect 18892 14550 18920 15030
rect 20076 14952 20128 14958
rect 20076 14894 20128 14900
rect 18880 14544 18932 14550
rect 18880 14486 18932 14492
rect 18696 14408 18748 14414
rect 18696 14350 18748 14356
rect 18420 14272 18472 14278
rect 18420 14214 18472 14220
rect 18144 14000 18196 14006
rect 18144 13942 18196 13948
rect 18156 13394 18184 13942
rect 18144 13388 18196 13394
rect 18144 13330 18196 13336
rect 18052 13184 18104 13190
rect 18052 13126 18104 13132
rect 18156 12850 18184 13330
rect 17224 12844 17276 12850
rect 17224 12786 17276 12792
rect 18144 12844 18196 12850
rect 18144 12786 18196 12792
rect 17960 12776 18012 12782
rect 17960 12718 18012 12724
rect 17370 12540 17678 12549
rect 17370 12538 17376 12540
rect 17432 12538 17456 12540
rect 17512 12538 17536 12540
rect 17592 12538 17616 12540
rect 17672 12538 17678 12540
rect 17432 12486 17434 12538
rect 17614 12486 17616 12538
rect 17370 12484 17376 12486
rect 17432 12484 17456 12486
rect 17512 12484 17536 12486
rect 17592 12484 17616 12486
rect 17672 12484 17678 12486
rect 17370 12475 17678 12484
rect 17224 12300 17276 12306
rect 17224 12242 17276 12248
rect 17132 12096 17184 12102
rect 17132 12038 17184 12044
rect 17040 11688 17092 11694
rect 17040 11630 17092 11636
rect 16856 11552 16908 11558
rect 16856 11494 16908 11500
rect 16764 11144 16816 11150
rect 16764 11086 16816 11092
rect 16580 10804 16632 10810
rect 16580 10746 16632 10752
rect 16776 10198 16804 11086
rect 16868 10742 16896 11494
rect 17052 10810 17080 11630
rect 17144 11354 17172 12038
rect 17132 11348 17184 11354
rect 17132 11290 17184 11296
rect 17144 10810 17172 11290
rect 17236 11014 17264 12242
rect 17972 12238 18000 12718
rect 17500 12232 17552 12238
rect 17500 12174 17552 12180
rect 17960 12232 18012 12238
rect 17960 12174 18012 12180
rect 17512 11694 17540 12174
rect 17500 11688 17552 11694
rect 17500 11630 17552 11636
rect 17370 11452 17678 11461
rect 17370 11450 17376 11452
rect 17432 11450 17456 11452
rect 17512 11450 17536 11452
rect 17592 11450 17616 11452
rect 17672 11450 17678 11452
rect 17432 11398 17434 11450
rect 17614 11398 17616 11450
rect 17370 11396 17376 11398
rect 17432 11396 17456 11398
rect 17512 11396 17536 11398
rect 17592 11396 17616 11398
rect 17672 11396 17678 11398
rect 17370 11387 17678 11396
rect 17868 11348 17920 11354
rect 17868 11290 17920 11296
rect 17224 11008 17276 11014
rect 17224 10950 17276 10956
rect 17040 10804 17092 10810
rect 17040 10746 17092 10752
rect 17132 10804 17184 10810
rect 17132 10746 17184 10752
rect 16856 10736 16908 10742
rect 16856 10678 16908 10684
rect 17236 10674 17264 10950
rect 17224 10668 17276 10674
rect 17224 10610 17276 10616
rect 17370 10364 17678 10373
rect 17370 10362 17376 10364
rect 17432 10362 17456 10364
rect 17512 10362 17536 10364
rect 17592 10362 17616 10364
rect 17672 10362 17678 10364
rect 17432 10310 17434 10362
rect 17614 10310 17616 10362
rect 17370 10308 17376 10310
rect 17432 10308 17456 10310
rect 17512 10308 17536 10310
rect 17592 10308 17616 10310
rect 17672 10308 17678 10310
rect 17370 10299 17678 10308
rect 16764 10192 16816 10198
rect 16764 10134 16816 10140
rect 16776 9518 16804 10134
rect 16764 9512 16816 9518
rect 16764 9454 16816 9460
rect 16396 9444 16448 9450
rect 16396 9386 16448 9392
rect 16948 9376 17000 9382
rect 16948 9318 17000 9324
rect 17776 9376 17828 9382
rect 17776 9318 17828 9324
rect 16120 9172 16172 9178
rect 16120 9114 16172 9120
rect 15660 8628 15712 8634
rect 15660 8570 15712 8576
rect 15476 5364 15528 5370
rect 15476 5306 15528 5312
rect 15672 4622 15700 8570
rect 16132 8498 16160 9114
rect 16960 9042 16988 9318
rect 17370 9276 17678 9285
rect 17370 9274 17376 9276
rect 17432 9274 17456 9276
rect 17512 9274 17536 9276
rect 17592 9274 17616 9276
rect 17672 9274 17678 9276
rect 17432 9222 17434 9274
rect 17614 9222 17616 9274
rect 17370 9220 17376 9222
rect 17432 9220 17456 9222
rect 17512 9220 17536 9222
rect 17592 9220 17616 9222
rect 17672 9220 17678 9222
rect 17370 9211 17678 9220
rect 16948 9036 17000 9042
rect 16948 8978 17000 8984
rect 16856 8968 16908 8974
rect 16856 8910 16908 8916
rect 17132 8968 17184 8974
rect 17132 8910 17184 8916
rect 16212 8832 16264 8838
rect 16212 8774 16264 8780
rect 16120 8492 16172 8498
rect 16120 8434 16172 8440
rect 16132 7886 16160 8434
rect 16224 8430 16252 8774
rect 16212 8424 16264 8430
rect 16212 8366 16264 8372
rect 16120 7880 16172 7886
rect 16120 7822 16172 7828
rect 16868 7546 16896 8910
rect 17144 8566 17172 8910
rect 17788 8906 17816 9318
rect 17776 8900 17828 8906
rect 17776 8842 17828 8848
rect 17132 8560 17184 8566
rect 17132 8502 17184 8508
rect 17224 8560 17276 8566
rect 17224 8502 17276 8508
rect 17144 7886 17172 8502
rect 17236 8294 17264 8502
rect 17224 8288 17276 8294
rect 17224 8230 17276 8236
rect 17370 8188 17678 8197
rect 17370 8186 17376 8188
rect 17432 8186 17456 8188
rect 17512 8186 17536 8188
rect 17592 8186 17616 8188
rect 17672 8186 17678 8188
rect 17432 8134 17434 8186
rect 17614 8134 17616 8186
rect 17370 8132 17376 8134
rect 17432 8132 17456 8134
rect 17512 8132 17536 8134
rect 17592 8132 17616 8134
rect 17672 8132 17678 8134
rect 17370 8123 17678 8132
rect 17132 7880 17184 7886
rect 17132 7822 17184 7828
rect 16856 7540 16908 7546
rect 16856 7482 16908 7488
rect 16028 6112 16080 6118
rect 16028 6054 16080 6060
rect 16040 5710 16068 6054
rect 17144 5778 17172 7822
rect 17880 7546 17908 11290
rect 18432 10130 18460 14214
rect 18512 13864 18564 13870
rect 18512 13806 18564 13812
rect 18524 13530 18552 13806
rect 18512 13524 18564 13530
rect 18512 13466 18564 13472
rect 18512 12844 18564 12850
rect 18512 12786 18564 12792
rect 18524 12306 18552 12786
rect 18512 12300 18564 12306
rect 18512 12242 18564 12248
rect 18524 11150 18552 12242
rect 18708 12238 18736 14350
rect 19524 14272 19576 14278
rect 19524 14214 19576 14220
rect 19536 14006 19564 14214
rect 20088 14074 20116 14894
rect 20444 14816 20496 14822
rect 20444 14758 20496 14764
rect 22836 14816 22888 14822
rect 22836 14758 22888 14764
rect 25136 14816 25188 14822
rect 25136 14758 25188 14764
rect 20168 14340 20220 14346
rect 20168 14282 20220 14288
rect 20260 14340 20312 14346
rect 20260 14282 20312 14288
rect 20180 14074 20208 14282
rect 20076 14068 20128 14074
rect 20076 14010 20128 14016
rect 20168 14068 20220 14074
rect 20168 14010 20220 14016
rect 19524 14000 19576 14006
rect 19524 13942 19576 13948
rect 20272 13938 20300 14282
rect 20456 14006 20484 14758
rect 22560 14408 22612 14414
rect 22560 14350 22612 14356
rect 22376 14272 22428 14278
rect 22376 14214 22428 14220
rect 20444 14000 20496 14006
rect 20444 13942 20496 13948
rect 20260 13932 20312 13938
rect 20260 13874 20312 13880
rect 19984 13728 20036 13734
rect 19984 13670 20036 13676
rect 19996 13326 20024 13670
rect 20272 13462 20300 13874
rect 20456 13530 20484 13942
rect 20628 13932 20680 13938
rect 20628 13874 20680 13880
rect 21180 13932 21232 13938
rect 21180 13874 21232 13880
rect 20444 13524 20496 13530
rect 20444 13466 20496 13472
rect 20260 13456 20312 13462
rect 20260 13398 20312 13404
rect 20640 13326 20668 13874
rect 20812 13864 20864 13870
rect 20812 13806 20864 13812
rect 20720 13388 20772 13394
rect 20824 13376 20852 13806
rect 21192 13530 21220 13874
rect 21272 13864 21324 13870
rect 21272 13806 21324 13812
rect 21180 13524 21232 13530
rect 21180 13466 21232 13472
rect 20772 13348 20852 13376
rect 20720 13330 20772 13336
rect 19984 13320 20036 13326
rect 19984 13262 20036 13268
rect 20628 13320 20680 13326
rect 20628 13262 20680 13268
rect 18696 12232 18748 12238
rect 18696 12174 18748 12180
rect 18512 11144 18564 11150
rect 18512 11086 18564 11092
rect 18708 10810 18736 12174
rect 19996 11898 20024 13262
rect 20640 12646 20668 13262
rect 20720 13252 20772 13258
rect 20720 13194 20772 13200
rect 20628 12640 20680 12646
rect 20628 12582 20680 12588
rect 19984 11892 20036 11898
rect 19984 11834 20036 11840
rect 20640 11694 20668 12582
rect 20732 12442 20760 13194
rect 20824 12986 20852 13348
rect 20996 13184 21048 13190
rect 20996 13126 21048 13132
rect 20812 12980 20864 12986
rect 20812 12922 20864 12928
rect 20824 12782 20852 12922
rect 20904 12844 20956 12850
rect 20904 12786 20956 12792
rect 20812 12776 20864 12782
rect 20812 12718 20864 12724
rect 20720 12436 20772 12442
rect 20720 12378 20772 12384
rect 20916 12374 20944 12786
rect 20904 12368 20956 12374
rect 20904 12310 20956 12316
rect 21008 11762 21036 13126
rect 21088 12844 21140 12850
rect 21088 12786 21140 12792
rect 20996 11756 21048 11762
rect 20996 11698 21048 11704
rect 20260 11688 20312 11694
rect 20260 11630 20312 11636
rect 20628 11688 20680 11694
rect 20628 11630 20680 11636
rect 19708 11552 19760 11558
rect 19708 11494 19760 11500
rect 19720 11218 19748 11494
rect 19708 11212 19760 11218
rect 19708 11154 19760 11160
rect 18696 10804 18748 10810
rect 18696 10746 18748 10752
rect 20272 10742 20300 11630
rect 20996 11552 21048 11558
rect 20996 11494 21048 11500
rect 20812 11144 20864 11150
rect 20812 11086 20864 11092
rect 20824 10810 20852 11086
rect 20812 10804 20864 10810
rect 20812 10746 20864 10752
rect 20260 10736 20312 10742
rect 20260 10678 20312 10684
rect 19432 10668 19484 10674
rect 19432 10610 19484 10616
rect 20168 10668 20220 10674
rect 20168 10610 20220 10616
rect 18696 10464 18748 10470
rect 18696 10406 18748 10412
rect 18420 10124 18472 10130
rect 18420 10066 18472 10072
rect 17960 10056 18012 10062
rect 17960 9998 18012 10004
rect 17972 9586 18000 9998
rect 18052 9920 18104 9926
rect 18052 9862 18104 9868
rect 18420 9920 18472 9926
rect 18420 9862 18472 9868
rect 18064 9654 18092 9862
rect 18052 9648 18104 9654
rect 18052 9590 18104 9596
rect 17960 9580 18012 9586
rect 17960 9522 18012 9528
rect 17972 9178 18000 9522
rect 18432 9178 18460 9862
rect 18708 9586 18736 10406
rect 19156 10124 19208 10130
rect 19156 10066 19208 10072
rect 18696 9580 18748 9586
rect 18696 9522 18748 9528
rect 17960 9172 18012 9178
rect 17960 9114 18012 9120
rect 18420 9172 18472 9178
rect 18420 9114 18472 9120
rect 19064 9172 19116 9178
rect 19064 9114 19116 9120
rect 19076 8498 19104 9114
rect 19168 9042 19196 10066
rect 19444 9178 19472 10610
rect 19524 9920 19576 9926
rect 19524 9862 19576 9868
rect 19536 9654 19564 9862
rect 19524 9648 19576 9654
rect 19524 9590 19576 9596
rect 19432 9172 19484 9178
rect 19432 9114 19484 9120
rect 19156 9036 19208 9042
rect 19156 8978 19208 8984
rect 19064 8492 19116 8498
rect 19064 8434 19116 8440
rect 18604 8356 18656 8362
rect 18604 8298 18656 8304
rect 18144 7948 18196 7954
rect 18144 7890 18196 7896
rect 18156 7546 18184 7890
rect 17868 7540 17920 7546
rect 17868 7482 17920 7488
rect 18144 7540 18196 7546
rect 18144 7482 18196 7488
rect 18616 7478 18644 8298
rect 17224 7472 17276 7478
rect 17224 7414 17276 7420
rect 18604 7472 18656 7478
rect 18604 7414 18656 7420
rect 17236 6798 17264 7414
rect 18328 7336 18380 7342
rect 18328 7278 18380 7284
rect 17370 7100 17678 7109
rect 17370 7098 17376 7100
rect 17432 7098 17456 7100
rect 17512 7098 17536 7100
rect 17592 7098 17616 7100
rect 17672 7098 17678 7100
rect 17432 7046 17434 7098
rect 17614 7046 17616 7098
rect 17370 7044 17376 7046
rect 17432 7044 17456 7046
rect 17512 7044 17536 7046
rect 17592 7044 17616 7046
rect 17672 7044 17678 7046
rect 17370 7035 17678 7044
rect 17224 6792 17276 6798
rect 17224 6734 17276 6740
rect 17774 6352 17830 6361
rect 17774 6287 17830 6296
rect 17788 6254 17816 6287
rect 18340 6254 18368 7278
rect 18420 6928 18472 6934
rect 18420 6870 18472 6876
rect 18432 6798 18460 6870
rect 18616 6798 18644 7414
rect 18880 7404 18932 7410
rect 18880 7346 18932 7352
rect 18892 6866 18920 7346
rect 19168 7342 19196 8978
rect 19800 8492 19852 8498
rect 19800 8434 19852 8440
rect 19892 8492 19944 8498
rect 19892 8434 19944 8440
rect 19812 7954 19840 8434
rect 19800 7948 19852 7954
rect 19800 7890 19852 7896
rect 19904 7886 19932 8434
rect 20076 8288 20128 8294
rect 20076 8230 20128 8236
rect 19892 7880 19944 7886
rect 19892 7822 19944 7828
rect 19340 7744 19392 7750
rect 19340 7686 19392 7692
rect 19352 7546 19380 7686
rect 19340 7540 19392 7546
rect 19340 7482 19392 7488
rect 19156 7336 19208 7342
rect 19156 7278 19208 7284
rect 18788 6860 18840 6866
rect 18788 6802 18840 6808
rect 18880 6860 18932 6866
rect 18880 6802 18932 6808
rect 18420 6792 18472 6798
rect 18420 6734 18472 6740
rect 18512 6792 18564 6798
rect 18512 6734 18564 6740
rect 18604 6792 18656 6798
rect 18604 6734 18656 6740
rect 18432 6390 18460 6734
rect 18524 6662 18552 6734
rect 18512 6656 18564 6662
rect 18512 6598 18564 6604
rect 18420 6384 18472 6390
rect 18420 6326 18472 6332
rect 18604 6384 18656 6390
rect 18604 6326 18656 6332
rect 17776 6248 17828 6254
rect 17776 6190 17828 6196
rect 18328 6248 18380 6254
rect 18328 6190 18380 6196
rect 17370 6012 17678 6021
rect 17370 6010 17376 6012
rect 17432 6010 17456 6012
rect 17512 6010 17536 6012
rect 17592 6010 17616 6012
rect 17672 6010 17678 6012
rect 17432 5958 17434 6010
rect 17614 5958 17616 6010
rect 17370 5956 17376 5958
rect 17432 5956 17456 5958
rect 17512 5956 17536 5958
rect 17592 5956 17616 5958
rect 17672 5956 17678 5958
rect 17370 5947 17678 5956
rect 18340 5846 18368 6190
rect 18432 5914 18460 6326
rect 18420 5908 18472 5914
rect 18420 5850 18472 5856
rect 18328 5840 18380 5846
rect 18328 5782 18380 5788
rect 17132 5772 17184 5778
rect 17132 5714 17184 5720
rect 16028 5704 16080 5710
rect 16028 5646 16080 5652
rect 16764 5636 16816 5642
rect 16764 5578 16816 5584
rect 16580 5568 16632 5574
rect 16776 5522 16804 5578
rect 16632 5516 16804 5522
rect 16580 5510 16804 5516
rect 16592 5494 16804 5510
rect 17144 5302 17172 5714
rect 18616 5370 18644 6326
rect 18800 6322 18828 6802
rect 18788 6316 18840 6322
rect 18788 6258 18840 6264
rect 19168 6254 19196 7278
rect 19352 7002 19380 7482
rect 19904 7206 19932 7822
rect 19984 7744 20036 7750
rect 19984 7686 20036 7692
rect 19892 7200 19944 7206
rect 19892 7142 19944 7148
rect 19340 6996 19392 7002
rect 19340 6938 19392 6944
rect 19616 6792 19668 6798
rect 19892 6792 19944 6798
rect 19668 6752 19748 6780
rect 19616 6734 19668 6740
rect 19720 6322 19748 6752
rect 19892 6734 19944 6740
rect 19904 6458 19932 6734
rect 19892 6452 19944 6458
rect 19892 6394 19944 6400
rect 19904 6322 19932 6394
rect 19996 6322 20024 7686
rect 20088 7410 20116 8230
rect 20180 7546 20208 10610
rect 20720 9376 20772 9382
rect 20720 9318 20772 9324
rect 20732 8906 20760 9318
rect 21008 9110 21036 11494
rect 21100 11014 21128 12786
rect 21284 12714 21312 13806
rect 21548 13388 21600 13394
rect 21548 13330 21600 13336
rect 22008 13388 22060 13394
rect 22008 13330 22060 13336
rect 21456 13320 21508 13326
rect 21456 13262 21508 13268
rect 21468 12782 21496 13262
rect 21456 12776 21508 12782
rect 21456 12718 21508 12724
rect 21560 12714 21588 13330
rect 22020 12850 22048 13330
rect 22284 13320 22336 13326
rect 22284 13262 22336 13268
rect 22192 12980 22244 12986
rect 22192 12922 22244 12928
rect 22008 12844 22060 12850
rect 22008 12786 22060 12792
rect 22204 12782 22232 12922
rect 22192 12776 22244 12782
rect 22192 12718 22244 12724
rect 22296 12714 22324 13262
rect 21272 12708 21324 12714
rect 21272 12650 21324 12656
rect 21548 12708 21600 12714
rect 21548 12650 21600 12656
rect 22284 12708 22336 12714
rect 22284 12650 22336 12656
rect 22100 12640 22152 12646
rect 22100 12582 22152 12588
rect 21916 12436 21968 12442
rect 21968 12396 22048 12424
rect 21916 12378 21968 12384
rect 21824 12232 21876 12238
rect 21824 12174 21876 12180
rect 21456 12096 21508 12102
rect 21456 12038 21508 12044
rect 21468 11762 21496 12038
rect 21456 11756 21508 11762
rect 21456 11698 21508 11704
rect 21468 11354 21496 11698
rect 21836 11354 21864 12174
rect 21916 12164 21968 12170
rect 22020 12152 22048 12396
rect 22112 12306 22140 12582
rect 22100 12300 22152 12306
rect 22100 12242 22152 12248
rect 22100 12164 22152 12170
rect 22020 12124 22100 12152
rect 21916 12106 21968 12112
rect 22100 12106 22152 12112
rect 21928 11830 21956 12106
rect 21916 11824 21968 11830
rect 21916 11766 21968 11772
rect 22112 11762 22140 12106
rect 22296 11762 22324 12650
rect 22100 11756 22152 11762
rect 22100 11698 22152 11704
rect 22284 11756 22336 11762
rect 22284 11698 22336 11704
rect 21456 11348 21508 11354
rect 21456 11290 21508 11296
rect 21824 11348 21876 11354
rect 21824 11290 21876 11296
rect 21088 11008 21140 11014
rect 21088 10950 21140 10956
rect 21100 10810 21128 10950
rect 21088 10804 21140 10810
rect 21088 10746 21140 10752
rect 21180 10600 21232 10606
rect 21180 10542 21232 10548
rect 21192 10062 21220 10542
rect 22192 10464 22244 10470
rect 22192 10406 22244 10412
rect 21180 10056 21232 10062
rect 21180 9998 21232 10004
rect 22204 9994 22232 10406
rect 22192 9988 22244 9994
rect 22192 9930 22244 9936
rect 20996 9104 21048 9110
rect 20996 9046 21048 9052
rect 21916 9104 21968 9110
rect 21916 9046 21968 9052
rect 21548 8968 21600 8974
rect 21548 8910 21600 8916
rect 20720 8900 20772 8906
rect 20720 8842 20772 8848
rect 21088 8900 21140 8906
rect 21088 8842 21140 8848
rect 20260 8560 20312 8566
rect 20260 8502 20312 8508
rect 20272 7886 20300 8502
rect 20732 8498 20760 8842
rect 21100 8566 21128 8842
rect 21088 8560 21140 8566
rect 21088 8502 21140 8508
rect 20352 8492 20404 8498
rect 20352 8434 20404 8440
rect 20720 8492 20772 8498
rect 20720 8434 20772 8440
rect 20364 7954 20392 8434
rect 20352 7948 20404 7954
rect 20352 7890 20404 7896
rect 21100 7886 21128 8502
rect 21560 7954 21588 8910
rect 21548 7948 21600 7954
rect 21548 7890 21600 7896
rect 20260 7880 20312 7886
rect 20260 7822 20312 7828
rect 21088 7880 21140 7886
rect 21088 7822 21140 7828
rect 20720 7744 20772 7750
rect 20720 7686 20772 7692
rect 20996 7744 21048 7750
rect 20996 7686 21048 7692
rect 20168 7540 20220 7546
rect 20168 7482 20220 7488
rect 20732 7410 20760 7686
rect 21008 7546 21036 7686
rect 20996 7540 21048 7546
rect 20996 7482 21048 7488
rect 20076 7404 20128 7410
rect 20076 7346 20128 7352
rect 20720 7404 20772 7410
rect 20720 7346 20772 7352
rect 20996 7336 21048 7342
rect 20732 7262 20944 7290
rect 20996 7278 21048 7284
rect 20732 7206 20760 7262
rect 20720 7200 20772 7206
rect 20720 7142 20772 7148
rect 20812 7200 20864 7206
rect 20812 7142 20864 7148
rect 20720 6724 20772 6730
rect 20720 6666 20772 6672
rect 19708 6316 19760 6322
rect 19708 6258 19760 6264
rect 19892 6316 19944 6322
rect 19892 6258 19944 6264
rect 19984 6316 20036 6322
rect 19984 6258 20036 6264
rect 18972 6248 19024 6254
rect 18972 6190 19024 6196
rect 19156 6248 19208 6254
rect 19156 6190 19208 6196
rect 18696 5704 18748 5710
rect 18696 5646 18748 5652
rect 18604 5364 18656 5370
rect 18604 5306 18656 5312
rect 17132 5296 17184 5302
rect 17132 5238 17184 5244
rect 18420 5296 18472 5302
rect 18420 5238 18472 5244
rect 15660 4616 15712 4622
rect 15660 4558 15712 4564
rect 17144 4554 17172 5238
rect 17370 4924 17678 4933
rect 17370 4922 17376 4924
rect 17432 4922 17456 4924
rect 17512 4922 17536 4924
rect 17592 4922 17616 4924
rect 17672 4922 17678 4924
rect 17432 4870 17434 4922
rect 17614 4870 17616 4922
rect 17370 4868 17376 4870
rect 17432 4868 17456 4870
rect 17512 4868 17536 4870
rect 17592 4868 17616 4870
rect 17672 4868 17678 4870
rect 17370 4859 17678 4868
rect 18432 4826 18460 5238
rect 18420 4820 18472 4826
rect 18420 4762 18472 4768
rect 18708 4622 18736 5646
rect 18984 4758 19012 6190
rect 19168 5846 19196 6190
rect 19720 6118 19748 6258
rect 20352 6248 20404 6254
rect 20352 6190 20404 6196
rect 19248 6112 19300 6118
rect 19248 6054 19300 6060
rect 19708 6112 19760 6118
rect 19708 6054 19760 6060
rect 19156 5840 19208 5846
rect 19156 5782 19208 5788
rect 19260 5234 19288 6054
rect 20364 5778 20392 6190
rect 20732 5930 20760 6666
rect 20824 6458 20852 7142
rect 20812 6452 20864 6458
rect 20812 6394 20864 6400
rect 20916 6186 20944 7262
rect 21008 6662 21036 7278
rect 20996 6656 21048 6662
rect 20996 6598 21048 6604
rect 21456 6656 21508 6662
rect 21456 6598 21508 6604
rect 20996 6452 21048 6458
rect 20996 6394 21048 6400
rect 20812 6180 20864 6186
rect 20812 6122 20864 6128
rect 20904 6180 20956 6186
rect 20904 6122 20956 6128
rect 20824 6066 20852 6122
rect 21008 6066 21036 6394
rect 21468 6390 21496 6598
rect 21456 6384 21508 6390
rect 21456 6326 21508 6332
rect 21560 6322 21588 7890
rect 21928 7478 21956 9046
rect 22008 8492 22060 8498
rect 22008 8434 22060 8440
rect 22020 7750 22048 8434
rect 22192 8288 22244 8294
rect 22192 8230 22244 8236
rect 22008 7744 22060 7750
rect 22008 7686 22060 7692
rect 21916 7472 21968 7478
rect 21916 7414 21968 7420
rect 21824 6792 21876 6798
rect 21652 6740 21824 6746
rect 21652 6734 21876 6740
rect 21928 6780 21956 7414
rect 22204 7206 22232 8230
rect 22388 7970 22416 14214
rect 22572 13938 22600 14350
rect 22848 14278 22876 14758
rect 22836 14272 22888 14278
rect 22836 14214 22888 14220
rect 22843 14172 23151 14181
rect 22843 14170 22849 14172
rect 22905 14170 22929 14172
rect 22985 14170 23009 14172
rect 23065 14170 23089 14172
rect 23145 14170 23151 14172
rect 22905 14118 22907 14170
rect 23087 14118 23089 14170
rect 22843 14116 22849 14118
rect 22905 14116 22929 14118
rect 22985 14116 23009 14118
rect 23065 14116 23089 14118
rect 23145 14116 23151 14118
rect 22843 14107 23151 14116
rect 25148 14074 25176 14758
rect 25136 14068 25188 14074
rect 25136 14010 25188 14016
rect 22468 13932 22520 13938
rect 22468 13874 22520 13880
rect 22560 13932 22612 13938
rect 22560 13874 22612 13880
rect 22480 12986 22508 13874
rect 24768 13728 24820 13734
rect 24768 13670 24820 13676
rect 22652 13388 22704 13394
rect 22652 13330 22704 13336
rect 22664 13258 22692 13330
rect 24584 13320 24636 13326
rect 24584 13262 24636 13268
rect 22652 13252 22704 13258
rect 22652 13194 22704 13200
rect 22468 12980 22520 12986
rect 22468 12922 22520 12928
rect 22664 12646 22692 13194
rect 22843 13084 23151 13093
rect 22843 13082 22849 13084
rect 22905 13082 22929 13084
rect 22985 13082 23009 13084
rect 23065 13082 23089 13084
rect 23145 13082 23151 13084
rect 22905 13030 22907 13082
rect 23087 13030 23089 13082
rect 22843 13028 22849 13030
rect 22905 13028 22929 13030
rect 22985 13028 23009 13030
rect 23065 13028 23089 13030
rect 23145 13028 23151 13030
rect 22843 13019 23151 13028
rect 23112 12708 23164 12714
rect 23112 12650 23164 12656
rect 22652 12640 22704 12646
rect 22652 12582 22704 12588
rect 23124 12238 23152 12650
rect 24596 12306 24624 13262
rect 24780 12889 24808 13670
rect 24766 12880 24822 12889
rect 24766 12815 24822 12824
rect 25228 12844 25280 12850
rect 25228 12786 25280 12792
rect 25964 12844 26016 12850
rect 25964 12786 26016 12792
rect 24676 12776 24728 12782
rect 24676 12718 24728 12724
rect 24584 12300 24636 12306
rect 24584 12242 24636 12248
rect 23112 12232 23164 12238
rect 23112 12174 23164 12180
rect 22744 12096 22796 12102
rect 22744 12038 22796 12044
rect 22756 11898 22784 12038
rect 22843 11996 23151 12005
rect 22843 11994 22849 11996
rect 22905 11994 22929 11996
rect 22985 11994 23009 11996
rect 23065 11994 23089 11996
rect 23145 11994 23151 11996
rect 22905 11942 22907 11994
rect 23087 11942 23089 11994
rect 22843 11940 22849 11942
rect 22905 11940 22929 11942
rect 22985 11940 23009 11942
rect 23065 11940 23089 11942
rect 23145 11940 23151 11942
rect 22843 11931 23151 11940
rect 22744 11892 22796 11898
rect 22744 11834 22796 11840
rect 22836 11756 22888 11762
rect 22836 11698 22888 11704
rect 22652 11552 22704 11558
rect 22652 11494 22704 11500
rect 22664 11150 22692 11494
rect 22848 11286 22876 11698
rect 22836 11280 22888 11286
rect 22836 11222 22888 11228
rect 24688 11150 24716 12718
rect 24860 12300 24912 12306
rect 24860 12242 24912 12248
rect 24872 11694 24900 12242
rect 25136 12096 25188 12102
rect 25136 12038 25188 12044
rect 25148 11830 25176 12038
rect 25044 11824 25096 11830
rect 25044 11766 25096 11772
rect 25136 11824 25188 11830
rect 25136 11766 25188 11772
rect 24860 11688 24912 11694
rect 24860 11630 24912 11636
rect 24768 11620 24820 11626
rect 24768 11562 24820 11568
rect 24780 11218 24808 11562
rect 24768 11212 24820 11218
rect 24768 11154 24820 11160
rect 22652 11144 22704 11150
rect 22652 11086 22704 11092
rect 24676 11144 24728 11150
rect 24676 11086 24728 11092
rect 23204 11008 23256 11014
rect 23204 10950 23256 10956
rect 22843 10908 23151 10917
rect 22843 10906 22849 10908
rect 22905 10906 22929 10908
rect 22985 10906 23009 10908
rect 23065 10906 23089 10908
rect 23145 10906 23151 10908
rect 22905 10854 22907 10906
rect 23087 10854 23089 10906
rect 22843 10852 22849 10854
rect 22905 10852 22929 10854
rect 22985 10852 23009 10854
rect 23065 10852 23089 10854
rect 23145 10852 23151 10854
rect 22843 10843 23151 10852
rect 22652 10804 22704 10810
rect 22652 10746 22704 10752
rect 22560 10600 22612 10606
rect 22560 10542 22612 10548
rect 22572 9586 22600 10542
rect 22664 9722 22692 10746
rect 23216 10742 23244 10950
rect 24780 10742 24808 11154
rect 23204 10736 23256 10742
rect 23204 10678 23256 10684
rect 24676 10736 24728 10742
rect 24676 10678 24728 10684
rect 24768 10736 24820 10742
rect 24768 10678 24820 10684
rect 24584 10600 24636 10606
rect 24584 10542 24636 10548
rect 24596 10266 24624 10542
rect 24688 10266 24716 10678
rect 24584 10260 24636 10266
rect 24584 10202 24636 10208
rect 24676 10260 24728 10266
rect 24676 10202 24728 10208
rect 22744 10192 22796 10198
rect 22744 10134 22796 10140
rect 22652 9716 22704 9722
rect 22652 9658 22704 9664
rect 22756 9654 22784 10134
rect 24872 10130 24900 11630
rect 25056 11218 25084 11766
rect 25044 11212 25096 11218
rect 25044 11154 25096 11160
rect 25240 11014 25268 12786
rect 25976 12730 26004 12786
rect 25884 12702 26004 12730
rect 25884 12442 25912 12702
rect 25872 12436 25924 12442
rect 25872 12378 25924 12384
rect 25504 12164 25556 12170
rect 25504 12106 25556 12112
rect 25516 11354 25544 12106
rect 25884 11898 25912 12378
rect 26148 12232 26200 12238
rect 26068 12192 26148 12220
rect 25872 11892 25924 11898
rect 25872 11834 25924 11840
rect 25504 11348 25556 11354
rect 25504 11290 25556 11296
rect 26068 11150 26096 12192
rect 26148 12174 26200 12180
rect 26148 11756 26200 11762
rect 26148 11698 26200 11704
rect 26160 11354 26188 11698
rect 26148 11348 26200 11354
rect 26148 11290 26200 11296
rect 25320 11144 25372 11150
rect 25320 11086 25372 11092
rect 25412 11144 25464 11150
rect 25412 11086 25464 11092
rect 25504 11144 25556 11150
rect 25504 11086 25556 11092
rect 26056 11144 26108 11150
rect 26056 11086 26108 11092
rect 24952 11008 25004 11014
rect 25228 11008 25280 11014
rect 24952 10950 25004 10956
rect 25148 10956 25228 10962
rect 25148 10950 25280 10956
rect 24964 10198 24992 10950
rect 25148 10934 25268 10950
rect 24952 10192 25004 10198
rect 24952 10134 25004 10140
rect 24860 10124 24912 10130
rect 24860 10066 24912 10072
rect 23572 9920 23624 9926
rect 23572 9862 23624 9868
rect 22843 9820 23151 9829
rect 22843 9818 22849 9820
rect 22905 9818 22929 9820
rect 22985 9818 23009 9820
rect 23065 9818 23089 9820
rect 23145 9818 23151 9820
rect 22905 9766 22907 9818
rect 23087 9766 23089 9818
rect 22843 9764 22849 9766
rect 22905 9764 22929 9766
rect 22985 9764 23009 9766
rect 23065 9764 23089 9766
rect 23145 9764 23151 9766
rect 22843 9755 23151 9764
rect 23584 9654 23612 9862
rect 25148 9722 25176 10934
rect 25332 10810 25360 11086
rect 25228 10804 25280 10810
rect 25228 10746 25280 10752
rect 25320 10804 25372 10810
rect 25320 10746 25372 10752
rect 25240 10690 25268 10746
rect 25424 10690 25452 11086
rect 25240 10662 25452 10690
rect 25424 10538 25452 10662
rect 25412 10532 25464 10538
rect 25412 10474 25464 10480
rect 25320 10464 25372 10470
rect 25320 10406 25372 10412
rect 25332 9926 25360 10406
rect 25516 10062 25544 11086
rect 26252 11082 26280 15030
rect 26608 14952 26660 14958
rect 26608 14894 26660 14900
rect 26424 14340 26476 14346
rect 26424 14282 26476 14288
rect 26516 14340 26568 14346
rect 26516 14282 26568 14288
rect 26332 13932 26384 13938
rect 26332 13874 26384 13880
rect 26344 13530 26372 13874
rect 26436 13530 26464 14282
rect 26528 14006 26556 14282
rect 26516 14000 26568 14006
rect 26516 13942 26568 13948
rect 26332 13524 26384 13530
rect 26332 13466 26384 13472
rect 26424 13524 26476 13530
rect 26424 13466 26476 13472
rect 26344 13394 26372 13466
rect 26332 13388 26384 13394
rect 26332 13330 26384 13336
rect 26528 12306 26556 13942
rect 26516 12300 26568 12306
rect 26516 12242 26568 12248
rect 26240 11076 26292 11082
rect 26240 11018 26292 11024
rect 26056 11008 26108 11014
rect 26056 10950 26108 10956
rect 25780 10736 25832 10742
rect 25780 10678 25832 10684
rect 25504 10056 25556 10062
rect 25504 9998 25556 10004
rect 25320 9920 25372 9926
rect 25320 9862 25372 9868
rect 25136 9716 25188 9722
rect 25136 9658 25188 9664
rect 25332 9654 25360 9862
rect 22744 9648 22796 9654
rect 22744 9590 22796 9596
rect 23572 9648 23624 9654
rect 23572 9590 23624 9596
rect 25320 9648 25372 9654
rect 25320 9590 25372 9596
rect 22560 9580 22612 9586
rect 22560 9522 22612 9528
rect 25044 9376 25096 9382
rect 25044 9318 25096 9324
rect 25056 9042 25084 9318
rect 25044 9036 25096 9042
rect 25044 8978 25096 8984
rect 24584 8968 24636 8974
rect 24584 8910 24636 8916
rect 22744 8900 22796 8906
rect 22744 8842 22796 8848
rect 22652 8832 22704 8838
rect 22652 8774 22704 8780
rect 22388 7942 22508 7970
rect 22376 7880 22428 7886
rect 22376 7822 22428 7828
rect 22388 7546 22416 7822
rect 22376 7540 22428 7546
rect 22376 7482 22428 7488
rect 22192 7200 22244 7206
rect 22192 7142 22244 7148
rect 22008 6792 22060 6798
rect 21928 6752 22008 6780
rect 21652 6730 21864 6734
rect 21640 6724 21864 6730
rect 21692 6718 21864 6724
rect 21640 6666 21692 6672
rect 21548 6316 21600 6322
rect 21548 6258 21600 6264
rect 21180 6248 21232 6254
rect 21180 6190 21232 6196
rect 20824 6038 21036 6066
rect 20640 5902 20760 5930
rect 20824 5914 20944 5930
rect 20824 5908 20956 5914
rect 20824 5902 20904 5908
rect 20352 5772 20404 5778
rect 20352 5714 20404 5720
rect 20640 5710 20668 5902
rect 20536 5704 20588 5710
rect 20456 5652 20536 5658
rect 20456 5646 20588 5652
rect 20628 5704 20680 5710
rect 20824 5658 20852 5902
rect 20904 5850 20956 5856
rect 21008 5710 21036 6038
rect 20628 5646 20680 5652
rect 20456 5630 20576 5646
rect 20732 5630 20852 5658
rect 20996 5704 21048 5710
rect 20996 5646 21048 5652
rect 20456 5574 20484 5630
rect 20444 5568 20496 5574
rect 20732 5522 20760 5630
rect 21192 5574 21220 6190
rect 21560 5914 21588 6258
rect 21548 5908 21600 5914
rect 21548 5850 21600 5856
rect 20444 5510 20496 5516
rect 20548 5494 20760 5522
rect 20996 5568 21048 5574
rect 20996 5510 21048 5516
rect 21180 5568 21232 5574
rect 21180 5510 21232 5516
rect 19248 5228 19300 5234
rect 19248 5170 19300 5176
rect 18972 4752 19024 4758
rect 18972 4694 19024 4700
rect 20548 4690 20576 5494
rect 21008 5234 21036 5510
rect 21192 5234 21220 5510
rect 21836 5370 21864 6718
rect 21928 6458 21956 6752
rect 22008 6734 22060 6740
rect 21916 6452 21968 6458
rect 21916 6394 21968 6400
rect 21916 5908 21968 5914
rect 21916 5850 21968 5856
rect 21928 5710 21956 5850
rect 21916 5704 21968 5710
rect 21916 5646 21968 5652
rect 21824 5364 21876 5370
rect 21824 5306 21876 5312
rect 20996 5228 21048 5234
rect 20996 5170 21048 5176
rect 21180 5228 21232 5234
rect 21180 5170 21232 5176
rect 20536 4684 20588 4690
rect 20536 4626 20588 4632
rect 20812 4684 20864 4690
rect 20812 4626 20864 4632
rect 17960 4616 18012 4622
rect 17960 4558 18012 4564
rect 18696 4616 18748 4622
rect 18696 4558 18748 4564
rect 17132 4548 17184 4554
rect 17132 4490 17184 4496
rect 17868 4548 17920 4554
rect 17868 4490 17920 4496
rect 17592 4208 17644 4214
rect 17592 4150 17644 4156
rect 16764 4140 16816 4146
rect 16764 4082 16816 4088
rect 14280 4072 14332 4078
rect 14280 4014 14332 4020
rect 14556 4072 14608 4078
rect 14556 4014 14608 4020
rect 15292 4072 15344 4078
rect 15292 4014 15344 4020
rect 14568 3534 14596 4014
rect 15844 3936 15896 3942
rect 15844 3878 15896 3884
rect 14556 3528 14608 3534
rect 14556 3470 14608 3476
rect 14832 3528 14884 3534
rect 14832 3470 14884 3476
rect 14464 3392 14516 3398
rect 14464 3334 14516 3340
rect 14476 3058 14504 3334
rect 14844 3058 14872 3470
rect 15856 3126 15884 3878
rect 16580 3460 16632 3466
rect 16580 3402 16632 3408
rect 16592 3126 16620 3402
rect 15844 3120 15896 3126
rect 15844 3062 15896 3068
rect 16580 3120 16632 3126
rect 16580 3062 16632 3068
rect 14464 3052 14516 3058
rect 14464 2994 14516 3000
rect 14832 3052 14884 3058
rect 14832 2994 14884 3000
rect 16776 2990 16804 4082
rect 17604 3942 17632 4150
rect 17880 4078 17908 4490
rect 17972 4146 18000 4558
rect 19432 4480 19484 4486
rect 19432 4422 19484 4428
rect 19444 4214 19472 4422
rect 19432 4208 19484 4214
rect 19432 4150 19484 4156
rect 17960 4140 18012 4146
rect 17960 4082 18012 4088
rect 17868 4072 17920 4078
rect 17868 4014 17920 4020
rect 17592 3936 17644 3942
rect 17592 3878 17644 3884
rect 17370 3836 17678 3845
rect 17370 3834 17376 3836
rect 17432 3834 17456 3836
rect 17512 3834 17536 3836
rect 17592 3834 17616 3836
rect 17672 3834 17678 3836
rect 17432 3782 17434 3834
rect 17614 3782 17616 3834
rect 17370 3780 17376 3782
rect 17432 3780 17456 3782
rect 17512 3780 17536 3782
rect 17592 3780 17616 3782
rect 17672 3780 17678 3782
rect 17370 3771 17678 3780
rect 16868 3590 17080 3618
rect 16868 3194 16896 3590
rect 17052 3534 17080 3590
rect 17880 3534 17908 4014
rect 20548 3534 20576 4626
rect 20720 4548 20772 4554
rect 20720 4490 20772 4496
rect 20732 4214 20760 4490
rect 20720 4208 20772 4214
rect 20720 4150 20772 4156
rect 20824 4078 20852 4626
rect 22100 4548 22152 4554
rect 22100 4490 22152 4496
rect 22112 4146 22140 4490
rect 22100 4140 22152 4146
rect 22100 4082 22152 4088
rect 20812 4072 20864 4078
rect 20812 4014 20864 4020
rect 16948 3528 17000 3534
rect 16948 3470 17000 3476
rect 17040 3528 17092 3534
rect 17040 3470 17092 3476
rect 17868 3528 17920 3534
rect 17868 3470 17920 3476
rect 20536 3528 20588 3534
rect 20536 3470 20588 3476
rect 16960 3194 16988 3470
rect 17040 3392 17092 3398
rect 17040 3334 17092 3340
rect 16856 3188 16908 3194
rect 16856 3130 16908 3136
rect 16948 3188 17000 3194
rect 16948 3130 17000 3136
rect 16764 2984 16816 2990
rect 16764 2926 16816 2932
rect 14188 2848 14240 2854
rect 14188 2790 14240 2796
rect 12808 2508 12860 2514
rect 12808 2450 12860 2456
rect 1308 2440 1360 2446
rect 1308 2382 1360 2388
rect 4160 2440 4212 2446
rect 4160 2382 4212 2388
rect 4528 2440 4580 2446
rect 4528 2382 4580 2388
rect 5724 2440 5776 2446
rect 5724 2382 5776 2388
rect 7748 2440 7800 2446
rect 7748 2382 7800 2388
rect 9588 2440 9640 2446
rect 9588 2382 9640 2388
rect 11060 2440 11112 2446
rect 11060 2382 11112 2388
rect 12900 2440 12952 2446
rect 12900 2382 12952 2388
rect 938 1456 994 1465
rect 938 1391 994 1400
rect 1320 800 1348 2382
rect 4172 950 4200 2382
rect 3240 944 3292 950
rect 3240 886 3292 892
rect 4160 944 4212 950
rect 4160 886 4212 892
rect 3252 800 3280 886
rect 4540 800 4568 2382
rect 6460 2304 6512 2310
rect 6460 2246 6512 2252
rect 6472 800 6500 2246
rect 7760 800 7788 2382
rect 9680 2304 9732 2310
rect 9680 2246 9732 2252
rect 9692 800 9720 2246
rect 11072 898 11100 2382
rect 11896 2204 12204 2213
rect 11896 2202 11902 2204
rect 11958 2202 11982 2204
rect 12038 2202 12062 2204
rect 12118 2202 12142 2204
rect 12198 2202 12204 2204
rect 11958 2150 11960 2202
rect 12140 2150 12142 2202
rect 11896 2148 11902 2150
rect 11958 2148 11982 2150
rect 12038 2148 12062 2150
rect 12118 2148 12142 2150
rect 12198 2148 12204 2150
rect 11896 2139 12204 2148
rect 10980 870 11100 898
rect 10980 800 11008 870
rect 12912 800 12940 2382
rect 14200 800 14228 2790
rect 16776 2446 16804 2926
rect 17052 2774 17080 3334
rect 17880 3126 17908 3470
rect 18880 3460 18932 3466
rect 18880 3402 18932 3408
rect 22100 3460 22152 3466
rect 22100 3402 22152 3408
rect 18604 3392 18656 3398
rect 18604 3334 18656 3340
rect 17868 3120 17920 3126
rect 17868 3062 17920 3068
rect 18616 3058 18644 3334
rect 18892 3058 18920 3402
rect 22112 3194 22140 3402
rect 22100 3188 22152 3194
rect 22100 3130 22152 3136
rect 22480 3058 22508 7942
rect 22664 7410 22692 8774
rect 22756 7546 22784 8842
rect 24032 8832 24084 8838
rect 24032 8774 24084 8780
rect 22843 8732 23151 8741
rect 22843 8730 22849 8732
rect 22905 8730 22929 8732
rect 22985 8730 23009 8732
rect 23065 8730 23089 8732
rect 23145 8730 23151 8732
rect 22905 8678 22907 8730
rect 23087 8678 23089 8730
rect 22843 8676 22849 8678
rect 22905 8676 22929 8678
rect 22985 8676 23009 8678
rect 23065 8676 23089 8678
rect 23145 8676 23151 8678
rect 22843 8667 23151 8676
rect 24044 8566 24072 8774
rect 24032 8560 24084 8566
rect 24032 8502 24084 8508
rect 23388 8492 23440 8498
rect 23388 8434 23440 8440
rect 22843 7644 23151 7653
rect 22843 7642 22849 7644
rect 22905 7642 22929 7644
rect 22985 7642 23009 7644
rect 23065 7642 23089 7644
rect 23145 7642 23151 7644
rect 22905 7590 22907 7642
rect 23087 7590 23089 7642
rect 22843 7588 22849 7590
rect 22905 7588 22929 7590
rect 22985 7588 23009 7590
rect 23065 7588 23089 7590
rect 23145 7588 23151 7590
rect 22843 7579 23151 7588
rect 22744 7540 22796 7546
rect 22744 7482 22796 7488
rect 22652 7404 22704 7410
rect 22652 7346 22704 7352
rect 22652 6792 22704 6798
rect 22652 6734 22704 6740
rect 22664 6458 22692 6734
rect 22843 6556 23151 6565
rect 22843 6554 22849 6556
rect 22905 6554 22929 6556
rect 22985 6554 23009 6556
rect 23065 6554 23089 6556
rect 23145 6554 23151 6556
rect 22905 6502 22907 6554
rect 23087 6502 23089 6554
rect 22843 6500 22849 6502
rect 22905 6500 22929 6502
rect 22985 6500 23009 6502
rect 23065 6500 23089 6502
rect 23145 6500 23151 6502
rect 22843 6491 23151 6500
rect 22652 6452 22704 6458
rect 22652 6394 22704 6400
rect 22843 5468 23151 5477
rect 22843 5466 22849 5468
rect 22905 5466 22929 5468
rect 22985 5466 23009 5468
rect 23065 5466 23089 5468
rect 23145 5466 23151 5468
rect 22905 5414 22907 5466
rect 23087 5414 23089 5466
rect 22843 5412 22849 5414
rect 22905 5412 22929 5414
rect 22985 5412 23009 5414
rect 23065 5412 23089 5414
rect 23145 5412 23151 5414
rect 22843 5403 23151 5412
rect 23296 5228 23348 5234
rect 23296 5170 23348 5176
rect 23204 4480 23256 4486
rect 23204 4422 23256 4428
rect 22843 4380 23151 4389
rect 22843 4378 22849 4380
rect 22905 4378 22929 4380
rect 22985 4378 23009 4380
rect 23065 4378 23089 4380
rect 23145 4378 23151 4380
rect 22905 4326 22907 4378
rect 23087 4326 23089 4378
rect 22843 4324 22849 4326
rect 22905 4324 22929 4326
rect 22985 4324 23009 4326
rect 23065 4324 23089 4326
rect 23145 4324 23151 4326
rect 22843 4315 23151 4324
rect 23216 4146 23244 4422
rect 23204 4140 23256 4146
rect 23204 4082 23256 4088
rect 23308 4010 23336 5170
rect 23296 4004 23348 4010
rect 23296 3946 23348 3952
rect 23400 3602 23428 8434
rect 23940 8016 23992 8022
rect 23940 7958 23992 7964
rect 23756 7404 23808 7410
rect 23756 7346 23808 7352
rect 23768 3942 23796 7346
rect 23952 7342 23980 7958
rect 24044 7954 24072 8502
rect 24032 7948 24084 7954
rect 24032 7890 24084 7896
rect 23940 7336 23992 7342
rect 23940 7278 23992 7284
rect 23952 4214 23980 7278
rect 24596 6798 24624 8910
rect 25516 7886 25544 9998
rect 25792 9586 25820 10678
rect 26068 10674 26096 10950
rect 26148 10804 26200 10810
rect 26148 10746 26200 10752
rect 26056 10668 26108 10674
rect 26056 10610 26108 10616
rect 26160 9602 26188 10746
rect 26424 9988 26476 9994
rect 26424 9930 26476 9936
rect 26436 9722 26464 9930
rect 26424 9716 26476 9722
rect 26424 9658 26476 9664
rect 26160 9586 26280 9602
rect 25596 9580 25648 9586
rect 25596 9522 25648 9528
rect 25780 9580 25832 9586
rect 26160 9580 26292 9586
rect 26160 9574 26240 9580
rect 25780 9522 25832 9528
rect 26240 9522 26292 9528
rect 25608 8634 25636 9522
rect 25792 9042 25820 9522
rect 26620 9042 26648 14894
rect 27252 14612 27304 14618
rect 27252 14554 27304 14560
rect 27160 13932 27212 13938
rect 27160 13874 27212 13880
rect 26976 13728 27028 13734
rect 26976 13670 27028 13676
rect 26988 13326 27016 13670
rect 27172 13326 27200 13874
rect 26976 13320 27028 13326
rect 26976 13262 27028 13268
rect 27160 13320 27212 13326
rect 27160 13262 27212 13268
rect 26884 13252 26936 13258
rect 26884 13194 26936 13200
rect 26896 12442 26924 13194
rect 27172 12986 27200 13262
rect 27160 12980 27212 12986
rect 27160 12922 27212 12928
rect 26884 12436 26936 12442
rect 26884 12378 26936 12384
rect 27264 10674 27292 14554
rect 27528 14272 27580 14278
rect 27528 14214 27580 14220
rect 27540 14074 27568 14214
rect 27436 14068 27488 14074
rect 27436 14010 27488 14016
rect 27528 14068 27580 14074
rect 27528 14010 27580 14016
rect 27448 13802 27476 14010
rect 27528 13932 27580 13938
rect 27528 13874 27580 13880
rect 27436 13796 27488 13802
rect 27436 13738 27488 13744
rect 27448 10810 27476 13738
rect 27436 10804 27488 10810
rect 27436 10746 27488 10752
rect 27252 10668 27304 10674
rect 27252 10610 27304 10616
rect 27540 9110 27568 13874
rect 27632 13870 27660 16526
rect 28317 15804 28625 15813
rect 28317 15802 28323 15804
rect 28379 15802 28403 15804
rect 28459 15802 28483 15804
rect 28539 15802 28563 15804
rect 28619 15802 28625 15804
rect 28379 15750 28381 15802
rect 28561 15750 28563 15802
rect 28317 15748 28323 15750
rect 28379 15748 28403 15750
rect 28459 15748 28483 15750
rect 28539 15748 28563 15750
rect 28619 15748 28625 15750
rect 28317 15739 28625 15748
rect 28317 14716 28625 14725
rect 28317 14714 28323 14716
rect 28379 14714 28403 14716
rect 28459 14714 28483 14716
rect 28539 14714 28563 14716
rect 28619 14714 28625 14716
rect 28379 14662 28381 14714
rect 28561 14662 28563 14714
rect 28317 14660 28323 14662
rect 28379 14660 28403 14662
rect 28459 14660 28483 14662
rect 28539 14660 28563 14662
rect 28619 14660 28625 14662
rect 28317 14651 28625 14660
rect 30288 14612 30340 14618
rect 30288 14554 30340 14560
rect 29184 14408 29236 14414
rect 29184 14350 29236 14356
rect 29196 14006 29224 14350
rect 30300 14006 30328 14554
rect 29184 14000 29236 14006
rect 29184 13942 29236 13948
rect 30288 14000 30340 14006
rect 30288 13942 30340 13948
rect 27620 13864 27672 13870
rect 27620 13806 27672 13812
rect 28317 13628 28625 13637
rect 28317 13626 28323 13628
rect 28379 13626 28403 13628
rect 28459 13626 28483 13628
rect 28539 13626 28563 13628
rect 28619 13626 28625 13628
rect 28379 13574 28381 13626
rect 28561 13574 28563 13626
rect 28317 13572 28323 13574
rect 28379 13572 28403 13574
rect 28459 13572 28483 13574
rect 28539 13572 28563 13574
rect 28619 13572 28625 13574
rect 28317 13563 28625 13572
rect 28908 13320 28960 13326
rect 28908 13262 28960 13268
rect 28317 12540 28625 12549
rect 28317 12538 28323 12540
rect 28379 12538 28403 12540
rect 28459 12538 28483 12540
rect 28539 12538 28563 12540
rect 28619 12538 28625 12540
rect 28379 12486 28381 12538
rect 28561 12486 28563 12538
rect 28317 12484 28323 12486
rect 28379 12484 28403 12486
rect 28459 12484 28483 12486
rect 28539 12484 28563 12486
rect 28619 12484 28625 12486
rect 28317 12475 28625 12484
rect 28920 12306 28948 13262
rect 29196 12850 29224 13942
rect 29920 13864 29972 13870
rect 29920 13806 29972 13812
rect 29932 13734 29960 13806
rect 29920 13728 29972 13734
rect 29920 13670 29972 13676
rect 29932 13326 29960 13670
rect 30300 13462 30328 13942
rect 30564 13932 30616 13938
rect 30564 13874 30616 13880
rect 30840 13932 30892 13938
rect 30840 13874 30892 13880
rect 30576 13462 30604 13874
rect 30852 13530 30880 13874
rect 30840 13524 30892 13530
rect 30840 13466 30892 13472
rect 30288 13456 30340 13462
rect 30288 13398 30340 13404
rect 30564 13456 30616 13462
rect 30564 13398 30616 13404
rect 30944 13394 30972 16934
rect 31760 15360 31812 15366
rect 31760 15302 31812 15308
rect 31576 14884 31628 14890
rect 31576 14826 31628 14832
rect 31392 14816 31444 14822
rect 31392 14758 31444 14764
rect 31404 14414 31432 14758
rect 31392 14408 31444 14414
rect 31392 14350 31444 14356
rect 31588 14074 31616 14826
rect 31576 14068 31628 14074
rect 31576 14010 31628 14016
rect 31772 13954 31800 15302
rect 32232 15094 32260 16934
rect 34796 16788 34848 16794
rect 34796 16730 34848 16736
rect 33790 16348 34098 16357
rect 33790 16346 33796 16348
rect 33852 16346 33876 16348
rect 33932 16346 33956 16348
rect 34012 16346 34036 16348
rect 34092 16346 34098 16348
rect 33852 16294 33854 16346
rect 34034 16294 34036 16346
rect 33790 16292 33796 16294
rect 33852 16292 33876 16294
rect 33932 16292 33956 16294
rect 34012 16292 34036 16294
rect 34092 16292 34098 16294
rect 33790 16283 34098 16292
rect 32956 15700 33008 15706
rect 32956 15642 33008 15648
rect 32680 15428 32732 15434
rect 32680 15370 32732 15376
rect 32496 15360 32548 15366
rect 32496 15302 32548 15308
rect 32220 15088 32272 15094
rect 32220 15030 32272 15036
rect 31852 14952 31904 14958
rect 31852 14894 31904 14900
rect 31496 13938 31800 13954
rect 31496 13932 31812 13938
rect 31496 13926 31760 13932
rect 31496 13462 31524 13926
rect 31760 13874 31812 13880
rect 31760 13796 31812 13802
rect 31760 13738 31812 13744
rect 31772 13462 31800 13738
rect 31484 13456 31536 13462
rect 31484 13398 31536 13404
rect 31760 13456 31812 13462
rect 31760 13398 31812 13404
rect 30932 13388 30984 13394
rect 30932 13330 30984 13336
rect 29920 13320 29972 13326
rect 29920 13262 29972 13268
rect 30564 13320 30616 13326
rect 30564 13262 30616 13268
rect 29184 12844 29236 12850
rect 29184 12786 29236 12792
rect 29460 12844 29512 12850
rect 29460 12786 29512 12792
rect 28908 12300 28960 12306
rect 28908 12242 28960 12248
rect 28317 11452 28625 11461
rect 28317 11450 28323 11452
rect 28379 11450 28403 11452
rect 28459 11450 28483 11452
rect 28539 11450 28563 11452
rect 28619 11450 28625 11452
rect 28379 11398 28381 11450
rect 28561 11398 28563 11450
rect 28317 11396 28323 11398
rect 28379 11396 28403 11398
rect 28459 11396 28483 11398
rect 28539 11396 28563 11398
rect 28619 11396 28625 11398
rect 28317 11387 28625 11396
rect 28920 11286 28948 12242
rect 28908 11280 28960 11286
rect 28908 11222 28960 11228
rect 29196 11150 29224 12786
rect 29472 11898 29500 12786
rect 30576 12646 30604 13262
rect 30932 13252 30984 13258
rect 30932 13194 30984 13200
rect 30564 12640 30616 12646
rect 30564 12582 30616 12588
rect 30576 12434 30604 12582
rect 30576 12406 30696 12434
rect 29552 12368 29604 12374
rect 29552 12310 29604 12316
rect 29460 11892 29512 11898
rect 29460 11834 29512 11840
rect 29564 11762 29592 12310
rect 29736 12232 29788 12238
rect 29736 12174 29788 12180
rect 29644 12164 29696 12170
rect 29644 12106 29696 12112
rect 29552 11756 29604 11762
rect 29552 11698 29604 11704
rect 29656 11694 29684 12106
rect 29748 11898 29776 12174
rect 29736 11892 29788 11898
rect 29736 11834 29788 11840
rect 30668 11830 30696 12406
rect 30944 12170 30972 13194
rect 31496 12918 31524 13398
rect 31864 13258 31892 14894
rect 32232 14822 32260 15030
rect 32508 15026 32536 15302
rect 32496 15020 32548 15026
rect 32496 14962 32548 14968
rect 32692 14958 32720 15370
rect 32968 14958 32996 15642
rect 33790 15260 34098 15269
rect 33790 15258 33796 15260
rect 33852 15258 33876 15260
rect 33932 15258 33956 15260
rect 34012 15258 34036 15260
rect 34092 15258 34098 15260
rect 33852 15206 33854 15258
rect 34034 15206 34036 15258
rect 33790 15204 33796 15206
rect 33852 15204 33876 15206
rect 33932 15204 33956 15206
rect 34012 15204 34036 15206
rect 34092 15204 34098 15206
rect 33790 15195 34098 15204
rect 33508 15088 33560 15094
rect 33508 15030 33560 15036
rect 33968 15088 34020 15094
rect 33968 15030 34020 15036
rect 32312 14952 32364 14958
rect 32680 14952 32732 14958
rect 32312 14894 32364 14900
rect 32586 14920 32642 14929
rect 32220 14816 32272 14822
rect 32220 14758 32272 14764
rect 32324 14346 32352 14894
rect 32680 14894 32732 14900
rect 32956 14952 33008 14958
rect 32956 14894 33008 14900
rect 32586 14855 32588 14864
rect 32640 14855 32642 14864
rect 32588 14826 32640 14832
rect 32692 14618 32720 14894
rect 32772 14816 32824 14822
rect 32772 14758 32824 14764
rect 32680 14612 32732 14618
rect 32680 14554 32732 14560
rect 32312 14340 32364 14346
rect 32312 14282 32364 14288
rect 32692 14278 32720 14554
rect 32680 14272 32732 14278
rect 32680 14214 32732 14220
rect 32692 14006 32720 14214
rect 32680 14000 32732 14006
rect 32680 13942 32732 13948
rect 32680 13728 32732 13734
rect 32680 13670 32732 13676
rect 32128 13524 32180 13530
rect 32128 13466 32180 13472
rect 31852 13252 31904 13258
rect 31852 13194 31904 13200
rect 31944 12980 31996 12986
rect 31944 12922 31996 12928
rect 31484 12912 31536 12918
rect 31484 12854 31536 12860
rect 31574 12880 31630 12889
rect 31496 12458 31524 12854
rect 31574 12815 31576 12824
rect 31628 12815 31630 12824
rect 31576 12786 31628 12792
rect 31956 12646 31984 12922
rect 32140 12714 32168 13466
rect 32404 13456 32456 13462
rect 32404 13398 32456 13404
rect 32416 13258 32444 13398
rect 32692 13326 32720 13670
rect 32784 13326 32812 14758
rect 32968 14482 32996 14894
rect 33416 14816 33468 14822
rect 33416 14758 33468 14764
rect 32956 14476 33008 14482
rect 32956 14418 33008 14424
rect 32968 13938 32996 14418
rect 33232 14272 33284 14278
rect 33232 14214 33284 14220
rect 32956 13932 33008 13938
rect 32956 13874 33008 13880
rect 32680 13320 32732 13326
rect 32494 13288 32550 13297
rect 32404 13252 32456 13258
rect 32680 13262 32732 13268
rect 32772 13320 32824 13326
rect 32772 13262 32824 13268
rect 33140 13320 33192 13326
rect 33140 13262 33192 13268
rect 32494 13223 32496 13232
rect 32404 13194 32456 13200
rect 32548 13223 32550 13232
rect 32496 13194 32548 13200
rect 32508 12782 32536 13194
rect 32680 13184 32732 13190
rect 32680 13126 32732 13132
rect 32692 12850 32720 13126
rect 33048 12980 33100 12986
rect 33048 12922 33100 12928
rect 32588 12844 32640 12850
rect 32588 12786 32640 12792
rect 32680 12844 32732 12850
rect 32680 12786 32732 12792
rect 32496 12776 32548 12782
rect 32600 12753 32628 12786
rect 32496 12718 32548 12724
rect 32586 12744 32642 12753
rect 32128 12708 32180 12714
rect 32586 12679 32642 12688
rect 32128 12650 32180 12656
rect 31944 12640 31996 12646
rect 31944 12582 31996 12588
rect 31208 12436 31260 12442
rect 31496 12430 31800 12458
rect 31208 12378 31260 12384
rect 30932 12164 30984 12170
rect 30932 12106 30984 12112
rect 30656 11824 30708 11830
rect 30656 11766 30708 11772
rect 29644 11688 29696 11694
rect 29644 11630 29696 11636
rect 30288 11688 30340 11694
rect 30288 11630 30340 11636
rect 29644 11552 29696 11558
rect 29644 11494 29696 11500
rect 29656 11354 29684 11494
rect 29644 11348 29696 11354
rect 29644 11290 29696 11296
rect 30300 11150 30328 11630
rect 29184 11144 29236 11150
rect 29184 11086 29236 11092
rect 29736 11144 29788 11150
rect 29736 11086 29788 11092
rect 30288 11144 30340 11150
rect 30288 11086 30340 11092
rect 30656 11144 30708 11150
rect 30656 11086 30708 11092
rect 27620 10668 27672 10674
rect 27620 10610 27672 10616
rect 28724 10668 28776 10674
rect 28724 10610 28776 10616
rect 27632 9518 27660 10610
rect 28317 10364 28625 10373
rect 28317 10362 28323 10364
rect 28379 10362 28403 10364
rect 28459 10362 28483 10364
rect 28539 10362 28563 10364
rect 28619 10362 28625 10364
rect 28379 10310 28381 10362
rect 28561 10310 28563 10362
rect 28317 10308 28323 10310
rect 28379 10308 28403 10310
rect 28459 10308 28483 10310
rect 28539 10308 28563 10310
rect 28619 10308 28625 10310
rect 28317 10299 28625 10308
rect 27620 9512 27672 9518
rect 27620 9454 27672 9460
rect 28317 9276 28625 9285
rect 28317 9274 28323 9276
rect 28379 9274 28403 9276
rect 28459 9274 28483 9276
rect 28539 9274 28563 9276
rect 28619 9274 28625 9276
rect 28379 9222 28381 9274
rect 28561 9222 28563 9274
rect 28317 9220 28323 9222
rect 28379 9220 28403 9222
rect 28459 9220 28483 9222
rect 28539 9220 28563 9222
rect 28619 9220 28625 9222
rect 28317 9211 28625 9220
rect 27528 9104 27580 9110
rect 27528 9046 27580 9052
rect 25780 9036 25832 9042
rect 25780 8978 25832 8984
rect 26608 9036 26660 9042
rect 26608 8978 26660 8984
rect 27344 9036 27396 9042
rect 27344 8978 27396 8984
rect 25688 8900 25740 8906
rect 25688 8842 25740 8848
rect 25596 8628 25648 8634
rect 25596 8570 25648 8576
rect 25700 8090 25728 8842
rect 25964 8832 26016 8838
rect 25964 8774 26016 8780
rect 25976 8634 26004 8774
rect 25964 8628 26016 8634
rect 25964 8570 26016 8576
rect 25688 8084 25740 8090
rect 25688 8026 25740 8032
rect 25976 7954 26004 8570
rect 26148 8424 26200 8430
rect 26148 8366 26200 8372
rect 25964 7948 26016 7954
rect 25964 7890 26016 7896
rect 25504 7880 25556 7886
rect 25504 7822 25556 7828
rect 25516 7410 25544 7822
rect 25504 7404 25556 7410
rect 25504 7346 25556 7352
rect 25596 7200 25648 7206
rect 25596 7142 25648 7148
rect 24032 6792 24084 6798
rect 24032 6734 24084 6740
rect 24584 6792 24636 6798
rect 24584 6734 24636 6740
rect 24044 6458 24072 6734
rect 24032 6452 24084 6458
rect 24032 6394 24084 6400
rect 24400 6180 24452 6186
rect 24400 6122 24452 6128
rect 24412 5914 24440 6122
rect 24400 5908 24452 5914
rect 24400 5850 24452 5856
rect 24412 5370 24440 5850
rect 24596 5778 24624 6734
rect 25608 6730 25636 7142
rect 25596 6724 25648 6730
rect 25596 6666 25648 6672
rect 25228 6656 25280 6662
rect 25228 6598 25280 6604
rect 25240 6458 25268 6598
rect 25228 6452 25280 6458
rect 25228 6394 25280 6400
rect 26160 6254 26188 8366
rect 25320 6248 25372 6254
rect 25318 6216 25320 6225
rect 26148 6248 26200 6254
rect 25372 6216 25374 6225
rect 26148 6190 26200 6196
rect 25318 6151 25374 6160
rect 26792 6180 26844 6186
rect 26792 6122 26844 6128
rect 26332 6112 26384 6118
rect 26332 6054 26384 6060
rect 24584 5772 24636 5778
rect 24584 5714 24636 5720
rect 24400 5364 24452 5370
rect 24400 5306 24452 5312
rect 24596 5302 24624 5714
rect 26344 5710 26372 6054
rect 26804 5778 26832 6122
rect 26792 5772 26844 5778
rect 26792 5714 26844 5720
rect 26332 5704 26384 5710
rect 26332 5646 26384 5652
rect 24584 5296 24636 5302
rect 24584 5238 24636 5244
rect 26804 4690 26832 5714
rect 27356 5030 27384 8978
rect 27710 8936 27766 8945
rect 27710 8871 27712 8880
rect 27764 8871 27766 8880
rect 27712 8842 27764 8848
rect 27620 8832 27672 8838
rect 27620 8774 27672 8780
rect 27632 8498 27660 8774
rect 28736 8566 28764 10610
rect 29748 10470 29776 11086
rect 30668 10810 30696 11086
rect 30944 11014 30972 12106
rect 31220 12102 31248 12378
rect 31772 12374 31800 12430
rect 31760 12368 31812 12374
rect 31760 12310 31812 12316
rect 31956 12238 31984 12582
rect 32140 12306 32168 12650
rect 32128 12300 32180 12306
rect 32128 12242 32180 12248
rect 32496 12300 32548 12306
rect 32496 12242 32548 12248
rect 31760 12232 31812 12238
rect 31760 12174 31812 12180
rect 31944 12232 31996 12238
rect 31944 12174 31996 12180
rect 31208 12096 31260 12102
rect 31208 12038 31260 12044
rect 31220 11830 31248 12038
rect 31208 11824 31260 11830
rect 31208 11766 31260 11772
rect 31772 11694 31800 12174
rect 31956 11762 31984 12174
rect 32128 12164 32180 12170
rect 32128 12106 32180 12112
rect 32140 11830 32168 12106
rect 32128 11824 32180 11830
rect 32128 11766 32180 11772
rect 31852 11756 31904 11762
rect 31852 11698 31904 11704
rect 31944 11756 31996 11762
rect 31944 11698 31996 11704
rect 31760 11688 31812 11694
rect 31760 11630 31812 11636
rect 31760 11552 31812 11558
rect 31760 11494 31812 11500
rect 30932 11008 30984 11014
rect 30932 10950 30984 10956
rect 30944 10810 30972 10950
rect 30656 10804 30708 10810
rect 30656 10746 30708 10752
rect 30932 10804 30984 10810
rect 30932 10746 30984 10752
rect 31300 10668 31352 10674
rect 31300 10610 31352 10616
rect 29736 10464 29788 10470
rect 29736 10406 29788 10412
rect 29748 10062 29776 10406
rect 29000 10056 29052 10062
rect 29000 9998 29052 10004
rect 29736 10056 29788 10062
rect 29828 10056 29880 10062
rect 29736 9998 29788 10004
rect 29826 10024 29828 10033
rect 30932 10056 30984 10062
rect 29880 10024 29882 10033
rect 29012 9654 29040 9998
rect 30932 9998 30984 10004
rect 29826 9959 29882 9968
rect 30656 9920 30708 9926
rect 30656 9862 30708 9868
rect 30668 9654 30696 9862
rect 29000 9648 29052 9654
rect 29000 9590 29052 9596
rect 29184 9648 29236 9654
rect 29184 9590 29236 9596
rect 30656 9648 30708 9654
rect 30656 9590 30708 9596
rect 29196 9110 29224 9590
rect 29828 9376 29880 9382
rect 29828 9318 29880 9324
rect 29840 9110 29868 9318
rect 29184 9104 29236 9110
rect 29184 9046 29236 9052
rect 29828 9104 29880 9110
rect 29828 9046 29880 9052
rect 30668 9042 30696 9590
rect 30944 9450 30972 9998
rect 31312 9722 31340 10610
rect 31772 10062 31800 11494
rect 31864 11354 31892 11698
rect 31852 11348 31904 11354
rect 31852 11290 31904 11296
rect 32508 11150 32536 12242
rect 32600 11150 32628 12679
rect 33060 12374 33088 12922
rect 33048 12368 33100 12374
rect 33048 12310 33100 12316
rect 32772 12164 32824 12170
rect 32772 12106 32824 12112
rect 32784 11830 32812 12106
rect 33152 12102 33180 13262
rect 33244 12918 33272 14214
rect 33428 13938 33456 14758
rect 33520 14414 33548 15030
rect 33600 15020 33652 15026
rect 33600 14962 33652 14968
rect 33612 14618 33640 14962
rect 33980 14929 34008 15030
rect 33966 14920 34022 14929
rect 33966 14855 34022 14864
rect 34520 14884 34572 14890
rect 34520 14826 34572 14832
rect 33600 14612 33652 14618
rect 33600 14554 33652 14560
rect 33508 14408 33560 14414
rect 33508 14350 33560 14356
rect 33520 14074 33548 14350
rect 33790 14172 34098 14181
rect 33790 14170 33796 14172
rect 33852 14170 33876 14172
rect 33932 14170 33956 14172
rect 34012 14170 34036 14172
rect 34092 14170 34098 14172
rect 33852 14118 33854 14170
rect 34034 14118 34036 14170
rect 33790 14116 33796 14118
rect 33852 14116 33876 14118
rect 33932 14116 33956 14118
rect 34012 14116 34036 14118
rect 34092 14116 34098 14118
rect 33790 14107 34098 14116
rect 33508 14068 33560 14074
rect 33508 14010 33560 14016
rect 33692 14000 33744 14006
rect 33692 13942 33744 13948
rect 33416 13932 33468 13938
rect 33416 13874 33468 13880
rect 33416 13524 33468 13530
rect 33416 13466 33468 13472
rect 33428 12918 33456 13466
rect 33232 12912 33284 12918
rect 33232 12854 33284 12860
rect 33416 12912 33468 12918
rect 33416 12854 33468 12860
rect 33506 12880 33562 12889
rect 33506 12815 33562 12824
rect 33520 12714 33548 12815
rect 33508 12708 33560 12714
rect 33508 12650 33560 12656
rect 33324 12436 33376 12442
rect 33324 12378 33376 12384
rect 33232 12232 33284 12238
rect 33232 12174 33284 12180
rect 33140 12096 33192 12102
rect 33140 12038 33192 12044
rect 32772 11824 32824 11830
rect 32772 11766 32824 11772
rect 32784 11558 32812 11766
rect 32772 11552 32824 11558
rect 32772 11494 32824 11500
rect 33152 11218 33180 12038
rect 33244 11354 33272 12174
rect 33336 11558 33364 12378
rect 33520 11898 33548 12650
rect 33508 11892 33560 11898
rect 33508 11834 33560 11840
rect 33704 11694 33732 13942
rect 33790 13084 34098 13093
rect 33790 13082 33796 13084
rect 33852 13082 33876 13084
rect 33932 13082 33956 13084
rect 34012 13082 34036 13084
rect 34092 13082 34098 13084
rect 33852 13030 33854 13082
rect 34034 13030 34036 13082
rect 33790 13028 33796 13030
rect 33852 13028 33876 13030
rect 33932 13028 33956 13030
rect 34012 13028 34036 13030
rect 34092 13028 34098 13030
rect 33790 13019 34098 13028
rect 34532 12434 34560 14826
rect 34808 14074 34836 16730
rect 34900 15162 34928 16934
rect 34888 15156 34940 15162
rect 34888 15098 34940 15104
rect 37832 15088 37884 15094
rect 37832 15030 37884 15036
rect 36544 15020 36596 15026
rect 36544 14962 36596 14968
rect 36912 15020 36964 15026
rect 36912 14962 36964 14968
rect 34888 14816 34940 14822
rect 34888 14758 34940 14764
rect 34900 14414 34928 14758
rect 36452 14544 36504 14550
rect 36452 14486 36504 14492
rect 34888 14408 34940 14414
rect 34888 14350 34940 14356
rect 35164 14408 35216 14414
rect 35164 14350 35216 14356
rect 34796 14068 34848 14074
rect 34796 14010 34848 14016
rect 34808 13938 34836 14010
rect 34796 13932 34848 13938
rect 34796 13874 34848 13880
rect 34532 12406 34744 12434
rect 33790 11996 34098 12005
rect 33790 11994 33796 11996
rect 33852 11994 33876 11996
rect 33932 11994 33956 11996
rect 34012 11994 34036 11996
rect 34092 11994 34098 11996
rect 33852 11942 33854 11994
rect 34034 11942 34036 11994
rect 33790 11940 33796 11942
rect 33852 11940 33876 11942
rect 33932 11940 33956 11942
rect 34012 11940 34036 11942
rect 34092 11940 34098 11942
rect 33790 11931 34098 11940
rect 33508 11688 33560 11694
rect 33508 11630 33560 11636
rect 33692 11688 33744 11694
rect 33692 11630 33744 11636
rect 33324 11552 33376 11558
rect 33324 11494 33376 11500
rect 33232 11348 33284 11354
rect 33232 11290 33284 11296
rect 33140 11212 33192 11218
rect 33140 11154 33192 11160
rect 32496 11144 32548 11150
rect 32496 11086 32548 11092
rect 32588 11144 32640 11150
rect 32588 11086 32640 11092
rect 32680 11144 32732 11150
rect 32680 11086 32732 11092
rect 32404 11076 32456 11082
rect 32404 11018 32456 11024
rect 32416 10810 32444 11018
rect 32692 11014 32720 11086
rect 32680 11008 32732 11014
rect 32680 10950 32732 10956
rect 32404 10804 32456 10810
rect 32404 10746 32456 10752
rect 31852 10124 31904 10130
rect 31852 10066 31904 10072
rect 31760 10056 31812 10062
rect 31760 9998 31812 10004
rect 31300 9716 31352 9722
rect 31300 9658 31352 9664
rect 30932 9444 30984 9450
rect 30932 9386 30984 9392
rect 31668 9376 31720 9382
rect 31668 9318 31720 9324
rect 30656 9036 30708 9042
rect 30656 8978 30708 8984
rect 29000 8968 29052 8974
rect 29000 8910 29052 8916
rect 31576 8968 31628 8974
rect 31576 8910 31628 8916
rect 28908 8900 28960 8906
rect 28908 8842 28960 8848
rect 28724 8560 28776 8566
rect 28724 8502 28776 8508
rect 27620 8492 27672 8498
rect 27620 8434 27672 8440
rect 28172 8288 28224 8294
rect 28172 8230 28224 8236
rect 27618 7984 27674 7993
rect 27618 7919 27620 7928
rect 27672 7919 27674 7928
rect 27620 7890 27672 7896
rect 28184 7342 28212 8230
rect 28317 8188 28625 8197
rect 28317 8186 28323 8188
rect 28379 8186 28403 8188
rect 28459 8186 28483 8188
rect 28539 8186 28563 8188
rect 28619 8186 28625 8188
rect 28379 8134 28381 8186
rect 28561 8134 28563 8186
rect 28317 8132 28323 8134
rect 28379 8132 28403 8134
rect 28459 8132 28483 8134
rect 28539 8132 28563 8134
rect 28619 8132 28625 8134
rect 28317 8123 28625 8132
rect 28172 7336 28224 7342
rect 28172 7278 28224 7284
rect 27988 6656 28040 6662
rect 27988 6598 28040 6604
rect 28000 6390 28028 6598
rect 27988 6384 28040 6390
rect 27988 6326 28040 6332
rect 27896 6316 27948 6322
rect 27896 6258 27948 6264
rect 27908 5846 27936 6258
rect 27988 6248 28040 6254
rect 27988 6190 28040 6196
rect 27896 5840 27948 5846
rect 27896 5782 27948 5788
rect 28000 5778 28028 6190
rect 28184 6186 28212 7278
rect 28317 7100 28625 7109
rect 28317 7098 28323 7100
rect 28379 7098 28403 7100
rect 28459 7098 28483 7100
rect 28539 7098 28563 7100
rect 28619 7098 28625 7100
rect 28379 7046 28381 7098
rect 28561 7046 28563 7098
rect 28317 7044 28323 7046
rect 28379 7044 28403 7046
rect 28459 7044 28483 7046
rect 28539 7044 28563 7046
rect 28619 7044 28625 7046
rect 28317 7035 28625 7044
rect 28172 6180 28224 6186
rect 28172 6122 28224 6128
rect 27988 5772 28040 5778
rect 27988 5714 28040 5720
rect 27436 5704 27488 5710
rect 27436 5646 27488 5652
rect 27344 5024 27396 5030
rect 27344 4966 27396 4972
rect 26792 4684 26844 4690
rect 26792 4626 26844 4632
rect 23940 4208 23992 4214
rect 23940 4150 23992 4156
rect 23756 3936 23808 3942
rect 23756 3878 23808 3884
rect 23768 3670 23796 3878
rect 26884 3732 26936 3738
rect 26884 3674 26936 3680
rect 23756 3664 23808 3670
rect 23756 3606 23808 3612
rect 23388 3596 23440 3602
rect 23388 3538 23440 3544
rect 22843 3292 23151 3301
rect 22843 3290 22849 3292
rect 22905 3290 22929 3292
rect 22985 3290 23009 3292
rect 23065 3290 23089 3292
rect 23145 3290 23151 3292
rect 22905 3238 22907 3290
rect 23087 3238 23089 3290
rect 22843 3236 22849 3238
rect 22905 3236 22929 3238
rect 22985 3236 23009 3238
rect 23065 3236 23089 3238
rect 23145 3236 23151 3238
rect 22843 3227 23151 3236
rect 26896 3194 26924 3674
rect 26884 3188 26936 3194
rect 26884 3130 26936 3136
rect 18604 3052 18656 3058
rect 18604 2994 18656 3000
rect 18880 3052 18932 3058
rect 18880 2994 18932 3000
rect 22468 3052 22520 3058
rect 22468 2994 22520 3000
rect 22652 2848 22704 2854
rect 22652 2790 22704 2796
rect 17052 2746 17172 2774
rect 17144 2650 17172 2746
rect 17370 2748 17678 2757
rect 17370 2746 17376 2748
rect 17432 2746 17456 2748
rect 17512 2746 17536 2748
rect 17592 2746 17616 2748
rect 17672 2746 17678 2748
rect 17432 2694 17434 2746
rect 17614 2694 17616 2746
rect 17370 2692 17376 2694
rect 17432 2692 17456 2694
rect 17512 2692 17536 2694
rect 17592 2692 17616 2694
rect 17672 2692 17678 2694
rect 17370 2683 17678 2692
rect 17132 2644 17184 2650
rect 17132 2586 17184 2592
rect 22664 2446 22692 2790
rect 27356 2650 27384 4966
rect 27448 4010 27476 5646
rect 27804 4820 27856 4826
rect 27804 4762 27856 4768
rect 27816 4214 27844 4762
rect 27896 4548 27948 4554
rect 27896 4490 27948 4496
rect 27804 4208 27856 4214
rect 27804 4150 27856 4156
rect 27908 4146 27936 4490
rect 27896 4140 27948 4146
rect 27896 4082 27948 4088
rect 28000 4078 28028 5714
rect 28184 5370 28212 6122
rect 28317 6012 28625 6021
rect 28317 6010 28323 6012
rect 28379 6010 28403 6012
rect 28459 6010 28483 6012
rect 28539 6010 28563 6012
rect 28619 6010 28625 6012
rect 28379 5958 28381 6010
rect 28561 5958 28563 6010
rect 28317 5956 28323 5958
rect 28379 5956 28403 5958
rect 28459 5956 28483 5958
rect 28539 5956 28563 5958
rect 28619 5956 28625 5958
rect 28317 5947 28625 5956
rect 28264 5568 28316 5574
rect 28264 5510 28316 5516
rect 28172 5364 28224 5370
rect 28172 5306 28224 5312
rect 28276 5114 28304 5510
rect 28736 5302 28764 8502
rect 28920 8430 28948 8842
rect 28908 8424 28960 8430
rect 28908 8366 28960 8372
rect 29012 8022 29040 8910
rect 31484 8900 31536 8906
rect 31484 8842 31536 8848
rect 30196 8832 30248 8838
rect 30196 8774 30248 8780
rect 30288 8832 30340 8838
rect 30288 8774 30340 8780
rect 30208 8634 30236 8774
rect 30196 8628 30248 8634
rect 30196 8570 30248 8576
rect 29736 8492 29788 8498
rect 29736 8434 29788 8440
rect 30196 8492 30248 8498
rect 30196 8434 30248 8440
rect 29184 8288 29236 8294
rect 29184 8230 29236 8236
rect 29000 8016 29052 8022
rect 29000 7958 29052 7964
rect 29196 7886 29224 8230
rect 29748 8090 29776 8434
rect 29736 8084 29788 8090
rect 29736 8026 29788 8032
rect 30208 8022 30236 8434
rect 30196 8016 30248 8022
rect 30196 7958 30248 7964
rect 29184 7880 29236 7886
rect 29184 7822 29236 7828
rect 28816 7404 28868 7410
rect 28816 7346 28868 7352
rect 28828 7002 28856 7346
rect 30012 7200 30064 7206
rect 30012 7142 30064 7148
rect 28816 6996 28868 7002
rect 28816 6938 28868 6944
rect 30024 6798 30052 7142
rect 30012 6792 30064 6798
rect 30012 6734 30064 6740
rect 29736 6724 29788 6730
rect 29736 6666 29788 6672
rect 29748 5914 29776 6666
rect 30194 6352 30250 6361
rect 30194 6287 30250 6296
rect 30104 6112 30156 6118
rect 30104 6054 30156 6060
rect 29736 5908 29788 5914
rect 29736 5850 29788 5856
rect 30116 5710 30144 6054
rect 30104 5704 30156 5710
rect 30104 5646 30156 5652
rect 30208 5642 30236 6287
rect 30196 5636 30248 5642
rect 30196 5578 30248 5584
rect 28724 5296 28776 5302
rect 28724 5238 28776 5244
rect 28184 5086 28304 5114
rect 28184 4622 28212 5086
rect 28317 4924 28625 4933
rect 28317 4922 28323 4924
rect 28379 4922 28403 4924
rect 28459 4922 28483 4924
rect 28539 4922 28563 4924
rect 28619 4922 28625 4924
rect 28379 4870 28381 4922
rect 28561 4870 28563 4922
rect 28317 4868 28323 4870
rect 28379 4868 28403 4870
rect 28459 4868 28483 4870
rect 28539 4868 28563 4870
rect 28619 4868 28625 4870
rect 28317 4859 28625 4868
rect 28172 4616 28224 4622
rect 28172 4558 28224 4564
rect 27988 4072 28040 4078
rect 27988 4014 28040 4020
rect 27436 4004 27488 4010
rect 27436 3946 27488 3952
rect 28317 3836 28625 3845
rect 28317 3834 28323 3836
rect 28379 3834 28403 3836
rect 28459 3834 28483 3836
rect 28539 3834 28563 3836
rect 28619 3834 28625 3836
rect 28379 3782 28381 3834
rect 28561 3782 28563 3834
rect 28317 3780 28323 3782
rect 28379 3780 28403 3782
rect 28459 3780 28483 3782
rect 28539 3780 28563 3782
rect 28619 3780 28625 3782
rect 28317 3771 28625 3780
rect 28317 2748 28625 2757
rect 28317 2746 28323 2748
rect 28379 2746 28403 2748
rect 28459 2746 28483 2748
rect 28539 2746 28563 2748
rect 28619 2746 28625 2748
rect 28379 2694 28381 2746
rect 28561 2694 28563 2746
rect 28317 2692 28323 2694
rect 28379 2692 28403 2694
rect 28459 2692 28483 2694
rect 28539 2692 28563 2694
rect 28619 2692 28625 2694
rect 28317 2683 28625 2692
rect 27344 2644 27396 2650
rect 27344 2586 27396 2592
rect 30208 2582 30236 5578
rect 30300 3398 30328 8774
rect 31496 8634 31524 8842
rect 31484 8628 31536 8634
rect 31484 8570 31536 8576
rect 31588 8498 31616 8910
rect 31680 8498 31708 9318
rect 31576 8492 31628 8498
rect 31576 8434 31628 8440
rect 31668 8492 31720 8498
rect 31668 8434 31720 8440
rect 31024 7880 31076 7886
rect 31024 7822 31076 7828
rect 30748 7540 30800 7546
rect 30748 7482 30800 7488
rect 30472 7336 30524 7342
rect 30472 7278 30524 7284
rect 30484 5778 30512 7278
rect 30760 6798 30788 7482
rect 30748 6792 30800 6798
rect 30748 6734 30800 6740
rect 30472 5772 30524 5778
rect 30472 5714 30524 5720
rect 31036 3942 31064 7822
rect 31208 7336 31260 7342
rect 31208 7278 31260 7284
rect 31220 5370 31248 7278
rect 31208 5364 31260 5370
rect 31208 5306 31260 5312
rect 31220 4690 31248 5306
rect 31484 5024 31536 5030
rect 31484 4966 31536 4972
rect 31496 4690 31524 4966
rect 31208 4684 31260 4690
rect 31208 4626 31260 4632
rect 31484 4684 31536 4690
rect 31484 4626 31536 4632
rect 31220 4570 31248 4626
rect 31128 4542 31248 4570
rect 31024 3936 31076 3942
rect 31024 3878 31076 3884
rect 31128 3534 31156 4542
rect 31668 3936 31720 3942
rect 31668 3878 31720 3884
rect 31116 3528 31168 3534
rect 31116 3470 31168 3476
rect 31680 3466 31708 3878
rect 31668 3460 31720 3466
rect 31668 3402 31720 3408
rect 30288 3392 30340 3398
rect 30288 3334 30340 3340
rect 30196 2576 30248 2582
rect 30196 2518 30248 2524
rect 16120 2440 16172 2446
rect 16120 2382 16172 2388
rect 16764 2440 16816 2446
rect 16764 2382 16816 2388
rect 17408 2440 17460 2446
rect 17408 2382 17460 2388
rect 19340 2440 19392 2446
rect 19340 2382 19392 2388
rect 20720 2440 20772 2446
rect 20720 2382 20772 2388
rect 22652 2440 22704 2446
rect 22652 2382 22704 2388
rect 23848 2440 23900 2446
rect 23848 2382 23900 2388
rect 25780 2440 25832 2446
rect 25780 2382 25832 2388
rect 27068 2440 27120 2446
rect 27068 2382 27120 2388
rect 29000 2440 29052 2446
rect 29000 2382 29052 2388
rect 30380 2440 30432 2446
rect 30380 2382 30432 2388
rect 16132 800 16160 2382
rect 17420 800 17448 2382
rect 19352 800 19380 2382
rect 20732 898 20760 2382
rect 22560 2304 22612 2310
rect 22560 2246 22612 2252
rect 20640 870 20760 898
rect 20640 800 20668 870
rect 22572 800 22600 2246
rect 22843 2204 23151 2213
rect 22843 2202 22849 2204
rect 22905 2202 22929 2204
rect 22985 2202 23009 2204
rect 23065 2202 23089 2204
rect 23145 2202 23151 2204
rect 22905 2150 22907 2202
rect 23087 2150 23089 2202
rect 22843 2148 22849 2150
rect 22905 2148 22929 2150
rect 22985 2148 23009 2150
rect 23065 2148 23089 2150
rect 23145 2148 23151 2150
rect 22843 2139 23151 2148
rect 23860 800 23888 2382
rect 25792 800 25820 2382
rect 27080 800 27108 2382
rect 29012 800 29040 2382
rect 30392 898 30420 2382
rect 31864 2310 31892 10066
rect 32692 10062 32720 10950
rect 32864 10532 32916 10538
rect 32864 10474 32916 10480
rect 32680 10056 32732 10062
rect 32680 9998 32732 10004
rect 32772 10056 32824 10062
rect 32772 9998 32824 10004
rect 32496 9920 32548 9926
rect 32496 9862 32548 9868
rect 32508 9586 32536 9862
rect 32784 9654 32812 9998
rect 32772 9648 32824 9654
rect 32772 9590 32824 9596
rect 32496 9580 32548 9586
rect 32496 9522 32548 9528
rect 32680 9104 32732 9110
rect 32680 9046 32732 9052
rect 32876 9058 32904 10474
rect 33520 10470 33548 11630
rect 33790 10908 34098 10917
rect 33790 10906 33796 10908
rect 33852 10906 33876 10908
rect 33932 10906 33956 10908
rect 34012 10906 34036 10908
rect 34092 10906 34098 10908
rect 33852 10854 33854 10906
rect 34034 10854 34036 10906
rect 33790 10852 33796 10854
rect 33852 10852 33876 10854
rect 33932 10852 33956 10854
rect 34012 10852 34036 10854
rect 34092 10852 34098 10854
rect 33790 10843 34098 10852
rect 33508 10464 33560 10470
rect 33508 10406 33560 10412
rect 33520 9654 33548 10406
rect 33790 9820 34098 9829
rect 33790 9818 33796 9820
rect 33852 9818 33876 9820
rect 33932 9818 33956 9820
rect 34012 9818 34036 9820
rect 34092 9818 34098 9820
rect 33852 9766 33854 9818
rect 34034 9766 34036 9818
rect 33790 9764 33796 9766
rect 33852 9764 33876 9766
rect 33932 9764 33956 9766
rect 34012 9764 34036 9766
rect 34092 9764 34098 9766
rect 33790 9755 34098 9764
rect 33508 9648 33560 9654
rect 33508 9590 33560 9596
rect 33692 9648 33744 9654
rect 33692 9590 33744 9596
rect 32956 9376 33008 9382
rect 32956 9318 33008 9324
rect 32968 9178 32996 9318
rect 33704 9178 33732 9590
rect 34336 9376 34388 9382
rect 34336 9318 34388 9324
rect 32956 9172 33008 9178
rect 32956 9114 33008 9120
rect 33692 9172 33744 9178
rect 33692 9114 33744 9120
rect 34152 9172 34204 9178
rect 34152 9114 34204 9120
rect 31944 8832 31996 8838
rect 31944 8774 31996 8780
rect 31956 6254 31984 8774
rect 32496 8560 32548 8566
rect 32496 8502 32548 8508
rect 32404 7744 32456 7750
rect 32404 7686 32456 7692
rect 32416 7478 32444 7686
rect 32404 7472 32456 7478
rect 32404 7414 32456 7420
rect 32508 6882 32536 8502
rect 32588 7880 32640 7886
rect 32588 7822 32640 7828
rect 32600 7002 32628 7822
rect 32692 7478 32720 9046
rect 32876 9030 32996 9058
rect 32968 8974 32996 9030
rect 32956 8968 33008 8974
rect 32956 8910 33008 8916
rect 32968 7954 32996 8910
rect 34164 8906 34192 9114
rect 34348 8974 34376 9318
rect 34520 9036 34572 9042
rect 34520 8978 34572 8984
rect 34336 8968 34388 8974
rect 34336 8910 34388 8916
rect 34152 8900 34204 8906
rect 34152 8842 34204 8848
rect 33790 8732 34098 8741
rect 33790 8730 33796 8732
rect 33852 8730 33876 8732
rect 33932 8730 33956 8732
rect 34012 8730 34036 8732
rect 34092 8730 34098 8732
rect 33852 8678 33854 8730
rect 34034 8678 34036 8730
rect 33790 8676 33796 8678
rect 33852 8676 33876 8678
rect 33932 8676 33956 8678
rect 34012 8676 34036 8678
rect 34092 8676 34098 8678
rect 33790 8667 34098 8676
rect 34532 8634 34560 8978
rect 34612 8968 34664 8974
rect 34612 8910 34664 8916
rect 34520 8628 34572 8634
rect 34520 8570 34572 8576
rect 34624 8498 34652 8910
rect 34520 8492 34572 8498
rect 34520 8434 34572 8440
rect 34612 8492 34664 8498
rect 34612 8434 34664 8440
rect 34532 8090 34560 8434
rect 34520 8084 34572 8090
rect 34520 8026 34572 8032
rect 32956 7948 33008 7954
rect 32956 7890 33008 7896
rect 33790 7644 34098 7653
rect 33790 7642 33796 7644
rect 33852 7642 33876 7644
rect 33932 7642 33956 7644
rect 34012 7642 34036 7644
rect 34092 7642 34098 7644
rect 33852 7590 33854 7642
rect 34034 7590 34036 7642
rect 33790 7588 33796 7590
rect 33852 7588 33876 7590
rect 33932 7588 33956 7590
rect 34012 7588 34036 7590
rect 34092 7588 34098 7590
rect 33790 7579 34098 7588
rect 32680 7472 32732 7478
rect 32680 7414 32732 7420
rect 32588 6996 32640 7002
rect 32588 6938 32640 6944
rect 32508 6854 32628 6882
rect 32692 6866 32720 7414
rect 33508 7200 33560 7206
rect 33508 7142 33560 7148
rect 32600 6730 32628 6854
rect 32680 6860 32732 6866
rect 32680 6802 32732 6808
rect 33048 6860 33100 6866
rect 33048 6802 33100 6808
rect 32588 6724 32640 6730
rect 32588 6666 32640 6672
rect 32220 6316 32272 6322
rect 32220 6258 32272 6264
rect 31944 6248 31996 6254
rect 31944 6190 31996 6196
rect 31956 5914 31984 6190
rect 32036 6112 32088 6118
rect 32036 6054 32088 6060
rect 31944 5908 31996 5914
rect 31944 5850 31996 5856
rect 32048 5710 32076 6054
rect 32232 5710 32260 6258
rect 32496 5908 32548 5914
rect 32496 5850 32548 5856
rect 31944 5704 31996 5710
rect 31944 5646 31996 5652
rect 32036 5704 32088 5710
rect 32036 5646 32088 5652
rect 32220 5704 32272 5710
rect 32220 5646 32272 5652
rect 31956 4010 31984 5646
rect 32128 5568 32180 5574
rect 32128 5510 32180 5516
rect 32140 5234 32168 5510
rect 32128 5228 32180 5234
rect 32128 5170 32180 5176
rect 32140 4593 32168 5170
rect 32232 5166 32260 5646
rect 32220 5160 32272 5166
rect 32220 5102 32272 5108
rect 32508 5098 32536 5850
rect 32496 5092 32548 5098
rect 32496 5034 32548 5040
rect 32126 4584 32182 4593
rect 32126 4519 32182 4528
rect 32140 4078 32168 4519
rect 32128 4072 32180 4078
rect 32128 4014 32180 4020
rect 31944 4004 31996 4010
rect 31944 3946 31996 3952
rect 32036 3936 32088 3942
rect 32036 3878 32088 3884
rect 32048 3738 32076 3878
rect 32036 3732 32088 3738
rect 32036 3674 32088 3680
rect 32600 2514 32628 6666
rect 32772 6656 32824 6662
rect 32772 6598 32824 6604
rect 32784 6474 32812 6598
rect 32784 6458 32904 6474
rect 32784 6452 32916 6458
rect 32784 6446 32864 6452
rect 32680 6112 32732 6118
rect 32680 6054 32732 6060
rect 32692 5234 32720 6054
rect 32784 5574 32812 6446
rect 32864 6394 32916 6400
rect 32954 6352 33010 6361
rect 33060 6322 33088 6802
rect 33520 6798 33548 7142
rect 34428 6860 34480 6866
rect 34428 6802 34480 6808
rect 33508 6792 33560 6798
rect 33692 6792 33744 6798
rect 33508 6734 33560 6740
rect 33612 6740 33692 6746
rect 33612 6734 33744 6740
rect 33140 6724 33192 6730
rect 33140 6666 33192 6672
rect 33612 6718 33732 6734
rect 33152 6322 33180 6666
rect 32954 6287 33010 6296
rect 33048 6316 33100 6322
rect 32864 6180 32916 6186
rect 32864 6122 32916 6128
rect 32772 5568 32824 5574
rect 32772 5510 32824 5516
rect 32876 5370 32904 6122
rect 32968 5710 32996 6287
rect 33048 6258 33100 6264
rect 33140 6316 33192 6322
rect 33140 6258 33192 6264
rect 33416 6316 33468 6322
rect 33416 6258 33468 6264
rect 32956 5704 33008 5710
rect 32956 5646 33008 5652
rect 32864 5364 32916 5370
rect 32864 5306 32916 5312
rect 32876 5234 32904 5306
rect 32680 5228 32732 5234
rect 32680 5170 32732 5176
rect 32864 5228 32916 5234
rect 32864 5170 32916 5176
rect 33152 4758 33180 6258
rect 33324 6180 33376 6186
rect 33324 6122 33376 6128
rect 33336 5234 33364 6122
rect 33428 5914 33456 6258
rect 33416 5908 33468 5914
rect 33416 5850 33468 5856
rect 33612 5846 33640 6718
rect 33692 6656 33744 6662
rect 33692 6598 33744 6604
rect 34152 6656 34204 6662
rect 34152 6598 34204 6604
rect 33704 5846 33732 6598
rect 33790 6556 34098 6565
rect 33790 6554 33796 6556
rect 33852 6554 33876 6556
rect 33932 6554 33956 6556
rect 34012 6554 34036 6556
rect 34092 6554 34098 6556
rect 33852 6502 33854 6554
rect 34034 6502 34036 6554
rect 33790 6500 33796 6502
rect 33852 6500 33876 6502
rect 33932 6500 33956 6502
rect 34012 6500 34036 6502
rect 34092 6500 34098 6502
rect 33790 6491 34098 6500
rect 34060 6316 34112 6322
rect 34060 6258 34112 6264
rect 33968 6248 34020 6254
rect 33968 6190 34020 6196
rect 33600 5840 33652 5846
rect 33600 5782 33652 5788
rect 33692 5840 33744 5846
rect 33692 5782 33744 5788
rect 33692 5704 33744 5710
rect 33692 5646 33744 5652
rect 33324 5228 33376 5234
rect 33324 5170 33376 5176
rect 33336 4758 33364 5170
rect 33704 4826 33732 5646
rect 33980 5574 34008 6190
rect 34072 5642 34100 6258
rect 34164 5914 34192 6598
rect 34336 6452 34388 6458
rect 34336 6394 34388 6400
rect 34242 6352 34298 6361
rect 34242 6287 34244 6296
rect 34296 6287 34298 6296
rect 34244 6258 34296 6264
rect 34348 6254 34376 6394
rect 34336 6248 34388 6254
rect 34336 6190 34388 6196
rect 34440 5914 34468 6802
rect 34152 5908 34204 5914
rect 34152 5850 34204 5856
rect 34428 5908 34480 5914
rect 34428 5850 34480 5856
rect 34060 5636 34112 5642
rect 34060 5578 34112 5584
rect 34152 5636 34204 5642
rect 34152 5578 34204 5584
rect 33968 5568 34020 5574
rect 33968 5510 34020 5516
rect 33790 5468 34098 5477
rect 33790 5466 33796 5468
rect 33852 5466 33876 5468
rect 33932 5466 33956 5468
rect 34012 5466 34036 5468
rect 34092 5466 34098 5468
rect 33852 5414 33854 5466
rect 34034 5414 34036 5466
rect 33790 5412 33796 5414
rect 33852 5412 33876 5414
rect 33932 5412 33956 5414
rect 34012 5412 34036 5414
rect 34092 5412 34098 5414
rect 33790 5403 34098 5412
rect 34164 5370 34192 5578
rect 34624 5370 34652 8434
rect 34716 7954 34744 12406
rect 35176 12102 35204 14350
rect 36360 14272 36412 14278
rect 36360 14214 36412 14220
rect 36268 14068 36320 14074
rect 36268 14010 36320 14016
rect 35440 13932 35492 13938
rect 35440 13874 35492 13880
rect 35348 12436 35400 12442
rect 35452 12434 35480 13874
rect 36084 13796 36136 13802
rect 36084 13738 36136 13744
rect 36096 13394 36124 13738
rect 36084 13388 36136 13394
rect 36084 13330 36136 13336
rect 36280 13326 36308 14010
rect 36372 14006 36400 14214
rect 36464 14074 36492 14486
rect 36556 14346 36584 14962
rect 36636 14816 36688 14822
rect 36636 14758 36688 14764
rect 36544 14340 36596 14346
rect 36544 14282 36596 14288
rect 36648 14074 36676 14758
rect 36820 14408 36872 14414
rect 36820 14350 36872 14356
rect 36452 14068 36504 14074
rect 36452 14010 36504 14016
rect 36636 14068 36688 14074
rect 36636 14010 36688 14016
rect 36360 14000 36412 14006
rect 36360 13942 36412 13948
rect 36464 13870 36492 14010
rect 36360 13864 36412 13870
rect 36360 13806 36412 13812
rect 36452 13864 36504 13870
rect 36452 13806 36504 13812
rect 36268 13320 36320 13326
rect 36268 13262 36320 13268
rect 35716 13252 35768 13258
rect 35716 13194 35768 13200
rect 35728 12850 35756 13194
rect 36372 13138 36400 13806
rect 36832 13802 36860 14350
rect 36924 14074 36952 14962
rect 37844 14822 37872 15030
rect 38948 14822 38976 16934
rect 39264 16892 39572 16901
rect 39264 16890 39270 16892
rect 39326 16890 39350 16892
rect 39406 16890 39430 16892
rect 39486 16890 39510 16892
rect 39566 16890 39572 16892
rect 39326 16838 39328 16890
rect 39508 16838 39510 16890
rect 39264 16836 39270 16838
rect 39326 16836 39350 16838
rect 39406 16836 39430 16838
rect 39486 16836 39510 16838
rect 39566 16836 39572 16838
rect 39264 16827 39572 16836
rect 40696 16454 40724 17138
rect 43732 16794 43760 17954
rect 43824 17202 43852 19200
rect 45006 19136 45062 19145
rect 45006 19071 45062 19080
rect 45020 18018 45048 19071
rect 45008 18012 45060 18018
rect 45008 17954 45060 17960
rect 44270 17776 44326 17785
rect 44270 17711 44326 17720
rect 44284 17338 44312 17711
rect 44737 17436 45045 17445
rect 44737 17434 44743 17436
rect 44799 17434 44823 17436
rect 44879 17434 44903 17436
rect 44959 17434 44983 17436
rect 45039 17434 45045 17436
rect 44799 17382 44801 17434
rect 44981 17382 44983 17434
rect 44737 17380 44743 17382
rect 44799 17380 44823 17382
rect 44879 17380 44903 17382
rect 44959 17380 44983 17382
rect 45039 17380 45045 17382
rect 44737 17371 45045 17380
rect 44272 17332 44324 17338
rect 44272 17274 44324 17280
rect 43812 17196 43864 17202
rect 43812 17138 43864 17144
rect 44088 17196 44140 17202
rect 44088 17138 44140 17144
rect 43720 16788 43772 16794
rect 43720 16730 43772 16736
rect 40684 16448 40736 16454
rect 40684 16390 40736 16396
rect 44100 16250 44128 17138
rect 45112 16794 45140 19200
rect 45100 16788 45152 16794
rect 45100 16730 45152 16736
rect 44737 16348 45045 16357
rect 44737 16346 44743 16348
rect 44799 16346 44823 16348
rect 44879 16346 44903 16348
rect 44959 16346 44983 16348
rect 45039 16346 45045 16348
rect 44799 16294 44801 16346
rect 44981 16294 44983 16346
rect 44737 16292 44743 16294
rect 44799 16292 44823 16294
rect 44879 16292 44903 16294
rect 44959 16292 44983 16294
rect 45039 16292 45045 16294
rect 44737 16283 45045 16292
rect 44088 16244 44140 16250
rect 44088 16186 44140 16192
rect 44364 15904 44416 15910
rect 44364 15846 44416 15852
rect 39264 15804 39572 15813
rect 39264 15802 39270 15804
rect 39326 15802 39350 15804
rect 39406 15802 39430 15804
rect 39486 15802 39510 15804
rect 39566 15802 39572 15804
rect 39326 15750 39328 15802
rect 39508 15750 39510 15802
rect 39264 15748 39270 15750
rect 39326 15748 39350 15750
rect 39406 15748 39430 15750
rect 39486 15748 39510 15750
rect 39566 15748 39572 15750
rect 39264 15739 39572 15748
rect 44376 15745 44404 15846
rect 44362 15736 44418 15745
rect 44362 15671 44418 15680
rect 44737 15260 45045 15269
rect 44737 15258 44743 15260
rect 44799 15258 44823 15260
rect 44879 15258 44903 15260
rect 44959 15258 44983 15260
rect 45039 15258 45045 15260
rect 44799 15206 44801 15258
rect 44981 15206 44983 15258
rect 44737 15204 44743 15206
rect 44799 15204 44823 15206
rect 44879 15204 44903 15206
rect 44959 15204 44983 15206
rect 45039 15204 45045 15206
rect 44737 15195 45045 15204
rect 37464 14816 37516 14822
rect 37464 14758 37516 14764
rect 37832 14816 37884 14822
rect 37832 14758 37884 14764
rect 38936 14816 38988 14822
rect 38936 14758 38988 14764
rect 37476 14414 37504 14758
rect 37464 14408 37516 14414
rect 37464 14350 37516 14356
rect 36912 14068 36964 14074
rect 36912 14010 36964 14016
rect 37280 14068 37332 14074
rect 37280 14010 37332 14016
rect 36820 13796 36872 13802
rect 36820 13738 36872 13744
rect 36636 13728 36688 13734
rect 36636 13670 36688 13676
rect 36004 13110 36400 13138
rect 36452 13184 36504 13190
rect 36452 13126 36504 13132
rect 35624 12844 35676 12850
rect 35624 12786 35676 12792
rect 35716 12844 35768 12850
rect 35716 12786 35768 12792
rect 35532 12436 35584 12442
rect 35452 12406 35532 12434
rect 35348 12378 35400 12384
rect 35636 12434 35664 12786
rect 35636 12406 35848 12434
rect 35532 12378 35584 12384
rect 35256 12368 35308 12374
rect 35256 12310 35308 12316
rect 35268 12170 35296 12310
rect 35256 12164 35308 12170
rect 35256 12106 35308 12112
rect 35164 12096 35216 12102
rect 35164 12038 35216 12044
rect 35360 12050 35388 12378
rect 35820 12374 35848 12406
rect 35808 12368 35860 12374
rect 35808 12310 35860 12316
rect 35716 12164 35768 12170
rect 35716 12106 35768 12112
rect 35624 12096 35676 12102
rect 35176 11150 35204 12038
rect 35360 12022 35480 12050
rect 35624 12038 35676 12044
rect 35452 11898 35480 12022
rect 35440 11892 35492 11898
rect 35440 11834 35492 11840
rect 35636 11830 35664 12038
rect 35728 11830 35756 12106
rect 35624 11824 35676 11830
rect 35624 11766 35676 11772
rect 35716 11824 35768 11830
rect 35716 11766 35768 11772
rect 35820 11762 35848 12310
rect 36004 12306 36032 13110
rect 36372 12918 36400 13110
rect 36176 12912 36228 12918
rect 36176 12854 36228 12860
rect 36360 12912 36412 12918
rect 36360 12854 36412 12860
rect 36084 12708 36136 12714
rect 36084 12650 36136 12656
rect 35992 12300 36044 12306
rect 35992 12242 36044 12248
rect 36096 11762 36124 12650
rect 36188 12238 36216 12854
rect 36464 12850 36492 13126
rect 36648 12850 36676 13670
rect 36832 13394 36860 13738
rect 37292 13530 37320 14010
rect 37648 14000 37700 14006
rect 37648 13942 37700 13948
rect 37556 13932 37608 13938
rect 37556 13874 37608 13880
rect 37464 13728 37516 13734
rect 37464 13670 37516 13676
rect 37280 13524 37332 13530
rect 37280 13466 37332 13472
rect 36820 13388 36872 13394
rect 36820 13330 36872 13336
rect 36268 12844 36320 12850
rect 36268 12786 36320 12792
rect 36452 12844 36504 12850
rect 36452 12786 36504 12792
rect 36636 12844 36688 12850
rect 36636 12786 36688 12792
rect 36280 12442 36308 12786
rect 36268 12436 36320 12442
rect 36268 12378 36320 12384
rect 36176 12232 36228 12238
rect 36176 12174 36228 12180
rect 36636 12232 36688 12238
rect 36636 12174 36688 12180
rect 36648 11898 36676 12174
rect 36544 11892 36596 11898
rect 36544 11834 36596 11840
rect 36636 11892 36688 11898
rect 36636 11834 36688 11840
rect 35256 11756 35308 11762
rect 35256 11698 35308 11704
rect 35808 11756 35860 11762
rect 35808 11698 35860 11704
rect 36084 11756 36136 11762
rect 36084 11698 36136 11704
rect 35268 11354 35296 11698
rect 35992 11688 36044 11694
rect 35992 11630 36044 11636
rect 35900 11552 35952 11558
rect 35900 11494 35952 11500
rect 35256 11348 35308 11354
rect 35256 11290 35308 11296
rect 35912 11218 35940 11494
rect 35900 11212 35952 11218
rect 35900 11154 35952 11160
rect 36004 11150 36032 11630
rect 36556 11626 36584 11834
rect 36636 11756 36688 11762
rect 36636 11698 36688 11704
rect 36544 11620 36596 11626
rect 36544 11562 36596 11568
rect 36452 11280 36504 11286
rect 36452 11222 36504 11228
rect 34980 11144 35032 11150
rect 35164 11144 35216 11150
rect 35032 11104 35164 11132
rect 34980 11086 35032 11092
rect 35164 11086 35216 11092
rect 35992 11144 36044 11150
rect 35992 11086 36044 11092
rect 36004 10674 36032 11086
rect 36464 11082 36492 11222
rect 36556 11150 36584 11562
rect 36544 11144 36596 11150
rect 36544 11086 36596 11092
rect 36648 11082 36676 11698
rect 36728 11552 36780 11558
rect 36728 11494 36780 11500
rect 36740 11354 36768 11494
rect 36728 11348 36780 11354
rect 36728 11290 36780 11296
rect 36452 11076 36504 11082
rect 36452 11018 36504 11024
rect 36636 11076 36688 11082
rect 36636 11018 36688 11024
rect 36360 11008 36412 11014
rect 36360 10950 36412 10956
rect 35992 10668 36044 10674
rect 35992 10610 36044 10616
rect 36372 10470 36400 10950
rect 36464 10810 36492 11018
rect 36452 10804 36504 10810
rect 36452 10746 36504 10752
rect 36832 10674 36860 13330
rect 37292 12238 37320 13466
rect 37476 13326 37504 13670
rect 37464 13320 37516 13326
rect 37464 13262 37516 13268
rect 37568 12986 37596 13874
rect 37556 12980 37608 12986
rect 37556 12922 37608 12928
rect 37660 12850 37688 13942
rect 37648 12844 37700 12850
rect 37648 12786 37700 12792
rect 37372 12640 37424 12646
rect 37372 12582 37424 12588
rect 37384 12238 37412 12582
rect 37280 12232 37332 12238
rect 37280 12174 37332 12180
rect 37372 12232 37424 12238
rect 37372 12174 37424 12180
rect 37660 11898 37688 12786
rect 37740 12164 37792 12170
rect 37740 12106 37792 12112
rect 37556 11892 37608 11898
rect 37556 11834 37608 11840
rect 37648 11892 37700 11898
rect 37648 11834 37700 11840
rect 37568 11694 37596 11834
rect 37752 11830 37780 12106
rect 37740 11824 37792 11830
rect 37740 11766 37792 11772
rect 37556 11688 37608 11694
rect 37556 11630 37608 11636
rect 37648 11620 37700 11626
rect 37648 11562 37700 11568
rect 37556 11552 37608 11558
rect 37556 11494 37608 11500
rect 37568 10674 37596 11494
rect 37660 11150 37688 11562
rect 37648 11144 37700 11150
rect 37648 11086 37700 11092
rect 36820 10668 36872 10674
rect 36820 10610 36872 10616
rect 37556 10668 37608 10674
rect 37556 10610 37608 10616
rect 36268 10464 36320 10470
rect 36268 10406 36320 10412
rect 36360 10464 36412 10470
rect 36360 10406 36412 10412
rect 36280 10130 36308 10406
rect 36832 10130 36860 10610
rect 36912 10464 36964 10470
rect 36912 10406 36964 10412
rect 36268 10124 36320 10130
rect 36268 10066 36320 10072
rect 36820 10124 36872 10130
rect 36820 10066 36872 10072
rect 36728 9988 36780 9994
rect 36728 9930 36780 9936
rect 36740 9722 36768 9930
rect 36728 9716 36780 9722
rect 36728 9658 36780 9664
rect 36924 9586 36952 10406
rect 36360 9580 36412 9586
rect 36360 9522 36412 9528
rect 36912 9580 36964 9586
rect 36912 9522 36964 9528
rect 37740 9580 37792 9586
rect 37740 9522 37792 9528
rect 34980 9512 35032 9518
rect 34980 9454 35032 9460
rect 34992 8838 35020 9454
rect 35716 9444 35768 9450
rect 35716 9386 35768 9392
rect 35728 9178 35756 9386
rect 36372 9178 36400 9522
rect 37556 9376 37608 9382
rect 37556 9318 37608 9324
rect 35716 9172 35768 9178
rect 35716 9114 35768 9120
rect 36360 9172 36412 9178
rect 36360 9114 36412 9120
rect 34980 8832 35032 8838
rect 34980 8774 35032 8780
rect 35728 8430 35756 9114
rect 35716 8424 35768 8430
rect 35716 8366 35768 8372
rect 35624 8356 35676 8362
rect 35624 8298 35676 8304
rect 34704 7948 34756 7954
rect 34704 7890 34756 7896
rect 35636 7886 35664 8298
rect 35728 7954 35756 8366
rect 35716 7948 35768 7954
rect 35716 7890 35768 7896
rect 35624 7880 35676 7886
rect 35624 7822 35676 7828
rect 35532 7744 35584 7750
rect 35532 7686 35584 7692
rect 35544 7410 35572 7686
rect 35636 7410 35664 7822
rect 35532 7404 35584 7410
rect 35532 7346 35584 7352
rect 35624 7404 35676 7410
rect 35624 7346 35676 7352
rect 36084 7404 36136 7410
rect 36084 7346 36136 7352
rect 35440 7336 35492 7342
rect 35440 7278 35492 7284
rect 35256 7200 35308 7206
rect 35256 7142 35308 7148
rect 35268 6798 35296 7142
rect 35452 6798 35480 7278
rect 35636 6866 35664 7346
rect 35900 7336 35952 7342
rect 35900 7278 35952 7284
rect 35624 6860 35676 6866
rect 35624 6802 35676 6808
rect 35912 6798 35940 7278
rect 35256 6792 35308 6798
rect 35256 6734 35308 6740
rect 35440 6792 35492 6798
rect 35440 6734 35492 6740
rect 35900 6792 35952 6798
rect 35900 6734 35952 6740
rect 34980 6656 35032 6662
rect 34980 6598 35032 6604
rect 34992 6322 35020 6598
rect 35452 6458 35480 6734
rect 36096 6730 36124 7346
rect 36372 7342 36400 9114
rect 37568 8974 37596 9318
rect 37464 8968 37516 8974
rect 37464 8910 37516 8916
rect 37556 8968 37608 8974
rect 37556 8910 37608 8916
rect 36360 7336 36412 7342
rect 36360 7278 36412 7284
rect 36268 7200 36320 7206
rect 36268 7142 36320 7148
rect 36084 6724 36136 6730
rect 36084 6666 36136 6672
rect 35440 6452 35492 6458
rect 35440 6394 35492 6400
rect 36280 6390 36308 7142
rect 37476 6866 37504 8910
rect 37752 8634 37780 9522
rect 37844 8634 37872 14758
rect 39264 14716 39572 14725
rect 39264 14714 39270 14716
rect 39326 14714 39350 14716
rect 39406 14714 39430 14716
rect 39486 14714 39510 14716
rect 39566 14714 39572 14716
rect 39326 14662 39328 14714
rect 39508 14662 39510 14714
rect 39264 14660 39270 14662
rect 39326 14660 39350 14662
rect 39406 14660 39430 14662
rect 39486 14660 39510 14662
rect 39566 14660 39572 14662
rect 39264 14651 39572 14660
rect 42708 14612 42760 14618
rect 42708 14554 42760 14560
rect 40960 14408 41012 14414
rect 40960 14350 41012 14356
rect 40500 14272 40552 14278
rect 40500 14214 40552 14220
rect 38384 13932 38436 13938
rect 38384 13874 38436 13880
rect 38396 13190 38424 13874
rect 38936 13864 38988 13870
rect 38936 13806 38988 13812
rect 38384 13184 38436 13190
rect 38384 13126 38436 13132
rect 38660 13184 38712 13190
rect 38660 13126 38712 13132
rect 38672 12850 38700 13126
rect 37924 12844 37976 12850
rect 37924 12786 37976 12792
rect 38660 12844 38712 12850
rect 38660 12786 38712 12792
rect 37936 12442 37964 12786
rect 38568 12708 38620 12714
rect 38568 12650 38620 12656
rect 37924 12436 37976 12442
rect 37924 12378 37976 12384
rect 38016 12368 38068 12374
rect 38016 12310 38068 12316
rect 37924 12232 37976 12238
rect 38028 12220 38056 12310
rect 38108 12232 38160 12238
rect 38028 12192 38108 12220
rect 37924 12174 37976 12180
rect 38108 12174 38160 12180
rect 37936 11082 37964 12174
rect 38108 12096 38160 12102
rect 38108 12038 38160 12044
rect 38384 12096 38436 12102
rect 38384 12038 38436 12044
rect 38120 11898 38148 12038
rect 38108 11892 38160 11898
rect 38108 11834 38160 11840
rect 38396 11762 38424 12038
rect 38580 11898 38608 12650
rect 38672 12434 38700 12786
rect 38672 12406 38792 12434
rect 38660 12368 38712 12374
rect 38660 12310 38712 12316
rect 38672 12170 38700 12310
rect 38764 12238 38792 12406
rect 38752 12232 38804 12238
rect 38752 12174 38804 12180
rect 38660 12164 38712 12170
rect 38660 12106 38712 12112
rect 38568 11892 38620 11898
rect 38568 11834 38620 11840
rect 38384 11756 38436 11762
rect 38384 11698 38436 11704
rect 38108 11688 38160 11694
rect 38108 11630 38160 11636
rect 38016 11144 38068 11150
rect 38016 11086 38068 11092
rect 37924 11076 37976 11082
rect 37924 11018 37976 11024
rect 38028 10266 38056 11086
rect 38016 10260 38068 10266
rect 38016 10202 38068 10208
rect 37924 8832 37976 8838
rect 37924 8774 37976 8780
rect 37740 8628 37792 8634
rect 37740 8570 37792 8576
rect 37832 8628 37884 8634
rect 37832 8570 37884 8576
rect 37936 8498 37964 8774
rect 37924 8492 37976 8498
rect 37924 8434 37976 8440
rect 37936 7954 37964 8434
rect 37924 7948 37976 7954
rect 37924 7890 37976 7896
rect 37464 6860 37516 6866
rect 37464 6802 37516 6808
rect 36268 6384 36320 6390
rect 36268 6326 36320 6332
rect 34980 6316 35032 6322
rect 34980 6258 35032 6264
rect 35900 6316 35952 6322
rect 35900 6258 35952 6264
rect 36084 6316 36136 6322
rect 36084 6258 36136 6264
rect 35348 6112 35400 6118
rect 35348 6054 35400 6060
rect 35360 5778 35388 6054
rect 35912 5914 35940 6258
rect 35992 6112 36044 6118
rect 35992 6054 36044 6060
rect 35900 5908 35952 5914
rect 35900 5850 35952 5856
rect 35348 5772 35400 5778
rect 35348 5714 35400 5720
rect 34152 5364 34204 5370
rect 34152 5306 34204 5312
rect 34612 5364 34664 5370
rect 34612 5306 34664 5312
rect 35440 5364 35492 5370
rect 35440 5306 35492 5312
rect 33692 4820 33744 4826
rect 33692 4762 33744 4768
rect 33140 4752 33192 4758
rect 33140 4694 33192 4700
rect 33324 4752 33376 4758
rect 33324 4694 33376 4700
rect 35452 4690 35480 5306
rect 35900 5092 35952 5098
rect 35900 5034 35952 5040
rect 35440 4684 35492 4690
rect 35440 4626 35492 4632
rect 32864 4616 32916 4622
rect 33876 4616 33928 4622
rect 32864 4558 32916 4564
rect 33874 4584 33876 4593
rect 33928 4584 33930 4593
rect 32876 4010 32904 4558
rect 33508 4548 33560 4554
rect 33874 4519 33930 4528
rect 35072 4548 35124 4554
rect 33508 4490 33560 4496
rect 35072 4490 35124 4496
rect 33140 4480 33192 4486
rect 33140 4422 33192 4428
rect 33152 4146 33180 4422
rect 33520 4146 33548 4490
rect 33790 4380 34098 4389
rect 33790 4378 33796 4380
rect 33852 4378 33876 4380
rect 33932 4378 33956 4380
rect 34012 4378 34036 4380
rect 34092 4378 34098 4380
rect 33852 4326 33854 4378
rect 34034 4326 34036 4378
rect 33790 4324 33796 4326
rect 33852 4324 33876 4326
rect 33932 4324 33956 4326
rect 34012 4324 34036 4326
rect 34092 4324 34098 4326
rect 33790 4315 34098 4324
rect 33140 4140 33192 4146
rect 33140 4082 33192 4088
rect 33508 4140 33560 4146
rect 33508 4082 33560 4088
rect 35084 4010 35112 4490
rect 35912 4146 35940 5034
rect 36004 5030 36032 6054
rect 36096 5574 36124 6258
rect 37476 5778 37504 6802
rect 37464 5772 37516 5778
rect 37464 5714 37516 5720
rect 37188 5636 37240 5642
rect 37188 5578 37240 5584
rect 36084 5568 36136 5574
rect 36084 5510 36136 5516
rect 36912 5568 36964 5574
rect 36912 5510 36964 5516
rect 36924 5370 36952 5510
rect 36912 5364 36964 5370
rect 36912 5306 36964 5312
rect 36268 5228 36320 5234
rect 36268 5170 36320 5176
rect 35992 5024 36044 5030
rect 35992 4966 36044 4972
rect 35900 4140 35952 4146
rect 35900 4082 35952 4088
rect 36280 4078 36308 5170
rect 37200 4826 37228 5578
rect 37372 5228 37424 5234
rect 37372 5170 37424 5176
rect 37188 4820 37240 4826
rect 37188 4762 37240 4768
rect 37384 4622 37412 5170
rect 37372 4616 37424 4622
rect 37372 4558 37424 4564
rect 37384 4146 37412 4558
rect 37476 4146 37504 5714
rect 38016 5636 38068 5642
rect 38016 5578 38068 5584
rect 38028 4826 38056 5578
rect 38016 4820 38068 4826
rect 38016 4762 38068 4768
rect 36360 4140 36412 4146
rect 36360 4082 36412 4088
rect 37372 4140 37424 4146
rect 37372 4082 37424 4088
rect 37464 4140 37516 4146
rect 37464 4082 37516 4088
rect 36268 4072 36320 4078
rect 36268 4014 36320 4020
rect 32864 4004 32916 4010
rect 32864 3946 32916 3952
rect 35072 4004 35124 4010
rect 35072 3946 35124 3952
rect 32876 3738 32904 3946
rect 36372 3942 36400 4082
rect 36360 3936 36412 3942
rect 36360 3878 36412 3884
rect 32864 3732 32916 3738
rect 32864 3674 32916 3680
rect 33508 3596 33560 3602
rect 33508 3538 33560 3544
rect 32588 2508 32640 2514
rect 32588 2450 32640 2456
rect 32220 2440 32272 2446
rect 32220 2382 32272 2388
rect 31852 2304 31904 2310
rect 31852 2246 31904 2252
rect 30300 870 30420 898
rect 30300 800 30328 870
rect 32232 800 32260 2382
rect 33520 800 33548 3538
rect 36372 3466 36400 3878
rect 37384 3534 37412 4082
rect 37372 3528 37424 3534
rect 37372 3470 37424 3476
rect 36360 3460 36412 3466
rect 36360 3402 36412 3408
rect 33790 3292 34098 3301
rect 33790 3290 33796 3292
rect 33852 3290 33876 3292
rect 33932 3290 33956 3292
rect 34012 3290 34036 3292
rect 34092 3290 34098 3292
rect 33852 3238 33854 3290
rect 34034 3238 34036 3290
rect 33790 3236 33796 3238
rect 33852 3236 33876 3238
rect 33932 3236 33956 3238
rect 34012 3236 34036 3238
rect 34092 3236 34098 3238
rect 33790 3227 34098 3236
rect 35532 2848 35584 2854
rect 35532 2790 35584 2796
rect 35544 2446 35572 2790
rect 38120 2650 38148 11630
rect 38292 11620 38344 11626
rect 38292 11562 38344 11568
rect 38304 11150 38332 11562
rect 38396 11286 38424 11698
rect 38384 11280 38436 11286
rect 38384 11222 38436 11228
rect 38476 11280 38528 11286
rect 38476 11222 38528 11228
rect 38488 11150 38516 11222
rect 38672 11150 38700 12106
rect 38764 11370 38792 12174
rect 38844 12096 38896 12102
rect 38844 12038 38896 12044
rect 38856 11762 38884 12038
rect 38948 11898 38976 13806
rect 39264 13628 39572 13637
rect 39264 13626 39270 13628
rect 39326 13626 39350 13628
rect 39406 13626 39430 13628
rect 39486 13626 39510 13628
rect 39566 13626 39572 13628
rect 39326 13574 39328 13626
rect 39508 13574 39510 13626
rect 39264 13572 39270 13574
rect 39326 13572 39350 13574
rect 39406 13572 39430 13574
rect 39486 13572 39510 13574
rect 39566 13572 39572 13574
rect 39264 13563 39572 13572
rect 40512 13326 40540 14214
rect 40592 13796 40644 13802
rect 40592 13738 40644 13744
rect 40604 13326 40632 13738
rect 40500 13320 40552 13326
rect 39394 13288 39450 13297
rect 40500 13262 40552 13268
rect 40592 13320 40644 13326
rect 40592 13262 40644 13268
rect 39394 13223 39450 13232
rect 40132 13252 40184 13258
rect 39408 12782 39436 13223
rect 40132 13194 40184 13200
rect 40040 12980 40092 12986
rect 40040 12922 40092 12928
rect 39764 12912 39816 12918
rect 39764 12854 39816 12860
rect 39396 12776 39448 12782
rect 39396 12718 39448 12724
rect 39264 12540 39572 12549
rect 39264 12538 39270 12540
rect 39326 12538 39350 12540
rect 39406 12538 39430 12540
rect 39486 12538 39510 12540
rect 39566 12538 39572 12540
rect 39326 12486 39328 12538
rect 39508 12486 39510 12538
rect 39264 12484 39270 12486
rect 39326 12484 39350 12486
rect 39406 12484 39430 12486
rect 39486 12484 39510 12486
rect 39566 12484 39572 12486
rect 39264 12475 39572 12484
rect 39132 12406 39344 12434
rect 39132 12238 39160 12406
rect 39212 12368 39264 12374
rect 39212 12310 39264 12316
rect 39224 12238 39252 12310
rect 39120 12232 39172 12238
rect 39120 12174 39172 12180
rect 39212 12232 39264 12238
rect 39212 12174 39264 12180
rect 39028 12164 39080 12170
rect 39028 12106 39080 12112
rect 38936 11892 38988 11898
rect 38936 11834 38988 11840
rect 38844 11756 38896 11762
rect 38844 11698 38896 11704
rect 38764 11342 38976 11370
rect 38948 11218 38976 11342
rect 38752 11212 38804 11218
rect 38752 11154 38804 11160
rect 38936 11212 38988 11218
rect 38936 11154 38988 11160
rect 38292 11144 38344 11150
rect 38292 11086 38344 11092
rect 38476 11144 38528 11150
rect 38476 11086 38528 11092
rect 38660 11144 38712 11150
rect 38660 11086 38712 11092
rect 38304 10554 38332 11086
rect 38660 10736 38712 10742
rect 38660 10678 38712 10684
rect 38304 10538 38516 10554
rect 38304 10532 38528 10538
rect 38304 10526 38476 10532
rect 38304 10266 38332 10526
rect 38476 10474 38528 10480
rect 38292 10260 38344 10266
rect 38292 10202 38344 10208
rect 38672 10062 38700 10678
rect 38764 10266 38792 11154
rect 38844 11144 38896 11150
rect 38844 11086 38896 11092
rect 38856 10810 38884 11086
rect 39040 10810 39068 12106
rect 39120 12096 39172 12102
rect 39120 12038 39172 12044
rect 39132 11286 39160 12038
rect 39210 11792 39266 11801
rect 39316 11778 39344 12406
rect 39266 11750 39344 11778
rect 39210 11727 39266 11736
rect 39224 11694 39252 11727
rect 39212 11688 39264 11694
rect 39212 11630 39264 11636
rect 39264 11452 39572 11461
rect 39264 11450 39270 11452
rect 39326 11450 39350 11452
rect 39406 11450 39430 11452
rect 39486 11450 39510 11452
rect 39566 11450 39572 11452
rect 39326 11398 39328 11450
rect 39508 11398 39510 11450
rect 39264 11396 39270 11398
rect 39326 11396 39350 11398
rect 39406 11396 39430 11398
rect 39486 11396 39510 11398
rect 39566 11396 39572 11398
rect 39264 11387 39572 11396
rect 39120 11280 39172 11286
rect 39120 11222 39172 11228
rect 39776 11150 39804 12854
rect 40052 12628 40080 12922
rect 40144 12782 40172 13194
rect 40408 13184 40460 13190
rect 40408 13126 40460 13132
rect 40316 12980 40368 12986
rect 40316 12922 40368 12928
rect 40132 12776 40184 12782
rect 40184 12736 40264 12764
rect 40132 12718 40184 12724
rect 40132 12640 40184 12646
rect 40052 12600 40132 12628
rect 40132 12582 40184 12588
rect 40236 12374 40264 12736
rect 40224 12368 40276 12374
rect 40224 12310 40276 12316
rect 40040 12300 40092 12306
rect 40040 12242 40092 12248
rect 40052 11626 40080 12242
rect 40328 12170 40356 12922
rect 40420 12306 40448 13126
rect 40512 12986 40540 13262
rect 40500 12980 40552 12986
rect 40500 12922 40552 12928
rect 40408 12300 40460 12306
rect 40408 12242 40460 12248
rect 40316 12164 40368 12170
rect 40316 12106 40368 12112
rect 40040 11620 40092 11626
rect 40040 11562 40092 11568
rect 40604 11218 40632 13262
rect 40972 12646 41000 14350
rect 41972 14272 42024 14278
rect 41972 14214 42024 14220
rect 41984 14006 42012 14214
rect 41972 14000 42024 14006
rect 41972 13942 42024 13948
rect 42064 13728 42116 13734
rect 42064 13670 42116 13676
rect 41972 13388 42024 13394
rect 41972 13330 42024 13336
rect 41052 13252 41104 13258
rect 41052 13194 41104 13200
rect 41696 13252 41748 13258
rect 41696 13194 41748 13200
rect 41064 12986 41092 13194
rect 41052 12980 41104 12986
rect 41052 12922 41104 12928
rect 41512 12844 41564 12850
rect 41512 12786 41564 12792
rect 40960 12640 41012 12646
rect 40960 12582 41012 12588
rect 41420 12232 41472 12238
rect 41420 12174 41472 12180
rect 40868 12096 40920 12102
rect 40868 12038 40920 12044
rect 40880 11830 40908 12038
rect 41432 11898 41460 12174
rect 41524 12170 41552 12786
rect 41708 12782 41736 13194
rect 41696 12776 41748 12782
rect 41880 12776 41932 12782
rect 41696 12718 41748 12724
rect 41878 12744 41880 12753
rect 41932 12744 41934 12753
rect 41984 12730 42012 13330
rect 42076 13326 42104 13670
rect 42720 13530 42748 14554
rect 42982 14512 43038 14521
rect 42982 14447 43038 14456
rect 42996 14414 43024 14447
rect 42984 14408 43036 14414
rect 42984 14350 43036 14356
rect 44270 14376 44326 14385
rect 44270 14311 44326 14320
rect 44284 14278 44312 14311
rect 44272 14272 44324 14278
rect 44272 14214 44324 14220
rect 44737 14172 45045 14181
rect 44737 14170 44743 14172
rect 44799 14170 44823 14172
rect 44879 14170 44903 14172
rect 44959 14170 44983 14172
rect 45039 14170 45045 14172
rect 44799 14118 44801 14170
rect 44981 14118 44983 14170
rect 44737 14116 44743 14118
rect 44799 14116 44823 14118
rect 44879 14116 44903 14118
rect 44959 14116 44983 14118
rect 45039 14116 45045 14118
rect 44737 14107 45045 14116
rect 42708 13524 42760 13530
rect 42708 13466 42760 13472
rect 42064 13320 42116 13326
rect 42064 13262 42116 13268
rect 42076 12986 42104 13262
rect 42340 13184 42392 13190
rect 42340 13126 42392 13132
rect 42064 12980 42116 12986
rect 42064 12922 42116 12928
rect 42352 12850 42380 13126
rect 44737 13084 45045 13093
rect 44737 13082 44743 13084
rect 44799 13082 44823 13084
rect 44879 13082 44903 13084
rect 44959 13082 44983 13084
rect 45039 13082 45045 13084
rect 44799 13030 44801 13082
rect 44981 13030 44983 13082
rect 44737 13028 44743 13030
rect 44799 13028 44823 13030
rect 44879 13028 44903 13030
rect 44959 13028 44983 13030
rect 45039 13028 45045 13030
rect 44737 13019 45045 13028
rect 42340 12844 42392 12850
rect 42340 12786 42392 12792
rect 41604 12640 41656 12646
rect 41604 12582 41656 12588
rect 41512 12164 41564 12170
rect 41512 12106 41564 12112
rect 41420 11892 41472 11898
rect 41420 11834 41472 11840
rect 40868 11824 40920 11830
rect 40868 11766 40920 11772
rect 41524 11762 41552 12106
rect 41616 11762 41644 12582
rect 41708 12434 41736 12718
rect 41934 12702 42012 12730
rect 41878 12679 41934 12688
rect 41708 12406 41828 12434
rect 41708 12306 41736 12406
rect 41696 12300 41748 12306
rect 41696 12242 41748 12248
rect 41696 12096 41748 12102
rect 41696 12038 41748 12044
rect 41512 11756 41564 11762
rect 41512 11698 41564 11704
rect 41604 11756 41656 11762
rect 41604 11698 41656 11704
rect 40592 11212 40644 11218
rect 40592 11154 40644 11160
rect 41708 11150 41736 12038
rect 41800 11830 41828 12406
rect 41984 12238 42012 12702
rect 45008 12640 45060 12646
rect 45008 12582 45060 12588
rect 45020 12345 45048 12582
rect 45006 12336 45062 12345
rect 45006 12271 45062 12280
rect 41972 12232 42024 12238
rect 41972 12174 42024 12180
rect 42248 12232 42300 12238
rect 42248 12174 42300 12180
rect 41788 11824 41840 11830
rect 41788 11766 41840 11772
rect 41984 11762 42012 12174
rect 42260 11830 42288 12174
rect 44737 11996 45045 12005
rect 44737 11994 44743 11996
rect 44799 11994 44823 11996
rect 44879 11994 44903 11996
rect 44959 11994 44983 11996
rect 45039 11994 45045 11996
rect 44799 11942 44801 11994
rect 44981 11942 44983 11994
rect 44737 11940 44743 11942
rect 44799 11940 44823 11942
rect 44879 11940 44903 11942
rect 44959 11940 44983 11942
rect 45039 11940 45045 11942
rect 44737 11931 45045 11940
rect 42248 11824 42300 11830
rect 42248 11766 42300 11772
rect 42800 11824 42852 11830
rect 42800 11766 42852 11772
rect 41972 11756 42024 11762
rect 41972 11698 42024 11704
rect 39764 11144 39816 11150
rect 39764 11086 39816 11092
rect 41696 11144 41748 11150
rect 41696 11086 41748 11092
rect 42812 11014 42840 11766
rect 43168 11688 43220 11694
rect 43168 11630 43220 11636
rect 42892 11076 42944 11082
rect 42892 11018 42944 11024
rect 42800 11008 42852 11014
rect 42800 10950 42852 10956
rect 38844 10804 38896 10810
rect 38844 10746 38896 10752
rect 39028 10804 39080 10810
rect 39028 10746 39080 10752
rect 42812 10674 42840 10950
rect 42800 10668 42852 10674
rect 42800 10610 42852 10616
rect 39264 10364 39572 10373
rect 39264 10362 39270 10364
rect 39326 10362 39350 10364
rect 39406 10362 39430 10364
rect 39486 10362 39510 10364
rect 39566 10362 39572 10364
rect 39326 10310 39328 10362
rect 39508 10310 39510 10362
rect 39264 10308 39270 10310
rect 39326 10308 39350 10310
rect 39406 10308 39430 10310
rect 39486 10308 39510 10310
rect 39566 10308 39572 10310
rect 39264 10299 39572 10308
rect 42904 10266 42932 11018
rect 43180 10810 43208 11630
rect 45008 11144 45060 11150
rect 45006 11112 45008 11121
rect 45060 11112 45062 11121
rect 45006 11047 45062 11056
rect 44737 10908 45045 10917
rect 44737 10906 44743 10908
rect 44799 10906 44823 10908
rect 44879 10906 44903 10908
rect 44959 10906 44983 10908
rect 45039 10906 45045 10908
rect 44799 10854 44801 10906
rect 44981 10854 44983 10906
rect 44737 10852 44743 10854
rect 44799 10852 44823 10854
rect 44879 10852 44903 10854
rect 44959 10852 44983 10854
rect 45039 10852 45045 10854
rect 44737 10843 45045 10852
rect 43168 10804 43220 10810
rect 43168 10746 43220 10752
rect 44456 10736 44508 10742
rect 44456 10678 44508 10684
rect 44272 10600 44324 10606
rect 44272 10542 44324 10548
rect 38752 10260 38804 10266
rect 38752 10202 38804 10208
rect 42892 10260 42944 10266
rect 42892 10202 42944 10208
rect 38660 10056 38712 10062
rect 38660 9998 38712 10004
rect 43444 10056 43496 10062
rect 43444 9998 43496 10004
rect 39264 9276 39572 9285
rect 39264 9274 39270 9276
rect 39326 9274 39350 9276
rect 39406 9274 39430 9276
rect 39486 9274 39510 9276
rect 39566 9274 39572 9276
rect 39326 9222 39328 9274
rect 39508 9222 39510 9274
rect 39264 9220 39270 9222
rect 39326 9220 39350 9222
rect 39406 9220 39430 9222
rect 39486 9220 39510 9222
rect 39566 9220 39572 9222
rect 39264 9211 39572 9220
rect 38936 8900 38988 8906
rect 38936 8842 38988 8848
rect 38948 7818 38976 8842
rect 42616 8492 42668 8498
rect 42616 8434 42668 8440
rect 41420 8356 41472 8362
rect 41420 8298 41472 8304
rect 39264 8188 39572 8197
rect 39264 8186 39270 8188
rect 39326 8186 39350 8188
rect 39406 8186 39430 8188
rect 39486 8186 39510 8188
rect 39566 8186 39572 8188
rect 39326 8134 39328 8186
rect 39508 8134 39510 8186
rect 39264 8132 39270 8134
rect 39326 8132 39350 8134
rect 39406 8132 39430 8134
rect 39486 8132 39510 8134
rect 39566 8132 39572 8134
rect 39264 8123 39572 8132
rect 40500 8084 40552 8090
rect 40500 8026 40552 8032
rect 39120 7880 39172 7886
rect 39120 7822 39172 7828
rect 39304 7880 39356 7886
rect 39304 7822 39356 7828
rect 40040 7880 40092 7886
rect 40040 7822 40092 7828
rect 38936 7812 38988 7818
rect 38936 7754 38988 7760
rect 38752 7744 38804 7750
rect 38752 7686 38804 7692
rect 38764 7478 38792 7686
rect 38948 7478 38976 7754
rect 38752 7472 38804 7478
rect 38752 7414 38804 7420
rect 38936 7472 38988 7478
rect 38936 7414 38988 7420
rect 39132 7002 39160 7822
rect 39316 7546 39344 7822
rect 39856 7812 39908 7818
rect 39856 7754 39908 7760
rect 39304 7540 39356 7546
rect 39304 7482 39356 7488
rect 39868 7410 39896 7754
rect 39856 7404 39908 7410
rect 39856 7346 39908 7352
rect 39264 7100 39572 7109
rect 39264 7098 39270 7100
rect 39326 7098 39350 7100
rect 39406 7098 39430 7100
rect 39486 7098 39510 7100
rect 39566 7098 39572 7100
rect 39326 7046 39328 7098
rect 39508 7046 39510 7098
rect 39264 7044 39270 7046
rect 39326 7044 39350 7046
rect 39406 7044 39430 7046
rect 39486 7044 39510 7046
rect 39566 7044 39572 7046
rect 39264 7035 39572 7044
rect 39120 6996 39172 7002
rect 39120 6938 39172 6944
rect 39488 6996 39540 7002
rect 39488 6938 39540 6944
rect 38476 6792 38528 6798
rect 38476 6734 38528 6740
rect 38488 6458 38516 6734
rect 38936 6724 38988 6730
rect 38936 6666 38988 6672
rect 38476 6452 38528 6458
rect 38476 6394 38528 6400
rect 38948 6390 38976 6666
rect 39500 6458 39528 6938
rect 39868 6934 39896 7346
rect 39948 7200 40000 7206
rect 39948 7142 40000 7148
rect 39856 6928 39908 6934
rect 39856 6870 39908 6876
rect 39960 6798 39988 7142
rect 40052 7002 40080 7822
rect 40316 7812 40368 7818
rect 40316 7754 40368 7760
rect 40224 7744 40276 7750
rect 40224 7686 40276 7692
rect 40236 7478 40264 7686
rect 40224 7472 40276 7478
rect 40224 7414 40276 7420
rect 40224 7336 40276 7342
rect 40224 7278 40276 7284
rect 40236 7002 40264 7278
rect 40328 7274 40356 7754
rect 40408 7744 40460 7750
rect 40408 7686 40460 7692
rect 40316 7268 40368 7274
rect 40316 7210 40368 7216
rect 40040 6996 40092 7002
rect 40040 6938 40092 6944
rect 40224 6996 40276 7002
rect 40224 6938 40276 6944
rect 39948 6792 40000 6798
rect 39948 6734 40000 6740
rect 39672 6656 39724 6662
rect 39672 6598 39724 6604
rect 39488 6452 39540 6458
rect 39488 6394 39540 6400
rect 38936 6384 38988 6390
rect 38936 6326 38988 6332
rect 38948 6254 38976 6326
rect 39500 6322 39528 6394
rect 39488 6316 39540 6322
rect 39488 6258 39540 6264
rect 38936 6248 38988 6254
rect 38936 6190 38988 6196
rect 38948 5930 38976 6190
rect 39120 6112 39172 6118
rect 39120 6054 39172 6060
rect 38948 5902 39068 5930
rect 39040 5846 39068 5902
rect 39028 5840 39080 5846
rect 39028 5782 39080 5788
rect 38660 5636 38712 5642
rect 38660 5578 38712 5584
rect 38672 5234 38700 5578
rect 39132 5370 39160 6054
rect 39264 6012 39572 6021
rect 39264 6010 39270 6012
rect 39326 6010 39350 6012
rect 39406 6010 39430 6012
rect 39486 6010 39510 6012
rect 39566 6010 39572 6012
rect 39326 5958 39328 6010
rect 39508 5958 39510 6010
rect 39264 5956 39270 5958
rect 39326 5956 39350 5958
rect 39406 5956 39430 5958
rect 39486 5956 39510 5958
rect 39566 5956 39572 5958
rect 39264 5947 39572 5956
rect 39684 5914 39712 6598
rect 40052 6322 40080 6938
rect 40132 6860 40184 6866
rect 40132 6802 40184 6808
rect 40144 6662 40172 6802
rect 40420 6746 40448 7686
rect 40512 7478 40540 8026
rect 41432 7886 41460 8298
rect 41420 7880 41472 7886
rect 41420 7822 41472 7828
rect 42524 7812 42576 7818
rect 42524 7754 42576 7760
rect 42536 7546 42564 7754
rect 42524 7540 42576 7546
rect 42524 7482 42576 7488
rect 40500 7472 40552 7478
rect 40500 7414 40552 7420
rect 40512 6934 40540 7414
rect 42628 7410 42656 8434
rect 42984 7812 43036 7818
rect 42984 7754 43036 7760
rect 42996 7546 43024 7754
rect 42984 7540 43036 7546
rect 42984 7482 43036 7488
rect 42616 7404 42668 7410
rect 42616 7346 42668 7352
rect 41236 7200 41288 7206
rect 41236 7142 41288 7148
rect 40500 6928 40552 6934
rect 40500 6870 40552 6876
rect 40328 6730 40448 6746
rect 40316 6724 40448 6730
rect 40368 6718 40448 6724
rect 40316 6666 40368 6672
rect 40132 6656 40184 6662
rect 40132 6598 40184 6604
rect 40408 6656 40460 6662
rect 40408 6598 40460 6604
rect 40224 6384 40276 6390
rect 40276 6332 40356 6338
rect 40224 6326 40356 6332
rect 40040 6316 40092 6322
rect 40236 6310 40356 6326
rect 40040 6258 40092 6264
rect 39672 5908 39724 5914
rect 39672 5850 39724 5856
rect 39120 5364 39172 5370
rect 39120 5306 39172 5312
rect 39684 5234 39712 5850
rect 40052 5846 40080 6258
rect 40132 6112 40184 6118
rect 40132 6054 40184 6060
rect 40224 6112 40276 6118
rect 40224 6054 40276 6060
rect 40144 5914 40172 6054
rect 40132 5908 40184 5914
rect 40132 5850 40184 5856
rect 40040 5840 40092 5846
rect 40040 5782 40092 5788
rect 40236 5778 40264 6054
rect 40328 5778 40356 6310
rect 40420 5914 40448 6598
rect 40512 6390 40540 6870
rect 41248 6866 41276 7142
rect 40776 6860 40828 6866
rect 40776 6802 40828 6808
rect 41236 6860 41288 6866
rect 41236 6802 41288 6808
rect 40684 6656 40736 6662
rect 40684 6598 40736 6604
rect 40500 6384 40552 6390
rect 40500 6326 40552 6332
rect 40592 6248 40644 6254
rect 40592 6190 40644 6196
rect 40408 5908 40460 5914
rect 40408 5850 40460 5856
rect 40500 5908 40552 5914
rect 40500 5850 40552 5856
rect 40224 5772 40276 5778
rect 40224 5714 40276 5720
rect 40316 5772 40368 5778
rect 40316 5714 40368 5720
rect 40132 5704 40184 5710
rect 40132 5646 40184 5652
rect 40144 5302 40172 5646
rect 40512 5370 40540 5850
rect 40604 5370 40632 6190
rect 40500 5364 40552 5370
rect 40500 5306 40552 5312
rect 40592 5364 40644 5370
rect 40592 5306 40644 5312
rect 40696 5302 40724 6598
rect 40132 5296 40184 5302
rect 40132 5238 40184 5244
rect 40684 5296 40736 5302
rect 40684 5238 40736 5244
rect 40788 5234 40816 6802
rect 42628 6798 42656 7346
rect 40868 6792 40920 6798
rect 40868 6734 40920 6740
rect 42616 6792 42668 6798
rect 42616 6734 42668 6740
rect 40880 6458 40908 6734
rect 42248 6656 42300 6662
rect 42248 6598 42300 6604
rect 40868 6452 40920 6458
rect 40868 6394 40920 6400
rect 40880 5914 40908 6394
rect 40868 5908 40920 5914
rect 40868 5850 40920 5856
rect 42260 5710 42288 6598
rect 42628 6322 42656 6734
rect 42616 6316 42668 6322
rect 42616 6258 42668 6264
rect 42248 5704 42300 5710
rect 42248 5646 42300 5652
rect 41144 5636 41196 5642
rect 41144 5578 41196 5584
rect 41052 5568 41104 5574
rect 41052 5510 41104 5516
rect 41064 5234 41092 5510
rect 38660 5228 38712 5234
rect 38660 5170 38712 5176
rect 39672 5228 39724 5234
rect 39672 5170 39724 5176
rect 40776 5228 40828 5234
rect 40776 5170 40828 5176
rect 41052 5228 41104 5234
rect 41052 5170 41104 5176
rect 41156 5098 41184 5578
rect 42984 5228 43036 5234
rect 42984 5170 43036 5176
rect 41144 5092 41196 5098
rect 41144 5034 41196 5040
rect 38844 5024 38896 5030
rect 38844 4966 38896 4972
rect 38856 4622 38884 4966
rect 39264 4924 39572 4933
rect 39264 4922 39270 4924
rect 39326 4922 39350 4924
rect 39406 4922 39430 4924
rect 39486 4922 39510 4924
rect 39566 4922 39572 4924
rect 39326 4870 39328 4922
rect 39508 4870 39510 4922
rect 39264 4868 39270 4870
rect 39326 4868 39350 4870
rect 39406 4868 39430 4870
rect 39486 4868 39510 4870
rect 39566 4868 39572 4870
rect 39264 4859 39572 4868
rect 38844 4616 38896 4622
rect 38844 4558 38896 4564
rect 42996 4282 43024 5170
rect 42984 4276 43036 4282
rect 42984 4218 43036 4224
rect 38200 4208 38252 4214
rect 38200 4150 38252 4156
rect 38212 3738 38240 4150
rect 39264 3836 39572 3845
rect 39264 3834 39270 3836
rect 39326 3834 39350 3836
rect 39406 3834 39430 3836
rect 39486 3834 39510 3836
rect 39566 3834 39572 3836
rect 39326 3782 39328 3834
rect 39508 3782 39510 3834
rect 39264 3780 39270 3782
rect 39326 3780 39350 3782
rect 39406 3780 39430 3782
rect 39486 3780 39510 3782
rect 39566 3780 39572 3782
rect 39264 3771 39572 3780
rect 38200 3732 38252 3738
rect 38200 3674 38252 3680
rect 39264 2748 39572 2757
rect 39264 2746 39270 2748
rect 39326 2746 39350 2748
rect 39406 2746 39430 2748
rect 39486 2746 39510 2748
rect 39566 2746 39572 2748
rect 39326 2694 39328 2746
rect 39508 2694 39510 2746
rect 39264 2692 39270 2694
rect 39326 2692 39350 2694
rect 39406 2692 39430 2694
rect 39486 2692 39510 2694
rect 39566 2692 39572 2694
rect 39264 2683 39572 2692
rect 43456 2650 43484 9998
rect 44088 9648 44140 9654
rect 44088 9590 44140 9596
rect 43996 7744 44048 7750
rect 43996 7686 44048 7692
rect 44008 7002 44036 7686
rect 43996 6996 44048 7002
rect 43996 6938 44048 6944
rect 44100 5710 44128 9590
rect 44178 8936 44234 8945
rect 44178 8871 44234 8880
rect 44192 8838 44220 8871
rect 44180 8832 44232 8838
rect 44180 8774 44232 8780
rect 44284 7546 44312 10542
rect 44364 8968 44416 8974
rect 44362 8936 44364 8945
rect 44416 8936 44418 8945
rect 44362 8871 44418 8880
rect 44272 7540 44324 7546
rect 44272 7482 44324 7488
rect 44362 7440 44418 7449
rect 44362 7375 44364 7384
rect 44416 7375 44418 7384
rect 44364 7346 44416 7352
rect 44088 5704 44140 5710
rect 44088 5646 44140 5652
rect 44088 5024 44140 5030
rect 44088 4966 44140 4972
rect 44100 4622 44128 4966
rect 44088 4616 44140 4622
rect 44088 4558 44140 4564
rect 44272 4480 44324 4486
rect 44272 4422 44324 4428
rect 44284 4185 44312 4422
rect 44270 4176 44326 4185
rect 44270 4111 44326 4120
rect 44088 3936 44140 3942
rect 44088 3878 44140 3884
rect 38108 2644 38160 2650
rect 38108 2586 38160 2592
rect 43444 2644 43496 2650
rect 43444 2586 43496 2592
rect 44100 2446 44128 3878
rect 44468 3194 44496 10678
rect 44737 9820 45045 9829
rect 44737 9818 44743 9820
rect 44799 9818 44823 9820
rect 44879 9818 44903 9820
rect 44959 9818 44983 9820
rect 45039 9818 45045 9820
rect 44799 9766 44801 9818
rect 44981 9766 44983 9818
rect 44737 9764 44743 9766
rect 44799 9764 44823 9766
rect 44879 9764 44903 9766
rect 44959 9764 44983 9766
rect 45039 9764 45045 9766
rect 44737 9755 45045 9764
rect 44737 8732 45045 8741
rect 44737 8730 44743 8732
rect 44799 8730 44823 8732
rect 44879 8730 44903 8732
rect 44959 8730 44983 8732
rect 45039 8730 45045 8732
rect 44799 8678 44801 8730
rect 44981 8678 44983 8730
rect 44737 8676 44743 8678
rect 44799 8676 44823 8678
rect 44879 8676 44903 8678
rect 44959 8676 44983 8678
rect 45039 8676 45045 8678
rect 44737 8667 45045 8676
rect 44737 7644 45045 7653
rect 44737 7642 44743 7644
rect 44799 7642 44823 7644
rect 44879 7642 44903 7644
rect 44959 7642 44983 7644
rect 45039 7642 45045 7644
rect 44799 7590 44801 7642
rect 44981 7590 44983 7642
rect 44737 7588 44743 7590
rect 44799 7588 44823 7590
rect 44879 7588 44903 7590
rect 44959 7588 44983 7590
rect 45039 7588 45045 7590
rect 44737 7579 45045 7588
rect 44737 6556 45045 6565
rect 44737 6554 44743 6556
rect 44799 6554 44823 6556
rect 44879 6554 44903 6556
rect 44959 6554 44983 6556
rect 45039 6554 45045 6556
rect 44799 6502 44801 6554
rect 44981 6502 44983 6554
rect 44737 6500 44743 6502
rect 44799 6500 44823 6502
rect 44879 6500 44903 6502
rect 44959 6500 44983 6502
rect 45039 6500 45045 6502
rect 44737 6491 45045 6500
rect 45006 5672 45062 5681
rect 45006 5607 45062 5616
rect 45020 5574 45048 5607
rect 45008 5568 45060 5574
rect 45008 5510 45060 5516
rect 44737 5468 45045 5477
rect 44737 5466 44743 5468
rect 44799 5466 44823 5468
rect 44879 5466 44903 5468
rect 44959 5466 44983 5468
rect 45039 5466 45045 5468
rect 44799 5414 44801 5466
rect 44981 5414 44983 5466
rect 44737 5412 44743 5414
rect 44799 5412 44823 5414
rect 44879 5412 44903 5414
rect 44959 5412 44983 5414
rect 45039 5412 45045 5414
rect 44737 5403 45045 5412
rect 44737 4380 45045 4389
rect 44737 4378 44743 4380
rect 44799 4378 44823 4380
rect 44879 4378 44903 4380
rect 44959 4378 44983 4380
rect 45039 4378 45045 4380
rect 44799 4326 44801 4378
rect 44981 4326 44983 4378
rect 44737 4324 44743 4326
rect 44799 4324 44823 4326
rect 44879 4324 44903 4326
rect 44959 4324 44983 4326
rect 45039 4324 45045 4326
rect 44737 4315 45045 4324
rect 44640 3528 44692 3534
rect 44640 3470 44692 3476
rect 44456 3188 44508 3194
rect 44456 3130 44508 3136
rect 35532 2440 35584 2446
rect 35532 2382 35584 2388
rect 37648 2440 37700 2446
rect 37648 2382 37700 2388
rect 38660 2440 38712 2446
rect 38660 2382 38712 2388
rect 40040 2440 40092 2446
rect 40040 2382 40092 2388
rect 43812 2440 43864 2446
rect 43812 2382 43864 2388
rect 44088 2440 44140 2446
rect 44088 2382 44140 2388
rect 35440 2304 35492 2310
rect 35440 2246 35492 2252
rect 33790 2204 34098 2213
rect 33790 2202 33796 2204
rect 33852 2202 33876 2204
rect 33932 2202 33956 2204
rect 34012 2202 34036 2204
rect 34092 2202 34098 2204
rect 33852 2150 33854 2202
rect 34034 2150 34036 2202
rect 33790 2148 33796 2150
rect 33852 2148 33876 2150
rect 33932 2148 33956 2150
rect 34012 2148 34036 2150
rect 34092 2148 34098 2150
rect 33790 2139 34098 2148
rect 35452 800 35480 2246
rect 37660 950 37688 2382
rect 36728 944 36780 950
rect 36728 886 36780 892
rect 37648 944 37700 950
rect 37648 886 37700 892
rect 36740 800 36768 886
rect 38672 800 38700 2382
rect 40052 898 40080 2382
rect 41880 2372 41932 2378
rect 41880 2314 41932 2320
rect 39960 870 40080 898
rect 39960 800 39988 870
rect 41892 800 41920 2314
rect 43824 800 43852 2382
rect 44272 2304 44324 2310
rect 44272 2246 44324 2252
rect 44284 2009 44312 2246
rect 44270 2000 44326 2009
rect 44270 1935 44326 1944
rect -10 0 102 800
rect 1278 0 1390 800
rect 3210 0 3322 800
rect 4498 0 4610 800
rect 6430 0 6542 800
rect 7718 0 7830 800
rect 9650 0 9762 800
rect 10938 0 11050 800
rect 12870 0 12982 800
rect 14158 0 14270 800
rect 16090 0 16202 800
rect 17378 0 17490 800
rect 19310 0 19422 800
rect 20598 0 20710 800
rect 22530 0 22642 800
rect 23818 0 23930 800
rect 25750 0 25862 800
rect 27038 0 27150 800
rect 28970 0 29082 800
rect 30258 0 30370 800
rect 32190 0 32302 800
rect 33478 0 33590 800
rect 35410 0 35522 800
rect 36698 0 36810 800
rect 38630 0 38742 800
rect 39918 0 40030 800
rect 41850 0 41962 800
rect 43782 0 43894 800
rect 44652 785 44680 3470
rect 44737 3292 45045 3301
rect 44737 3290 44743 3292
rect 44799 3290 44823 3292
rect 44879 3290 44903 3292
rect 44959 3290 44983 3292
rect 45039 3290 45045 3292
rect 44799 3238 44801 3290
rect 44981 3238 44983 3290
rect 44737 3236 44743 3238
rect 44799 3236 44823 3238
rect 44879 3236 44903 3238
rect 44959 3236 44983 3238
rect 45039 3236 45045 3238
rect 44737 3227 45045 3236
rect 45100 3052 45152 3058
rect 45100 2994 45152 3000
rect 44737 2204 45045 2213
rect 44737 2202 44743 2204
rect 44799 2202 44823 2204
rect 44879 2202 44903 2204
rect 44959 2202 44983 2204
rect 45039 2202 45045 2204
rect 44799 2150 44801 2202
rect 44981 2150 44983 2202
rect 44737 2148 44743 2150
rect 44799 2148 44823 2150
rect 44879 2148 44903 2150
rect 44959 2148 44983 2150
rect 45039 2148 45045 2150
rect 44737 2139 45045 2148
rect 45112 800 45140 2994
rect 44638 776 44694 785
rect 44638 711 44694 720
rect 45070 0 45182 800
<< via2 >>
rect 1030 18400 1086 18456
rect 938 17040 994 17096
rect 11902 17434 11958 17436
rect 11982 17434 12038 17436
rect 12062 17434 12118 17436
rect 12142 17434 12198 17436
rect 11902 17382 11948 17434
rect 11948 17382 11958 17434
rect 11982 17382 12012 17434
rect 12012 17382 12024 17434
rect 12024 17382 12038 17434
rect 12062 17382 12076 17434
rect 12076 17382 12088 17434
rect 12088 17382 12118 17434
rect 12142 17382 12152 17434
rect 12152 17382 12198 17434
rect 11902 17380 11958 17382
rect 11982 17380 12038 17382
rect 12062 17380 12118 17382
rect 12142 17380 12198 17382
rect 22849 17434 22905 17436
rect 22929 17434 22985 17436
rect 23009 17434 23065 17436
rect 23089 17434 23145 17436
rect 22849 17382 22895 17434
rect 22895 17382 22905 17434
rect 22929 17382 22959 17434
rect 22959 17382 22971 17434
rect 22971 17382 22985 17434
rect 23009 17382 23023 17434
rect 23023 17382 23035 17434
rect 23035 17382 23065 17434
rect 23089 17382 23099 17434
rect 23099 17382 23145 17434
rect 22849 17380 22905 17382
rect 22929 17380 22985 17382
rect 23009 17380 23065 17382
rect 23089 17380 23145 17382
rect 33796 17434 33852 17436
rect 33876 17434 33932 17436
rect 33956 17434 34012 17436
rect 34036 17434 34092 17436
rect 33796 17382 33842 17434
rect 33842 17382 33852 17434
rect 33876 17382 33906 17434
rect 33906 17382 33918 17434
rect 33918 17382 33932 17434
rect 33956 17382 33970 17434
rect 33970 17382 33982 17434
rect 33982 17382 34012 17434
rect 34036 17382 34046 17434
rect 34046 17382 34092 17434
rect 33796 17380 33852 17382
rect 33876 17380 33932 17382
rect 33956 17380 34012 17382
rect 34036 17380 34092 17382
rect 938 15000 994 15056
rect 938 13640 994 13696
rect 938 10260 994 10296
rect 938 10240 940 10260
rect 940 10240 992 10260
rect 992 10240 994 10260
rect 3146 12844 3202 12880
rect 3146 12824 3148 12844
rect 3148 12824 3200 12844
rect 3200 12824 3202 12844
rect 6429 16890 6485 16892
rect 6509 16890 6565 16892
rect 6589 16890 6645 16892
rect 6669 16890 6725 16892
rect 6429 16838 6475 16890
rect 6475 16838 6485 16890
rect 6509 16838 6539 16890
rect 6539 16838 6551 16890
rect 6551 16838 6565 16890
rect 6589 16838 6603 16890
rect 6603 16838 6615 16890
rect 6615 16838 6645 16890
rect 6669 16838 6679 16890
rect 6679 16838 6725 16890
rect 6429 16836 6485 16838
rect 6509 16836 6565 16838
rect 6589 16836 6645 16838
rect 6669 16836 6725 16838
rect 6429 15802 6485 15804
rect 6509 15802 6565 15804
rect 6589 15802 6645 15804
rect 6669 15802 6725 15804
rect 6429 15750 6475 15802
rect 6475 15750 6485 15802
rect 6509 15750 6539 15802
rect 6539 15750 6551 15802
rect 6551 15750 6565 15802
rect 6589 15750 6603 15802
rect 6603 15750 6615 15802
rect 6615 15750 6645 15802
rect 6669 15750 6679 15802
rect 6679 15750 6725 15802
rect 6429 15748 6485 15750
rect 6509 15748 6565 15750
rect 6589 15748 6645 15750
rect 6669 15748 6725 15750
rect 6429 14714 6485 14716
rect 6509 14714 6565 14716
rect 6589 14714 6645 14716
rect 6669 14714 6725 14716
rect 6429 14662 6475 14714
rect 6475 14662 6485 14714
rect 6509 14662 6539 14714
rect 6539 14662 6551 14714
rect 6551 14662 6565 14714
rect 6589 14662 6603 14714
rect 6603 14662 6615 14714
rect 6615 14662 6645 14714
rect 6669 14662 6679 14714
rect 6679 14662 6725 14714
rect 6429 14660 6485 14662
rect 6509 14660 6565 14662
rect 6589 14660 6645 14662
rect 6669 14660 6725 14662
rect 11902 16346 11958 16348
rect 11982 16346 12038 16348
rect 12062 16346 12118 16348
rect 12142 16346 12198 16348
rect 11902 16294 11948 16346
rect 11948 16294 11958 16346
rect 11982 16294 12012 16346
rect 12012 16294 12024 16346
rect 12024 16294 12038 16346
rect 12062 16294 12076 16346
rect 12076 16294 12088 16346
rect 12088 16294 12118 16346
rect 12142 16294 12152 16346
rect 12152 16294 12198 16346
rect 11902 16292 11958 16294
rect 11982 16292 12038 16294
rect 12062 16292 12118 16294
rect 12142 16292 12198 16294
rect 11902 15258 11958 15260
rect 11982 15258 12038 15260
rect 12062 15258 12118 15260
rect 12142 15258 12198 15260
rect 11902 15206 11948 15258
rect 11948 15206 11958 15258
rect 11982 15206 12012 15258
rect 12012 15206 12024 15258
rect 12024 15206 12038 15258
rect 12062 15206 12076 15258
rect 12076 15206 12088 15258
rect 12088 15206 12118 15258
rect 12142 15206 12152 15258
rect 12152 15206 12198 15258
rect 11902 15204 11958 15206
rect 11982 15204 12038 15206
rect 12062 15204 12118 15206
rect 12142 15204 12198 15206
rect 4066 11872 4122 11928
rect 4066 11600 4122 11656
rect 938 8200 994 8256
rect 938 6840 994 6896
rect 6429 13626 6485 13628
rect 6509 13626 6565 13628
rect 6589 13626 6645 13628
rect 6669 13626 6725 13628
rect 6429 13574 6475 13626
rect 6475 13574 6485 13626
rect 6509 13574 6539 13626
rect 6539 13574 6551 13626
rect 6551 13574 6565 13626
rect 6589 13574 6603 13626
rect 6603 13574 6615 13626
rect 6615 13574 6645 13626
rect 6669 13574 6679 13626
rect 6679 13574 6725 13626
rect 6429 13572 6485 13574
rect 6509 13572 6565 13574
rect 6589 13572 6645 13574
rect 6669 13572 6725 13574
rect 6429 12538 6485 12540
rect 6509 12538 6565 12540
rect 6589 12538 6645 12540
rect 6669 12538 6725 12540
rect 6429 12486 6475 12538
rect 6475 12486 6485 12538
rect 6509 12486 6539 12538
rect 6539 12486 6551 12538
rect 6551 12486 6565 12538
rect 6589 12486 6603 12538
rect 6603 12486 6615 12538
rect 6615 12486 6645 12538
rect 6669 12486 6679 12538
rect 6679 12486 6725 12538
rect 6429 12484 6485 12486
rect 6509 12484 6565 12486
rect 6589 12484 6645 12486
rect 6669 12484 6725 12486
rect 6429 11450 6485 11452
rect 6509 11450 6565 11452
rect 6589 11450 6645 11452
rect 6669 11450 6725 11452
rect 6429 11398 6475 11450
rect 6475 11398 6485 11450
rect 6509 11398 6539 11450
rect 6539 11398 6551 11450
rect 6551 11398 6565 11450
rect 6589 11398 6603 11450
rect 6603 11398 6615 11450
rect 6615 11398 6645 11450
rect 6669 11398 6679 11450
rect 6679 11398 6725 11450
rect 6429 11396 6485 11398
rect 6509 11396 6565 11398
rect 6589 11396 6645 11398
rect 6669 11396 6725 11398
rect 938 4800 994 4856
rect 6429 10362 6485 10364
rect 6509 10362 6565 10364
rect 6589 10362 6645 10364
rect 6669 10362 6725 10364
rect 6429 10310 6475 10362
rect 6475 10310 6485 10362
rect 6509 10310 6539 10362
rect 6539 10310 6551 10362
rect 6551 10310 6565 10362
rect 6589 10310 6603 10362
rect 6603 10310 6615 10362
rect 6615 10310 6645 10362
rect 6669 10310 6679 10362
rect 6679 10310 6725 10362
rect 6429 10308 6485 10310
rect 6509 10308 6565 10310
rect 6589 10308 6645 10310
rect 6669 10308 6725 10310
rect 11902 14170 11958 14172
rect 11982 14170 12038 14172
rect 12062 14170 12118 14172
rect 12142 14170 12198 14172
rect 11902 14118 11948 14170
rect 11948 14118 11958 14170
rect 11982 14118 12012 14170
rect 12012 14118 12024 14170
rect 12024 14118 12038 14170
rect 12062 14118 12076 14170
rect 12076 14118 12088 14170
rect 12088 14118 12118 14170
rect 12142 14118 12152 14170
rect 12152 14118 12198 14170
rect 11902 14116 11958 14118
rect 11982 14116 12038 14118
rect 12062 14116 12118 14118
rect 12142 14116 12198 14118
rect 6429 9274 6485 9276
rect 6509 9274 6565 9276
rect 6589 9274 6645 9276
rect 6669 9274 6725 9276
rect 6429 9222 6475 9274
rect 6475 9222 6485 9274
rect 6509 9222 6539 9274
rect 6539 9222 6551 9274
rect 6551 9222 6565 9274
rect 6589 9222 6603 9274
rect 6603 9222 6615 9274
rect 6615 9222 6645 9274
rect 6669 9222 6679 9274
rect 6679 9222 6725 9274
rect 6429 9220 6485 9222
rect 6509 9220 6565 9222
rect 6589 9220 6645 9222
rect 6669 9220 6725 9222
rect 6429 8186 6485 8188
rect 6509 8186 6565 8188
rect 6589 8186 6645 8188
rect 6669 8186 6725 8188
rect 6429 8134 6475 8186
rect 6475 8134 6485 8186
rect 6509 8134 6539 8186
rect 6539 8134 6551 8186
rect 6551 8134 6565 8186
rect 6589 8134 6603 8186
rect 6603 8134 6615 8186
rect 6615 8134 6645 8186
rect 6669 8134 6679 8186
rect 6679 8134 6725 8186
rect 6429 8132 6485 8134
rect 6509 8132 6565 8134
rect 6589 8132 6645 8134
rect 6669 8132 6725 8134
rect 6429 7098 6485 7100
rect 6509 7098 6565 7100
rect 6589 7098 6645 7100
rect 6669 7098 6725 7100
rect 6429 7046 6475 7098
rect 6475 7046 6485 7098
rect 6509 7046 6539 7098
rect 6539 7046 6551 7098
rect 6551 7046 6565 7098
rect 6589 7046 6603 7098
rect 6603 7046 6615 7098
rect 6615 7046 6645 7098
rect 6669 7046 6679 7098
rect 6679 7046 6725 7098
rect 6429 7044 6485 7046
rect 6509 7044 6565 7046
rect 6589 7044 6645 7046
rect 6669 7044 6725 7046
rect 6429 6010 6485 6012
rect 6509 6010 6565 6012
rect 6589 6010 6645 6012
rect 6669 6010 6725 6012
rect 6429 5958 6475 6010
rect 6475 5958 6485 6010
rect 6509 5958 6539 6010
rect 6539 5958 6551 6010
rect 6551 5958 6565 6010
rect 6589 5958 6603 6010
rect 6603 5958 6615 6010
rect 6615 5958 6645 6010
rect 6669 5958 6679 6010
rect 6679 5958 6725 6010
rect 6429 5956 6485 5958
rect 6509 5956 6565 5958
rect 6589 5956 6645 5958
rect 6669 5956 6725 5958
rect 6429 4922 6485 4924
rect 6509 4922 6565 4924
rect 6589 4922 6645 4924
rect 6669 4922 6725 4924
rect 6429 4870 6475 4922
rect 6475 4870 6485 4922
rect 6509 4870 6539 4922
rect 6539 4870 6551 4922
rect 6551 4870 6565 4922
rect 6589 4870 6603 4922
rect 6603 4870 6615 4922
rect 6615 4870 6645 4922
rect 6669 4870 6679 4922
rect 6679 4870 6725 4922
rect 6429 4868 6485 4870
rect 6509 4868 6565 4870
rect 6589 4868 6645 4870
rect 6669 4868 6725 4870
rect 6429 3834 6485 3836
rect 6509 3834 6565 3836
rect 6589 3834 6645 3836
rect 6669 3834 6725 3836
rect 6429 3782 6475 3834
rect 6475 3782 6485 3834
rect 6509 3782 6539 3834
rect 6539 3782 6551 3834
rect 6551 3782 6565 3834
rect 6589 3782 6603 3834
rect 6603 3782 6615 3834
rect 6615 3782 6645 3834
rect 6669 3782 6679 3834
rect 6679 3782 6725 3834
rect 6429 3780 6485 3782
rect 6509 3780 6565 3782
rect 6589 3780 6645 3782
rect 6669 3780 6725 3782
rect 938 3476 940 3496
rect 940 3476 992 3496
rect 992 3476 994 3496
rect 938 3440 994 3476
rect 11902 13082 11958 13084
rect 11982 13082 12038 13084
rect 12062 13082 12118 13084
rect 12142 13082 12198 13084
rect 11902 13030 11948 13082
rect 11948 13030 11958 13082
rect 11982 13030 12012 13082
rect 12012 13030 12024 13082
rect 12024 13030 12038 13082
rect 12062 13030 12076 13082
rect 12076 13030 12088 13082
rect 12088 13030 12118 13082
rect 12142 13030 12152 13082
rect 12152 13030 12198 13082
rect 11902 13028 11958 13030
rect 11982 13028 12038 13030
rect 12062 13028 12118 13030
rect 12142 13028 12198 13030
rect 11902 11994 11958 11996
rect 11982 11994 12038 11996
rect 12062 11994 12118 11996
rect 12142 11994 12198 11996
rect 11902 11942 11948 11994
rect 11948 11942 11958 11994
rect 11982 11942 12012 11994
rect 12012 11942 12024 11994
rect 12024 11942 12038 11994
rect 12062 11942 12076 11994
rect 12076 11942 12088 11994
rect 12088 11942 12118 11994
rect 12142 11942 12152 11994
rect 12152 11942 12198 11994
rect 11902 11940 11958 11942
rect 11982 11940 12038 11942
rect 12062 11940 12118 11942
rect 12142 11940 12198 11942
rect 11902 10906 11958 10908
rect 11982 10906 12038 10908
rect 12062 10906 12118 10908
rect 12142 10906 12198 10908
rect 11902 10854 11948 10906
rect 11948 10854 11958 10906
rect 11982 10854 12012 10906
rect 12012 10854 12024 10906
rect 12024 10854 12038 10906
rect 12062 10854 12076 10906
rect 12076 10854 12088 10906
rect 12088 10854 12118 10906
rect 12142 10854 12152 10906
rect 12152 10854 12198 10906
rect 11902 10852 11958 10854
rect 11982 10852 12038 10854
rect 12062 10852 12118 10854
rect 12142 10852 12198 10854
rect 12806 9968 12862 10024
rect 11902 9818 11958 9820
rect 11982 9818 12038 9820
rect 12062 9818 12118 9820
rect 12142 9818 12198 9820
rect 11902 9766 11948 9818
rect 11948 9766 11958 9818
rect 11982 9766 12012 9818
rect 12012 9766 12024 9818
rect 12024 9766 12038 9818
rect 12062 9766 12076 9818
rect 12076 9766 12088 9818
rect 12088 9766 12118 9818
rect 12142 9766 12152 9818
rect 12152 9766 12198 9818
rect 11902 9764 11958 9766
rect 11982 9764 12038 9766
rect 12062 9764 12118 9766
rect 12142 9764 12198 9766
rect 11902 8730 11958 8732
rect 11982 8730 12038 8732
rect 12062 8730 12118 8732
rect 12142 8730 12198 8732
rect 11902 8678 11948 8730
rect 11948 8678 11958 8730
rect 11982 8678 12012 8730
rect 12012 8678 12024 8730
rect 12024 8678 12038 8730
rect 12062 8678 12076 8730
rect 12076 8678 12088 8730
rect 12088 8678 12118 8730
rect 12142 8678 12152 8730
rect 12152 8678 12198 8730
rect 11902 8676 11958 8678
rect 11982 8676 12038 8678
rect 12062 8676 12118 8678
rect 12142 8676 12198 8678
rect 16302 14456 16358 14512
rect 11902 7642 11958 7644
rect 11982 7642 12038 7644
rect 12062 7642 12118 7644
rect 12142 7642 12198 7644
rect 11902 7590 11948 7642
rect 11948 7590 11958 7642
rect 11982 7590 12012 7642
rect 12012 7590 12024 7642
rect 12024 7590 12038 7642
rect 12062 7590 12076 7642
rect 12076 7590 12088 7642
rect 12088 7590 12118 7642
rect 12142 7590 12152 7642
rect 12152 7590 12198 7642
rect 11902 7588 11958 7590
rect 11982 7588 12038 7590
rect 12062 7588 12118 7590
rect 12142 7588 12198 7590
rect 11902 6554 11958 6556
rect 11982 6554 12038 6556
rect 12062 6554 12118 6556
rect 12142 6554 12198 6556
rect 11902 6502 11948 6554
rect 11948 6502 11958 6554
rect 11982 6502 12012 6554
rect 12012 6502 12024 6554
rect 12024 6502 12038 6554
rect 12062 6502 12076 6554
rect 12076 6502 12088 6554
rect 12088 6502 12118 6554
rect 12142 6502 12152 6554
rect 12152 6502 12198 6554
rect 11902 6500 11958 6502
rect 11982 6500 12038 6502
rect 12062 6500 12118 6502
rect 12142 6500 12198 6502
rect 12070 6316 12126 6352
rect 12070 6296 12072 6316
rect 12072 6296 12124 6316
rect 12124 6296 12126 6316
rect 11902 5466 11958 5468
rect 11982 5466 12038 5468
rect 12062 5466 12118 5468
rect 12142 5466 12198 5468
rect 11902 5414 11948 5466
rect 11948 5414 11958 5466
rect 11982 5414 12012 5466
rect 12012 5414 12024 5466
rect 12024 5414 12038 5466
rect 12062 5414 12076 5466
rect 12076 5414 12088 5466
rect 12088 5414 12118 5466
rect 12142 5414 12152 5466
rect 12152 5414 12198 5466
rect 11902 5412 11958 5414
rect 11982 5412 12038 5414
rect 12062 5412 12118 5414
rect 12142 5412 12198 5414
rect 11902 4378 11958 4380
rect 11982 4378 12038 4380
rect 12062 4378 12118 4380
rect 12142 4378 12198 4380
rect 11902 4326 11948 4378
rect 11948 4326 11958 4378
rect 11982 4326 12012 4378
rect 12012 4326 12024 4378
rect 12024 4326 12038 4378
rect 12062 4326 12076 4378
rect 12076 4326 12088 4378
rect 12088 4326 12118 4378
rect 12142 4326 12152 4378
rect 12152 4326 12198 4378
rect 11902 4324 11958 4326
rect 11982 4324 12038 4326
rect 12062 4324 12118 4326
rect 12142 4324 12198 4326
rect 11902 3290 11958 3292
rect 11982 3290 12038 3292
rect 12062 3290 12118 3292
rect 12142 3290 12198 3292
rect 11902 3238 11948 3290
rect 11948 3238 11958 3290
rect 11982 3238 12012 3290
rect 12012 3238 12024 3290
rect 12024 3238 12038 3290
rect 12062 3238 12076 3290
rect 12076 3238 12088 3290
rect 12088 3238 12118 3290
rect 12142 3238 12152 3290
rect 12152 3238 12198 3290
rect 11902 3236 11958 3238
rect 11982 3236 12038 3238
rect 12062 3236 12118 3238
rect 12142 3236 12198 3238
rect 6429 2746 6485 2748
rect 6509 2746 6565 2748
rect 6589 2746 6645 2748
rect 6669 2746 6725 2748
rect 6429 2694 6475 2746
rect 6475 2694 6485 2746
rect 6509 2694 6539 2746
rect 6539 2694 6551 2746
rect 6551 2694 6565 2746
rect 6589 2694 6603 2746
rect 6603 2694 6615 2746
rect 6615 2694 6645 2746
rect 6669 2694 6679 2746
rect 6679 2694 6725 2746
rect 6429 2692 6485 2694
rect 6509 2692 6565 2694
rect 6589 2692 6645 2694
rect 6669 2692 6725 2694
rect 14830 7928 14886 7984
rect 13634 6160 13690 6216
rect 17376 16890 17432 16892
rect 17456 16890 17512 16892
rect 17536 16890 17592 16892
rect 17616 16890 17672 16892
rect 17376 16838 17422 16890
rect 17422 16838 17432 16890
rect 17456 16838 17486 16890
rect 17486 16838 17498 16890
rect 17498 16838 17512 16890
rect 17536 16838 17550 16890
rect 17550 16838 17562 16890
rect 17562 16838 17592 16890
rect 17616 16838 17626 16890
rect 17626 16838 17672 16890
rect 17376 16836 17432 16838
rect 17456 16836 17512 16838
rect 17536 16836 17592 16838
rect 17616 16836 17672 16838
rect 22849 16346 22905 16348
rect 22929 16346 22985 16348
rect 23009 16346 23065 16348
rect 23089 16346 23145 16348
rect 22849 16294 22895 16346
rect 22895 16294 22905 16346
rect 22929 16294 22959 16346
rect 22959 16294 22971 16346
rect 22971 16294 22985 16346
rect 23009 16294 23023 16346
rect 23023 16294 23035 16346
rect 23035 16294 23065 16346
rect 23089 16294 23099 16346
rect 23099 16294 23145 16346
rect 22849 16292 22905 16294
rect 22929 16292 22985 16294
rect 23009 16292 23065 16294
rect 23089 16292 23145 16294
rect 17376 15802 17432 15804
rect 17456 15802 17512 15804
rect 17536 15802 17592 15804
rect 17616 15802 17672 15804
rect 17376 15750 17422 15802
rect 17422 15750 17432 15802
rect 17456 15750 17486 15802
rect 17486 15750 17498 15802
rect 17498 15750 17512 15802
rect 17536 15750 17550 15802
rect 17550 15750 17562 15802
rect 17562 15750 17592 15802
rect 17616 15750 17626 15802
rect 17626 15750 17672 15802
rect 17376 15748 17432 15750
rect 17456 15748 17512 15750
rect 17536 15748 17592 15750
rect 17616 15748 17672 15750
rect 22849 15258 22905 15260
rect 22929 15258 22985 15260
rect 23009 15258 23065 15260
rect 23089 15258 23145 15260
rect 22849 15206 22895 15258
rect 22895 15206 22905 15258
rect 22929 15206 22959 15258
rect 22959 15206 22971 15258
rect 22971 15206 22985 15258
rect 23009 15206 23023 15258
rect 23023 15206 23035 15258
rect 23035 15206 23065 15258
rect 23089 15206 23099 15258
rect 23099 15206 23145 15258
rect 22849 15204 22905 15206
rect 22929 15204 22985 15206
rect 23009 15204 23065 15206
rect 23089 15204 23145 15206
rect 28323 16890 28379 16892
rect 28403 16890 28459 16892
rect 28483 16890 28539 16892
rect 28563 16890 28619 16892
rect 28323 16838 28369 16890
rect 28369 16838 28379 16890
rect 28403 16838 28433 16890
rect 28433 16838 28445 16890
rect 28445 16838 28459 16890
rect 28483 16838 28497 16890
rect 28497 16838 28509 16890
rect 28509 16838 28539 16890
rect 28563 16838 28573 16890
rect 28573 16838 28619 16890
rect 28323 16836 28379 16838
rect 28403 16836 28459 16838
rect 28483 16836 28539 16838
rect 28563 16836 28619 16838
rect 17376 14714 17432 14716
rect 17456 14714 17512 14716
rect 17536 14714 17592 14716
rect 17616 14714 17672 14716
rect 17376 14662 17422 14714
rect 17422 14662 17432 14714
rect 17456 14662 17486 14714
rect 17486 14662 17498 14714
rect 17498 14662 17512 14714
rect 17536 14662 17550 14714
rect 17550 14662 17562 14714
rect 17562 14662 17592 14714
rect 17616 14662 17626 14714
rect 17626 14662 17672 14714
rect 17376 14660 17432 14662
rect 17456 14660 17512 14662
rect 17536 14660 17592 14662
rect 17616 14660 17672 14662
rect 17376 13626 17432 13628
rect 17456 13626 17512 13628
rect 17536 13626 17592 13628
rect 17616 13626 17672 13628
rect 17376 13574 17422 13626
rect 17422 13574 17432 13626
rect 17456 13574 17486 13626
rect 17486 13574 17498 13626
rect 17498 13574 17512 13626
rect 17536 13574 17550 13626
rect 17550 13574 17562 13626
rect 17562 13574 17592 13626
rect 17616 13574 17626 13626
rect 17626 13574 17672 13626
rect 17376 13572 17432 13574
rect 17456 13572 17512 13574
rect 17536 13572 17592 13574
rect 17616 13572 17672 13574
rect 17376 12538 17432 12540
rect 17456 12538 17512 12540
rect 17536 12538 17592 12540
rect 17616 12538 17672 12540
rect 17376 12486 17422 12538
rect 17422 12486 17432 12538
rect 17456 12486 17486 12538
rect 17486 12486 17498 12538
rect 17498 12486 17512 12538
rect 17536 12486 17550 12538
rect 17550 12486 17562 12538
rect 17562 12486 17592 12538
rect 17616 12486 17626 12538
rect 17626 12486 17672 12538
rect 17376 12484 17432 12486
rect 17456 12484 17512 12486
rect 17536 12484 17592 12486
rect 17616 12484 17672 12486
rect 17376 11450 17432 11452
rect 17456 11450 17512 11452
rect 17536 11450 17592 11452
rect 17616 11450 17672 11452
rect 17376 11398 17422 11450
rect 17422 11398 17432 11450
rect 17456 11398 17486 11450
rect 17486 11398 17498 11450
rect 17498 11398 17512 11450
rect 17536 11398 17550 11450
rect 17550 11398 17562 11450
rect 17562 11398 17592 11450
rect 17616 11398 17626 11450
rect 17626 11398 17672 11450
rect 17376 11396 17432 11398
rect 17456 11396 17512 11398
rect 17536 11396 17592 11398
rect 17616 11396 17672 11398
rect 17376 10362 17432 10364
rect 17456 10362 17512 10364
rect 17536 10362 17592 10364
rect 17616 10362 17672 10364
rect 17376 10310 17422 10362
rect 17422 10310 17432 10362
rect 17456 10310 17486 10362
rect 17486 10310 17498 10362
rect 17498 10310 17512 10362
rect 17536 10310 17550 10362
rect 17550 10310 17562 10362
rect 17562 10310 17592 10362
rect 17616 10310 17626 10362
rect 17626 10310 17672 10362
rect 17376 10308 17432 10310
rect 17456 10308 17512 10310
rect 17536 10308 17592 10310
rect 17616 10308 17672 10310
rect 17376 9274 17432 9276
rect 17456 9274 17512 9276
rect 17536 9274 17592 9276
rect 17616 9274 17672 9276
rect 17376 9222 17422 9274
rect 17422 9222 17432 9274
rect 17456 9222 17486 9274
rect 17486 9222 17498 9274
rect 17498 9222 17512 9274
rect 17536 9222 17550 9274
rect 17550 9222 17562 9274
rect 17562 9222 17592 9274
rect 17616 9222 17626 9274
rect 17626 9222 17672 9274
rect 17376 9220 17432 9222
rect 17456 9220 17512 9222
rect 17536 9220 17592 9222
rect 17616 9220 17672 9222
rect 17376 8186 17432 8188
rect 17456 8186 17512 8188
rect 17536 8186 17592 8188
rect 17616 8186 17672 8188
rect 17376 8134 17422 8186
rect 17422 8134 17432 8186
rect 17456 8134 17486 8186
rect 17486 8134 17498 8186
rect 17498 8134 17512 8186
rect 17536 8134 17550 8186
rect 17550 8134 17562 8186
rect 17562 8134 17592 8186
rect 17616 8134 17626 8186
rect 17626 8134 17672 8186
rect 17376 8132 17432 8134
rect 17456 8132 17512 8134
rect 17536 8132 17592 8134
rect 17616 8132 17672 8134
rect 17376 7098 17432 7100
rect 17456 7098 17512 7100
rect 17536 7098 17592 7100
rect 17616 7098 17672 7100
rect 17376 7046 17422 7098
rect 17422 7046 17432 7098
rect 17456 7046 17486 7098
rect 17486 7046 17498 7098
rect 17498 7046 17512 7098
rect 17536 7046 17550 7098
rect 17550 7046 17562 7098
rect 17562 7046 17592 7098
rect 17616 7046 17626 7098
rect 17626 7046 17672 7098
rect 17376 7044 17432 7046
rect 17456 7044 17512 7046
rect 17536 7044 17592 7046
rect 17616 7044 17672 7046
rect 17774 6296 17830 6352
rect 17376 6010 17432 6012
rect 17456 6010 17512 6012
rect 17536 6010 17592 6012
rect 17616 6010 17672 6012
rect 17376 5958 17422 6010
rect 17422 5958 17432 6010
rect 17456 5958 17486 6010
rect 17486 5958 17498 6010
rect 17498 5958 17512 6010
rect 17536 5958 17550 6010
rect 17550 5958 17562 6010
rect 17562 5958 17592 6010
rect 17616 5958 17626 6010
rect 17626 5958 17672 6010
rect 17376 5956 17432 5958
rect 17456 5956 17512 5958
rect 17536 5956 17592 5958
rect 17616 5956 17672 5958
rect 17376 4922 17432 4924
rect 17456 4922 17512 4924
rect 17536 4922 17592 4924
rect 17616 4922 17672 4924
rect 17376 4870 17422 4922
rect 17422 4870 17432 4922
rect 17456 4870 17486 4922
rect 17486 4870 17498 4922
rect 17498 4870 17512 4922
rect 17536 4870 17550 4922
rect 17550 4870 17562 4922
rect 17562 4870 17592 4922
rect 17616 4870 17626 4922
rect 17626 4870 17672 4922
rect 17376 4868 17432 4870
rect 17456 4868 17512 4870
rect 17536 4868 17592 4870
rect 17616 4868 17672 4870
rect 22849 14170 22905 14172
rect 22929 14170 22985 14172
rect 23009 14170 23065 14172
rect 23089 14170 23145 14172
rect 22849 14118 22895 14170
rect 22895 14118 22905 14170
rect 22929 14118 22959 14170
rect 22959 14118 22971 14170
rect 22971 14118 22985 14170
rect 23009 14118 23023 14170
rect 23023 14118 23035 14170
rect 23035 14118 23065 14170
rect 23089 14118 23099 14170
rect 23099 14118 23145 14170
rect 22849 14116 22905 14118
rect 22929 14116 22985 14118
rect 23009 14116 23065 14118
rect 23089 14116 23145 14118
rect 22849 13082 22905 13084
rect 22929 13082 22985 13084
rect 23009 13082 23065 13084
rect 23089 13082 23145 13084
rect 22849 13030 22895 13082
rect 22895 13030 22905 13082
rect 22929 13030 22959 13082
rect 22959 13030 22971 13082
rect 22971 13030 22985 13082
rect 23009 13030 23023 13082
rect 23023 13030 23035 13082
rect 23035 13030 23065 13082
rect 23089 13030 23099 13082
rect 23099 13030 23145 13082
rect 22849 13028 22905 13030
rect 22929 13028 22985 13030
rect 23009 13028 23065 13030
rect 23089 13028 23145 13030
rect 24766 12824 24822 12880
rect 22849 11994 22905 11996
rect 22929 11994 22985 11996
rect 23009 11994 23065 11996
rect 23089 11994 23145 11996
rect 22849 11942 22895 11994
rect 22895 11942 22905 11994
rect 22929 11942 22959 11994
rect 22959 11942 22971 11994
rect 22971 11942 22985 11994
rect 23009 11942 23023 11994
rect 23023 11942 23035 11994
rect 23035 11942 23065 11994
rect 23089 11942 23099 11994
rect 23099 11942 23145 11994
rect 22849 11940 22905 11942
rect 22929 11940 22985 11942
rect 23009 11940 23065 11942
rect 23089 11940 23145 11942
rect 22849 10906 22905 10908
rect 22929 10906 22985 10908
rect 23009 10906 23065 10908
rect 23089 10906 23145 10908
rect 22849 10854 22895 10906
rect 22895 10854 22905 10906
rect 22929 10854 22959 10906
rect 22959 10854 22971 10906
rect 22971 10854 22985 10906
rect 23009 10854 23023 10906
rect 23023 10854 23035 10906
rect 23035 10854 23065 10906
rect 23089 10854 23099 10906
rect 23099 10854 23145 10906
rect 22849 10852 22905 10854
rect 22929 10852 22985 10854
rect 23009 10852 23065 10854
rect 23089 10852 23145 10854
rect 22849 9818 22905 9820
rect 22929 9818 22985 9820
rect 23009 9818 23065 9820
rect 23089 9818 23145 9820
rect 22849 9766 22895 9818
rect 22895 9766 22905 9818
rect 22929 9766 22959 9818
rect 22959 9766 22971 9818
rect 22971 9766 22985 9818
rect 23009 9766 23023 9818
rect 23023 9766 23035 9818
rect 23035 9766 23065 9818
rect 23089 9766 23099 9818
rect 23099 9766 23145 9818
rect 22849 9764 22905 9766
rect 22929 9764 22985 9766
rect 23009 9764 23065 9766
rect 23089 9764 23145 9766
rect 17376 3834 17432 3836
rect 17456 3834 17512 3836
rect 17536 3834 17592 3836
rect 17616 3834 17672 3836
rect 17376 3782 17422 3834
rect 17422 3782 17432 3834
rect 17456 3782 17486 3834
rect 17486 3782 17498 3834
rect 17498 3782 17512 3834
rect 17536 3782 17550 3834
rect 17550 3782 17562 3834
rect 17562 3782 17592 3834
rect 17616 3782 17626 3834
rect 17626 3782 17672 3834
rect 17376 3780 17432 3782
rect 17456 3780 17512 3782
rect 17536 3780 17592 3782
rect 17616 3780 17672 3782
rect 938 1400 994 1456
rect 11902 2202 11958 2204
rect 11982 2202 12038 2204
rect 12062 2202 12118 2204
rect 12142 2202 12198 2204
rect 11902 2150 11948 2202
rect 11948 2150 11958 2202
rect 11982 2150 12012 2202
rect 12012 2150 12024 2202
rect 12024 2150 12038 2202
rect 12062 2150 12076 2202
rect 12076 2150 12088 2202
rect 12088 2150 12118 2202
rect 12142 2150 12152 2202
rect 12152 2150 12198 2202
rect 11902 2148 11958 2150
rect 11982 2148 12038 2150
rect 12062 2148 12118 2150
rect 12142 2148 12198 2150
rect 22849 8730 22905 8732
rect 22929 8730 22985 8732
rect 23009 8730 23065 8732
rect 23089 8730 23145 8732
rect 22849 8678 22895 8730
rect 22895 8678 22905 8730
rect 22929 8678 22959 8730
rect 22959 8678 22971 8730
rect 22971 8678 22985 8730
rect 23009 8678 23023 8730
rect 23023 8678 23035 8730
rect 23035 8678 23065 8730
rect 23089 8678 23099 8730
rect 23099 8678 23145 8730
rect 22849 8676 22905 8678
rect 22929 8676 22985 8678
rect 23009 8676 23065 8678
rect 23089 8676 23145 8678
rect 22849 7642 22905 7644
rect 22929 7642 22985 7644
rect 23009 7642 23065 7644
rect 23089 7642 23145 7644
rect 22849 7590 22895 7642
rect 22895 7590 22905 7642
rect 22929 7590 22959 7642
rect 22959 7590 22971 7642
rect 22971 7590 22985 7642
rect 23009 7590 23023 7642
rect 23023 7590 23035 7642
rect 23035 7590 23065 7642
rect 23089 7590 23099 7642
rect 23099 7590 23145 7642
rect 22849 7588 22905 7590
rect 22929 7588 22985 7590
rect 23009 7588 23065 7590
rect 23089 7588 23145 7590
rect 22849 6554 22905 6556
rect 22929 6554 22985 6556
rect 23009 6554 23065 6556
rect 23089 6554 23145 6556
rect 22849 6502 22895 6554
rect 22895 6502 22905 6554
rect 22929 6502 22959 6554
rect 22959 6502 22971 6554
rect 22971 6502 22985 6554
rect 23009 6502 23023 6554
rect 23023 6502 23035 6554
rect 23035 6502 23065 6554
rect 23089 6502 23099 6554
rect 23099 6502 23145 6554
rect 22849 6500 22905 6502
rect 22929 6500 22985 6502
rect 23009 6500 23065 6502
rect 23089 6500 23145 6502
rect 22849 5466 22905 5468
rect 22929 5466 22985 5468
rect 23009 5466 23065 5468
rect 23089 5466 23145 5468
rect 22849 5414 22895 5466
rect 22895 5414 22905 5466
rect 22929 5414 22959 5466
rect 22959 5414 22971 5466
rect 22971 5414 22985 5466
rect 23009 5414 23023 5466
rect 23023 5414 23035 5466
rect 23035 5414 23065 5466
rect 23089 5414 23099 5466
rect 23099 5414 23145 5466
rect 22849 5412 22905 5414
rect 22929 5412 22985 5414
rect 23009 5412 23065 5414
rect 23089 5412 23145 5414
rect 22849 4378 22905 4380
rect 22929 4378 22985 4380
rect 23009 4378 23065 4380
rect 23089 4378 23145 4380
rect 22849 4326 22895 4378
rect 22895 4326 22905 4378
rect 22929 4326 22959 4378
rect 22959 4326 22971 4378
rect 22971 4326 22985 4378
rect 23009 4326 23023 4378
rect 23023 4326 23035 4378
rect 23035 4326 23065 4378
rect 23089 4326 23099 4378
rect 23099 4326 23145 4378
rect 22849 4324 22905 4326
rect 22929 4324 22985 4326
rect 23009 4324 23065 4326
rect 23089 4324 23145 4326
rect 28323 15802 28379 15804
rect 28403 15802 28459 15804
rect 28483 15802 28539 15804
rect 28563 15802 28619 15804
rect 28323 15750 28369 15802
rect 28369 15750 28379 15802
rect 28403 15750 28433 15802
rect 28433 15750 28445 15802
rect 28445 15750 28459 15802
rect 28483 15750 28497 15802
rect 28497 15750 28509 15802
rect 28509 15750 28539 15802
rect 28563 15750 28573 15802
rect 28573 15750 28619 15802
rect 28323 15748 28379 15750
rect 28403 15748 28459 15750
rect 28483 15748 28539 15750
rect 28563 15748 28619 15750
rect 28323 14714 28379 14716
rect 28403 14714 28459 14716
rect 28483 14714 28539 14716
rect 28563 14714 28619 14716
rect 28323 14662 28369 14714
rect 28369 14662 28379 14714
rect 28403 14662 28433 14714
rect 28433 14662 28445 14714
rect 28445 14662 28459 14714
rect 28483 14662 28497 14714
rect 28497 14662 28509 14714
rect 28509 14662 28539 14714
rect 28563 14662 28573 14714
rect 28573 14662 28619 14714
rect 28323 14660 28379 14662
rect 28403 14660 28459 14662
rect 28483 14660 28539 14662
rect 28563 14660 28619 14662
rect 28323 13626 28379 13628
rect 28403 13626 28459 13628
rect 28483 13626 28539 13628
rect 28563 13626 28619 13628
rect 28323 13574 28369 13626
rect 28369 13574 28379 13626
rect 28403 13574 28433 13626
rect 28433 13574 28445 13626
rect 28445 13574 28459 13626
rect 28483 13574 28497 13626
rect 28497 13574 28509 13626
rect 28509 13574 28539 13626
rect 28563 13574 28573 13626
rect 28573 13574 28619 13626
rect 28323 13572 28379 13574
rect 28403 13572 28459 13574
rect 28483 13572 28539 13574
rect 28563 13572 28619 13574
rect 28323 12538 28379 12540
rect 28403 12538 28459 12540
rect 28483 12538 28539 12540
rect 28563 12538 28619 12540
rect 28323 12486 28369 12538
rect 28369 12486 28379 12538
rect 28403 12486 28433 12538
rect 28433 12486 28445 12538
rect 28445 12486 28459 12538
rect 28483 12486 28497 12538
rect 28497 12486 28509 12538
rect 28509 12486 28539 12538
rect 28563 12486 28573 12538
rect 28573 12486 28619 12538
rect 28323 12484 28379 12486
rect 28403 12484 28459 12486
rect 28483 12484 28539 12486
rect 28563 12484 28619 12486
rect 33796 16346 33852 16348
rect 33876 16346 33932 16348
rect 33956 16346 34012 16348
rect 34036 16346 34092 16348
rect 33796 16294 33842 16346
rect 33842 16294 33852 16346
rect 33876 16294 33906 16346
rect 33906 16294 33918 16346
rect 33918 16294 33932 16346
rect 33956 16294 33970 16346
rect 33970 16294 33982 16346
rect 33982 16294 34012 16346
rect 34036 16294 34046 16346
rect 34046 16294 34092 16346
rect 33796 16292 33852 16294
rect 33876 16292 33932 16294
rect 33956 16292 34012 16294
rect 34036 16292 34092 16294
rect 28323 11450 28379 11452
rect 28403 11450 28459 11452
rect 28483 11450 28539 11452
rect 28563 11450 28619 11452
rect 28323 11398 28369 11450
rect 28369 11398 28379 11450
rect 28403 11398 28433 11450
rect 28433 11398 28445 11450
rect 28445 11398 28459 11450
rect 28483 11398 28497 11450
rect 28497 11398 28509 11450
rect 28509 11398 28539 11450
rect 28563 11398 28573 11450
rect 28573 11398 28619 11450
rect 28323 11396 28379 11398
rect 28403 11396 28459 11398
rect 28483 11396 28539 11398
rect 28563 11396 28619 11398
rect 33796 15258 33852 15260
rect 33876 15258 33932 15260
rect 33956 15258 34012 15260
rect 34036 15258 34092 15260
rect 33796 15206 33842 15258
rect 33842 15206 33852 15258
rect 33876 15206 33906 15258
rect 33906 15206 33918 15258
rect 33918 15206 33932 15258
rect 33956 15206 33970 15258
rect 33970 15206 33982 15258
rect 33982 15206 34012 15258
rect 34036 15206 34046 15258
rect 34046 15206 34092 15258
rect 33796 15204 33852 15206
rect 33876 15204 33932 15206
rect 33956 15204 34012 15206
rect 34036 15204 34092 15206
rect 32586 14884 32642 14920
rect 32586 14864 32588 14884
rect 32588 14864 32640 14884
rect 32640 14864 32642 14884
rect 31574 12844 31630 12880
rect 31574 12824 31576 12844
rect 31576 12824 31628 12844
rect 31628 12824 31630 12844
rect 32494 13252 32550 13288
rect 32494 13232 32496 13252
rect 32496 13232 32548 13252
rect 32548 13232 32550 13252
rect 32586 12688 32642 12744
rect 28323 10362 28379 10364
rect 28403 10362 28459 10364
rect 28483 10362 28539 10364
rect 28563 10362 28619 10364
rect 28323 10310 28369 10362
rect 28369 10310 28379 10362
rect 28403 10310 28433 10362
rect 28433 10310 28445 10362
rect 28445 10310 28459 10362
rect 28483 10310 28497 10362
rect 28497 10310 28509 10362
rect 28509 10310 28539 10362
rect 28563 10310 28573 10362
rect 28573 10310 28619 10362
rect 28323 10308 28379 10310
rect 28403 10308 28459 10310
rect 28483 10308 28539 10310
rect 28563 10308 28619 10310
rect 28323 9274 28379 9276
rect 28403 9274 28459 9276
rect 28483 9274 28539 9276
rect 28563 9274 28619 9276
rect 28323 9222 28369 9274
rect 28369 9222 28379 9274
rect 28403 9222 28433 9274
rect 28433 9222 28445 9274
rect 28445 9222 28459 9274
rect 28483 9222 28497 9274
rect 28497 9222 28509 9274
rect 28509 9222 28539 9274
rect 28563 9222 28573 9274
rect 28573 9222 28619 9274
rect 28323 9220 28379 9222
rect 28403 9220 28459 9222
rect 28483 9220 28539 9222
rect 28563 9220 28619 9222
rect 25318 6196 25320 6216
rect 25320 6196 25372 6216
rect 25372 6196 25374 6216
rect 25318 6160 25374 6196
rect 27710 8900 27766 8936
rect 27710 8880 27712 8900
rect 27712 8880 27764 8900
rect 27764 8880 27766 8900
rect 29826 10004 29828 10024
rect 29828 10004 29880 10024
rect 29880 10004 29882 10024
rect 29826 9968 29882 10004
rect 33966 14864 34022 14920
rect 33796 14170 33852 14172
rect 33876 14170 33932 14172
rect 33956 14170 34012 14172
rect 34036 14170 34092 14172
rect 33796 14118 33842 14170
rect 33842 14118 33852 14170
rect 33876 14118 33906 14170
rect 33906 14118 33918 14170
rect 33918 14118 33932 14170
rect 33956 14118 33970 14170
rect 33970 14118 33982 14170
rect 33982 14118 34012 14170
rect 34036 14118 34046 14170
rect 34046 14118 34092 14170
rect 33796 14116 33852 14118
rect 33876 14116 33932 14118
rect 33956 14116 34012 14118
rect 34036 14116 34092 14118
rect 33506 12824 33562 12880
rect 33796 13082 33852 13084
rect 33876 13082 33932 13084
rect 33956 13082 34012 13084
rect 34036 13082 34092 13084
rect 33796 13030 33842 13082
rect 33842 13030 33852 13082
rect 33876 13030 33906 13082
rect 33906 13030 33918 13082
rect 33918 13030 33932 13082
rect 33956 13030 33970 13082
rect 33970 13030 33982 13082
rect 33982 13030 34012 13082
rect 34036 13030 34046 13082
rect 34046 13030 34092 13082
rect 33796 13028 33852 13030
rect 33876 13028 33932 13030
rect 33956 13028 34012 13030
rect 34036 13028 34092 13030
rect 33796 11994 33852 11996
rect 33876 11994 33932 11996
rect 33956 11994 34012 11996
rect 34036 11994 34092 11996
rect 33796 11942 33842 11994
rect 33842 11942 33852 11994
rect 33876 11942 33906 11994
rect 33906 11942 33918 11994
rect 33918 11942 33932 11994
rect 33956 11942 33970 11994
rect 33970 11942 33982 11994
rect 33982 11942 34012 11994
rect 34036 11942 34046 11994
rect 34046 11942 34092 11994
rect 33796 11940 33852 11942
rect 33876 11940 33932 11942
rect 33956 11940 34012 11942
rect 34036 11940 34092 11942
rect 27618 7948 27674 7984
rect 27618 7928 27620 7948
rect 27620 7928 27672 7948
rect 27672 7928 27674 7948
rect 28323 8186 28379 8188
rect 28403 8186 28459 8188
rect 28483 8186 28539 8188
rect 28563 8186 28619 8188
rect 28323 8134 28369 8186
rect 28369 8134 28379 8186
rect 28403 8134 28433 8186
rect 28433 8134 28445 8186
rect 28445 8134 28459 8186
rect 28483 8134 28497 8186
rect 28497 8134 28509 8186
rect 28509 8134 28539 8186
rect 28563 8134 28573 8186
rect 28573 8134 28619 8186
rect 28323 8132 28379 8134
rect 28403 8132 28459 8134
rect 28483 8132 28539 8134
rect 28563 8132 28619 8134
rect 28323 7098 28379 7100
rect 28403 7098 28459 7100
rect 28483 7098 28539 7100
rect 28563 7098 28619 7100
rect 28323 7046 28369 7098
rect 28369 7046 28379 7098
rect 28403 7046 28433 7098
rect 28433 7046 28445 7098
rect 28445 7046 28459 7098
rect 28483 7046 28497 7098
rect 28497 7046 28509 7098
rect 28509 7046 28539 7098
rect 28563 7046 28573 7098
rect 28573 7046 28619 7098
rect 28323 7044 28379 7046
rect 28403 7044 28459 7046
rect 28483 7044 28539 7046
rect 28563 7044 28619 7046
rect 22849 3290 22905 3292
rect 22929 3290 22985 3292
rect 23009 3290 23065 3292
rect 23089 3290 23145 3292
rect 22849 3238 22895 3290
rect 22895 3238 22905 3290
rect 22929 3238 22959 3290
rect 22959 3238 22971 3290
rect 22971 3238 22985 3290
rect 23009 3238 23023 3290
rect 23023 3238 23035 3290
rect 23035 3238 23065 3290
rect 23089 3238 23099 3290
rect 23099 3238 23145 3290
rect 22849 3236 22905 3238
rect 22929 3236 22985 3238
rect 23009 3236 23065 3238
rect 23089 3236 23145 3238
rect 17376 2746 17432 2748
rect 17456 2746 17512 2748
rect 17536 2746 17592 2748
rect 17616 2746 17672 2748
rect 17376 2694 17422 2746
rect 17422 2694 17432 2746
rect 17456 2694 17486 2746
rect 17486 2694 17498 2746
rect 17498 2694 17512 2746
rect 17536 2694 17550 2746
rect 17550 2694 17562 2746
rect 17562 2694 17592 2746
rect 17616 2694 17626 2746
rect 17626 2694 17672 2746
rect 17376 2692 17432 2694
rect 17456 2692 17512 2694
rect 17536 2692 17592 2694
rect 17616 2692 17672 2694
rect 28323 6010 28379 6012
rect 28403 6010 28459 6012
rect 28483 6010 28539 6012
rect 28563 6010 28619 6012
rect 28323 5958 28369 6010
rect 28369 5958 28379 6010
rect 28403 5958 28433 6010
rect 28433 5958 28445 6010
rect 28445 5958 28459 6010
rect 28483 5958 28497 6010
rect 28497 5958 28509 6010
rect 28509 5958 28539 6010
rect 28563 5958 28573 6010
rect 28573 5958 28619 6010
rect 28323 5956 28379 5958
rect 28403 5956 28459 5958
rect 28483 5956 28539 5958
rect 28563 5956 28619 5958
rect 30194 6296 30250 6352
rect 28323 4922 28379 4924
rect 28403 4922 28459 4924
rect 28483 4922 28539 4924
rect 28563 4922 28619 4924
rect 28323 4870 28369 4922
rect 28369 4870 28379 4922
rect 28403 4870 28433 4922
rect 28433 4870 28445 4922
rect 28445 4870 28459 4922
rect 28483 4870 28497 4922
rect 28497 4870 28509 4922
rect 28509 4870 28539 4922
rect 28563 4870 28573 4922
rect 28573 4870 28619 4922
rect 28323 4868 28379 4870
rect 28403 4868 28459 4870
rect 28483 4868 28539 4870
rect 28563 4868 28619 4870
rect 28323 3834 28379 3836
rect 28403 3834 28459 3836
rect 28483 3834 28539 3836
rect 28563 3834 28619 3836
rect 28323 3782 28369 3834
rect 28369 3782 28379 3834
rect 28403 3782 28433 3834
rect 28433 3782 28445 3834
rect 28445 3782 28459 3834
rect 28483 3782 28497 3834
rect 28497 3782 28509 3834
rect 28509 3782 28539 3834
rect 28563 3782 28573 3834
rect 28573 3782 28619 3834
rect 28323 3780 28379 3782
rect 28403 3780 28459 3782
rect 28483 3780 28539 3782
rect 28563 3780 28619 3782
rect 28323 2746 28379 2748
rect 28403 2746 28459 2748
rect 28483 2746 28539 2748
rect 28563 2746 28619 2748
rect 28323 2694 28369 2746
rect 28369 2694 28379 2746
rect 28403 2694 28433 2746
rect 28433 2694 28445 2746
rect 28445 2694 28459 2746
rect 28483 2694 28497 2746
rect 28497 2694 28509 2746
rect 28509 2694 28539 2746
rect 28563 2694 28573 2746
rect 28573 2694 28619 2746
rect 28323 2692 28379 2694
rect 28403 2692 28459 2694
rect 28483 2692 28539 2694
rect 28563 2692 28619 2694
rect 22849 2202 22905 2204
rect 22929 2202 22985 2204
rect 23009 2202 23065 2204
rect 23089 2202 23145 2204
rect 22849 2150 22895 2202
rect 22895 2150 22905 2202
rect 22929 2150 22959 2202
rect 22959 2150 22971 2202
rect 22971 2150 22985 2202
rect 23009 2150 23023 2202
rect 23023 2150 23035 2202
rect 23035 2150 23065 2202
rect 23089 2150 23099 2202
rect 23099 2150 23145 2202
rect 22849 2148 22905 2150
rect 22929 2148 22985 2150
rect 23009 2148 23065 2150
rect 23089 2148 23145 2150
rect 33796 10906 33852 10908
rect 33876 10906 33932 10908
rect 33956 10906 34012 10908
rect 34036 10906 34092 10908
rect 33796 10854 33842 10906
rect 33842 10854 33852 10906
rect 33876 10854 33906 10906
rect 33906 10854 33918 10906
rect 33918 10854 33932 10906
rect 33956 10854 33970 10906
rect 33970 10854 33982 10906
rect 33982 10854 34012 10906
rect 34036 10854 34046 10906
rect 34046 10854 34092 10906
rect 33796 10852 33852 10854
rect 33876 10852 33932 10854
rect 33956 10852 34012 10854
rect 34036 10852 34092 10854
rect 33796 9818 33852 9820
rect 33876 9818 33932 9820
rect 33956 9818 34012 9820
rect 34036 9818 34092 9820
rect 33796 9766 33842 9818
rect 33842 9766 33852 9818
rect 33876 9766 33906 9818
rect 33906 9766 33918 9818
rect 33918 9766 33932 9818
rect 33956 9766 33970 9818
rect 33970 9766 33982 9818
rect 33982 9766 34012 9818
rect 34036 9766 34046 9818
rect 34046 9766 34092 9818
rect 33796 9764 33852 9766
rect 33876 9764 33932 9766
rect 33956 9764 34012 9766
rect 34036 9764 34092 9766
rect 33796 8730 33852 8732
rect 33876 8730 33932 8732
rect 33956 8730 34012 8732
rect 34036 8730 34092 8732
rect 33796 8678 33842 8730
rect 33842 8678 33852 8730
rect 33876 8678 33906 8730
rect 33906 8678 33918 8730
rect 33918 8678 33932 8730
rect 33956 8678 33970 8730
rect 33970 8678 33982 8730
rect 33982 8678 34012 8730
rect 34036 8678 34046 8730
rect 34046 8678 34092 8730
rect 33796 8676 33852 8678
rect 33876 8676 33932 8678
rect 33956 8676 34012 8678
rect 34036 8676 34092 8678
rect 33796 7642 33852 7644
rect 33876 7642 33932 7644
rect 33956 7642 34012 7644
rect 34036 7642 34092 7644
rect 33796 7590 33842 7642
rect 33842 7590 33852 7642
rect 33876 7590 33906 7642
rect 33906 7590 33918 7642
rect 33918 7590 33932 7642
rect 33956 7590 33970 7642
rect 33970 7590 33982 7642
rect 33982 7590 34012 7642
rect 34036 7590 34046 7642
rect 34046 7590 34092 7642
rect 33796 7588 33852 7590
rect 33876 7588 33932 7590
rect 33956 7588 34012 7590
rect 34036 7588 34092 7590
rect 32126 4528 32182 4584
rect 32954 6296 33010 6352
rect 33796 6554 33852 6556
rect 33876 6554 33932 6556
rect 33956 6554 34012 6556
rect 34036 6554 34092 6556
rect 33796 6502 33842 6554
rect 33842 6502 33852 6554
rect 33876 6502 33906 6554
rect 33906 6502 33918 6554
rect 33918 6502 33932 6554
rect 33956 6502 33970 6554
rect 33970 6502 33982 6554
rect 33982 6502 34012 6554
rect 34036 6502 34046 6554
rect 34046 6502 34092 6554
rect 33796 6500 33852 6502
rect 33876 6500 33932 6502
rect 33956 6500 34012 6502
rect 34036 6500 34092 6502
rect 34242 6316 34298 6352
rect 34242 6296 34244 6316
rect 34244 6296 34296 6316
rect 34296 6296 34298 6316
rect 33796 5466 33852 5468
rect 33876 5466 33932 5468
rect 33956 5466 34012 5468
rect 34036 5466 34092 5468
rect 33796 5414 33842 5466
rect 33842 5414 33852 5466
rect 33876 5414 33906 5466
rect 33906 5414 33918 5466
rect 33918 5414 33932 5466
rect 33956 5414 33970 5466
rect 33970 5414 33982 5466
rect 33982 5414 34012 5466
rect 34036 5414 34046 5466
rect 34046 5414 34092 5466
rect 33796 5412 33852 5414
rect 33876 5412 33932 5414
rect 33956 5412 34012 5414
rect 34036 5412 34092 5414
rect 39270 16890 39326 16892
rect 39350 16890 39406 16892
rect 39430 16890 39486 16892
rect 39510 16890 39566 16892
rect 39270 16838 39316 16890
rect 39316 16838 39326 16890
rect 39350 16838 39380 16890
rect 39380 16838 39392 16890
rect 39392 16838 39406 16890
rect 39430 16838 39444 16890
rect 39444 16838 39456 16890
rect 39456 16838 39486 16890
rect 39510 16838 39520 16890
rect 39520 16838 39566 16890
rect 39270 16836 39326 16838
rect 39350 16836 39406 16838
rect 39430 16836 39486 16838
rect 39510 16836 39566 16838
rect 45006 19080 45062 19136
rect 44270 17720 44326 17776
rect 44743 17434 44799 17436
rect 44823 17434 44879 17436
rect 44903 17434 44959 17436
rect 44983 17434 45039 17436
rect 44743 17382 44789 17434
rect 44789 17382 44799 17434
rect 44823 17382 44853 17434
rect 44853 17382 44865 17434
rect 44865 17382 44879 17434
rect 44903 17382 44917 17434
rect 44917 17382 44929 17434
rect 44929 17382 44959 17434
rect 44983 17382 44993 17434
rect 44993 17382 45039 17434
rect 44743 17380 44799 17382
rect 44823 17380 44879 17382
rect 44903 17380 44959 17382
rect 44983 17380 45039 17382
rect 44743 16346 44799 16348
rect 44823 16346 44879 16348
rect 44903 16346 44959 16348
rect 44983 16346 45039 16348
rect 44743 16294 44789 16346
rect 44789 16294 44799 16346
rect 44823 16294 44853 16346
rect 44853 16294 44865 16346
rect 44865 16294 44879 16346
rect 44903 16294 44917 16346
rect 44917 16294 44929 16346
rect 44929 16294 44959 16346
rect 44983 16294 44993 16346
rect 44993 16294 45039 16346
rect 44743 16292 44799 16294
rect 44823 16292 44879 16294
rect 44903 16292 44959 16294
rect 44983 16292 45039 16294
rect 39270 15802 39326 15804
rect 39350 15802 39406 15804
rect 39430 15802 39486 15804
rect 39510 15802 39566 15804
rect 39270 15750 39316 15802
rect 39316 15750 39326 15802
rect 39350 15750 39380 15802
rect 39380 15750 39392 15802
rect 39392 15750 39406 15802
rect 39430 15750 39444 15802
rect 39444 15750 39456 15802
rect 39456 15750 39486 15802
rect 39510 15750 39520 15802
rect 39520 15750 39566 15802
rect 39270 15748 39326 15750
rect 39350 15748 39406 15750
rect 39430 15748 39486 15750
rect 39510 15748 39566 15750
rect 44362 15680 44418 15736
rect 44743 15258 44799 15260
rect 44823 15258 44879 15260
rect 44903 15258 44959 15260
rect 44983 15258 45039 15260
rect 44743 15206 44789 15258
rect 44789 15206 44799 15258
rect 44823 15206 44853 15258
rect 44853 15206 44865 15258
rect 44865 15206 44879 15258
rect 44903 15206 44917 15258
rect 44917 15206 44929 15258
rect 44929 15206 44959 15258
rect 44983 15206 44993 15258
rect 44993 15206 45039 15258
rect 44743 15204 44799 15206
rect 44823 15204 44879 15206
rect 44903 15204 44959 15206
rect 44983 15204 45039 15206
rect 39270 14714 39326 14716
rect 39350 14714 39406 14716
rect 39430 14714 39486 14716
rect 39510 14714 39566 14716
rect 39270 14662 39316 14714
rect 39316 14662 39326 14714
rect 39350 14662 39380 14714
rect 39380 14662 39392 14714
rect 39392 14662 39406 14714
rect 39430 14662 39444 14714
rect 39444 14662 39456 14714
rect 39456 14662 39486 14714
rect 39510 14662 39520 14714
rect 39520 14662 39566 14714
rect 39270 14660 39326 14662
rect 39350 14660 39406 14662
rect 39430 14660 39486 14662
rect 39510 14660 39566 14662
rect 33874 4564 33876 4584
rect 33876 4564 33928 4584
rect 33928 4564 33930 4584
rect 33874 4528 33930 4564
rect 33796 4378 33852 4380
rect 33876 4378 33932 4380
rect 33956 4378 34012 4380
rect 34036 4378 34092 4380
rect 33796 4326 33842 4378
rect 33842 4326 33852 4378
rect 33876 4326 33906 4378
rect 33906 4326 33918 4378
rect 33918 4326 33932 4378
rect 33956 4326 33970 4378
rect 33970 4326 33982 4378
rect 33982 4326 34012 4378
rect 34036 4326 34046 4378
rect 34046 4326 34092 4378
rect 33796 4324 33852 4326
rect 33876 4324 33932 4326
rect 33956 4324 34012 4326
rect 34036 4324 34092 4326
rect 33796 3290 33852 3292
rect 33876 3290 33932 3292
rect 33956 3290 34012 3292
rect 34036 3290 34092 3292
rect 33796 3238 33842 3290
rect 33842 3238 33852 3290
rect 33876 3238 33906 3290
rect 33906 3238 33918 3290
rect 33918 3238 33932 3290
rect 33956 3238 33970 3290
rect 33970 3238 33982 3290
rect 33982 3238 34012 3290
rect 34036 3238 34046 3290
rect 34046 3238 34092 3290
rect 33796 3236 33852 3238
rect 33876 3236 33932 3238
rect 33956 3236 34012 3238
rect 34036 3236 34092 3238
rect 39270 13626 39326 13628
rect 39350 13626 39406 13628
rect 39430 13626 39486 13628
rect 39510 13626 39566 13628
rect 39270 13574 39316 13626
rect 39316 13574 39326 13626
rect 39350 13574 39380 13626
rect 39380 13574 39392 13626
rect 39392 13574 39406 13626
rect 39430 13574 39444 13626
rect 39444 13574 39456 13626
rect 39456 13574 39486 13626
rect 39510 13574 39520 13626
rect 39520 13574 39566 13626
rect 39270 13572 39326 13574
rect 39350 13572 39406 13574
rect 39430 13572 39486 13574
rect 39510 13572 39566 13574
rect 39394 13232 39450 13288
rect 39270 12538 39326 12540
rect 39350 12538 39406 12540
rect 39430 12538 39486 12540
rect 39510 12538 39566 12540
rect 39270 12486 39316 12538
rect 39316 12486 39326 12538
rect 39350 12486 39380 12538
rect 39380 12486 39392 12538
rect 39392 12486 39406 12538
rect 39430 12486 39444 12538
rect 39444 12486 39456 12538
rect 39456 12486 39486 12538
rect 39510 12486 39520 12538
rect 39520 12486 39566 12538
rect 39270 12484 39326 12486
rect 39350 12484 39406 12486
rect 39430 12484 39486 12486
rect 39510 12484 39566 12486
rect 39210 11736 39266 11792
rect 39270 11450 39326 11452
rect 39350 11450 39406 11452
rect 39430 11450 39486 11452
rect 39510 11450 39566 11452
rect 39270 11398 39316 11450
rect 39316 11398 39326 11450
rect 39350 11398 39380 11450
rect 39380 11398 39392 11450
rect 39392 11398 39406 11450
rect 39430 11398 39444 11450
rect 39444 11398 39456 11450
rect 39456 11398 39486 11450
rect 39510 11398 39520 11450
rect 39520 11398 39566 11450
rect 39270 11396 39326 11398
rect 39350 11396 39406 11398
rect 39430 11396 39486 11398
rect 39510 11396 39566 11398
rect 41878 12724 41880 12744
rect 41880 12724 41932 12744
rect 41932 12724 41934 12744
rect 42982 14456 43038 14512
rect 44270 14320 44326 14376
rect 44743 14170 44799 14172
rect 44823 14170 44879 14172
rect 44903 14170 44959 14172
rect 44983 14170 45039 14172
rect 44743 14118 44789 14170
rect 44789 14118 44799 14170
rect 44823 14118 44853 14170
rect 44853 14118 44865 14170
rect 44865 14118 44879 14170
rect 44903 14118 44917 14170
rect 44917 14118 44929 14170
rect 44929 14118 44959 14170
rect 44983 14118 44993 14170
rect 44993 14118 45039 14170
rect 44743 14116 44799 14118
rect 44823 14116 44879 14118
rect 44903 14116 44959 14118
rect 44983 14116 45039 14118
rect 44743 13082 44799 13084
rect 44823 13082 44879 13084
rect 44903 13082 44959 13084
rect 44983 13082 45039 13084
rect 44743 13030 44789 13082
rect 44789 13030 44799 13082
rect 44823 13030 44853 13082
rect 44853 13030 44865 13082
rect 44865 13030 44879 13082
rect 44903 13030 44917 13082
rect 44917 13030 44929 13082
rect 44929 13030 44959 13082
rect 44983 13030 44993 13082
rect 44993 13030 45039 13082
rect 44743 13028 44799 13030
rect 44823 13028 44879 13030
rect 44903 13028 44959 13030
rect 44983 13028 45039 13030
rect 41878 12688 41934 12724
rect 45006 12280 45062 12336
rect 44743 11994 44799 11996
rect 44823 11994 44879 11996
rect 44903 11994 44959 11996
rect 44983 11994 45039 11996
rect 44743 11942 44789 11994
rect 44789 11942 44799 11994
rect 44823 11942 44853 11994
rect 44853 11942 44865 11994
rect 44865 11942 44879 11994
rect 44903 11942 44917 11994
rect 44917 11942 44929 11994
rect 44929 11942 44959 11994
rect 44983 11942 44993 11994
rect 44993 11942 45039 11994
rect 44743 11940 44799 11942
rect 44823 11940 44879 11942
rect 44903 11940 44959 11942
rect 44983 11940 45039 11942
rect 39270 10362 39326 10364
rect 39350 10362 39406 10364
rect 39430 10362 39486 10364
rect 39510 10362 39566 10364
rect 39270 10310 39316 10362
rect 39316 10310 39326 10362
rect 39350 10310 39380 10362
rect 39380 10310 39392 10362
rect 39392 10310 39406 10362
rect 39430 10310 39444 10362
rect 39444 10310 39456 10362
rect 39456 10310 39486 10362
rect 39510 10310 39520 10362
rect 39520 10310 39566 10362
rect 39270 10308 39326 10310
rect 39350 10308 39406 10310
rect 39430 10308 39486 10310
rect 39510 10308 39566 10310
rect 45006 11092 45008 11112
rect 45008 11092 45060 11112
rect 45060 11092 45062 11112
rect 45006 11056 45062 11092
rect 44743 10906 44799 10908
rect 44823 10906 44879 10908
rect 44903 10906 44959 10908
rect 44983 10906 45039 10908
rect 44743 10854 44789 10906
rect 44789 10854 44799 10906
rect 44823 10854 44853 10906
rect 44853 10854 44865 10906
rect 44865 10854 44879 10906
rect 44903 10854 44917 10906
rect 44917 10854 44929 10906
rect 44929 10854 44959 10906
rect 44983 10854 44993 10906
rect 44993 10854 45039 10906
rect 44743 10852 44799 10854
rect 44823 10852 44879 10854
rect 44903 10852 44959 10854
rect 44983 10852 45039 10854
rect 39270 9274 39326 9276
rect 39350 9274 39406 9276
rect 39430 9274 39486 9276
rect 39510 9274 39566 9276
rect 39270 9222 39316 9274
rect 39316 9222 39326 9274
rect 39350 9222 39380 9274
rect 39380 9222 39392 9274
rect 39392 9222 39406 9274
rect 39430 9222 39444 9274
rect 39444 9222 39456 9274
rect 39456 9222 39486 9274
rect 39510 9222 39520 9274
rect 39520 9222 39566 9274
rect 39270 9220 39326 9222
rect 39350 9220 39406 9222
rect 39430 9220 39486 9222
rect 39510 9220 39566 9222
rect 39270 8186 39326 8188
rect 39350 8186 39406 8188
rect 39430 8186 39486 8188
rect 39510 8186 39566 8188
rect 39270 8134 39316 8186
rect 39316 8134 39326 8186
rect 39350 8134 39380 8186
rect 39380 8134 39392 8186
rect 39392 8134 39406 8186
rect 39430 8134 39444 8186
rect 39444 8134 39456 8186
rect 39456 8134 39486 8186
rect 39510 8134 39520 8186
rect 39520 8134 39566 8186
rect 39270 8132 39326 8134
rect 39350 8132 39406 8134
rect 39430 8132 39486 8134
rect 39510 8132 39566 8134
rect 39270 7098 39326 7100
rect 39350 7098 39406 7100
rect 39430 7098 39486 7100
rect 39510 7098 39566 7100
rect 39270 7046 39316 7098
rect 39316 7046 39326 7098
rect 39350 7046 39380 7098
rect 39380 7046 39392 7098
rect 39392 7046 39406 7098
rect 39430 7046 39444 7098
rect 39444 7046 39456 7098
rect 39456 7046 39486 7098
rect 39510 7046 39520 7098
rect 39520 7046 39566 7098
rect 39270 7044 39326 7046
rect 39350 7044 39406 7046
rect 39430 7044 39486 7046
rect 39510 7044 39566 7046
rect 39270 6010 39326 6012
rect 39350 6010 39406 6012
rect 39430 6010 39486 6012
rect 39510 6010 39566 6012
rect 39270 5958 39316 6010
rect 39316 5958 39326 6010
rect 39350 5958 39380 6010
rect 39380 5958 39392 6010
rect 39392 5958 39406 6010
rect 39430 5958 39444 6010
rect 39444 5958 39456 6010
rect 39456 5958 39486 6010
rect 39510 5958 39520 6010
rect 39520 5958 39566 6010
rect 39270 5956 39326 5958
rect 39350 5956 39406 5958
rect 39430 5956 39486 5958
rect 39510 5956 39566 5958
rect 39270 4922 39326 4924
rect 39350 4922 39406 4924
rect 39430 4922 39486 4924
rect 39510 4922 39566 4924
rect 39270 4870 39316 4922
rect 39316 4870 39326 4922
rect 39350 4870 39380 4922
rect 39380 4870 39392 4922
rect 39392 4870 39406 4922
rect 39430 4870 39444 4922
rect 39444 4870 39456 4922
rect 39456 4870 39486 4922
rect 39510 4870 39520 4922
rect 39520 4870 39566 4922
rect 39270 4868 39326 4870
rect 39350 4868 39406 4870
rect 39430 4868 39486 4870
rect 39510 4868 39566 4870
rect 39270 3834 39326 3836
rect 39350 3834 39406 3836
rect 39430 3834 39486 3836
rect 39510 3834 39566 3836
rect 39270 3782 39316 3834
rect 39316 3782 39326 3834
rect 39350 3782 39380 3834
rect 39380 3782 39392 3834
rect 39392 3782 39406 3834
rect 39430 3782 39444 3834
rect 39444 3782 39456 3834
rect 39456 3782 39486 3834
rect 39510 3782 39520 3834
rect 39520 3782 39566 3834
rect 39270 3780 39326 3782
rect 39350 3780 39406 3782
rect 39430 3780 39486 3782
rect 39510 3780 39566 3782
rect 39270 2746 39326 2748
rect 39350 2746 39406 2748
rect 39430 2746 39486 2748
rect 39510 2746 39566 2748
rect 39270 2694 39316 2746
rect 39316 2694 39326 2746
rect 39350 2694 39380 2746
rect 39380 2694 39392 2746
rect 39392 2694 39406 2746
rect 39430 2694 39444 2746
rect 39444 2694 39456 2746
rect 39456 2694 39486 2746
rect 39510 2694 39520 2746
rect 39520 2694 39566 2746
rect 39270 2692 39326 2694
rect 39350 2692 39406 2694
rect 39430 2692 39486 2694
rect 39510 2692 39566 2694
rect 44178 8880 44234 8936
rect 44362 8916 44364 8936
rect 44364 8916 44416 8936
rect 44416 8916 44418 8936
rect 44362 8880 44418 8916
rect 44362 7404 44418 7440
rect 44362 7384 44364 7404
rect 44364 7384 44416 7404
rect 44416 7384 44418 7404
rect 44270 4120 44326 4176
rect 44743 9818 44799 9820
rect 44823 9818 44879 9820
rect 44903 9818 44959 9820
rect 44983 9818 45039 9820
rect 44743 9766 44789 9818
rect 44789 9766 44799 9818
rect 44823 9766 44853 9818
rect 44853 9766 44865 9818
rect 44865 9766 44879 9818
rect 44903 9766 44917 9818
rect 44917 9766 44929 9818
rect 44929 9766 44959 9818
rect 44983 9766 44993 9818
rect 44993 9766 45039 9818
rect 44743 9764 44799 9766
rect 44823 9764 44879 9766
rect 44903 9764 44959 9766
rect 44983 9764 45039 9766
rect 44743 8730 44799 8732
rect 44823 8730 44879 8732
rect 44903 8730 44959 8732
rect 44983 8730 45039 8732
rect 44743 8678 44789 8730
rect 44789 8678 44799 8730
rect 44823 8678 44853 8730
rect 44853 8678 44865 8730
rect 44865 8678 44879 8730
rect 44903 8678 44917 8730
rect 44917 8678 44929 8730
rect 44929 8678 44959 8730
rect 44983 8678 44993 8730
rect 44993 8678 45039 8730
rect 44743 8676 44799 8678
rect 44823 8676 44879 8678
rect 44903 8676 44959 8678
rect 44983 8676 45039 8678
rect 44743 7642 44799 7644
rect 44823 7642 44879 7644
rect 44903 7642 44959 7644
rect 44983 7642 45039 7644
rect 44743 7590 44789 7642
rect 44789 7590 44799 7642
rect 44823 7590 44853 7642
rect 44853 7590 44865 7642
rect 44865 7590 44879 7642
rect 44903 7590 44917 7642
rect 44917 7590 44929 7642
rect 44929 7590 44959 7642
rect 44983 7590 44993 7642
rect 44993 7590 45039 7642
rect 44743 7588 44799 7590
rect 44823 7588 44879 7590
rect 44903 7588 44959 7590
rect 44983 7588 45039 7590
rect 44743 6554 44799 6556
rect 44823 6554 44879 6556
rect 44903 6554 44959 6556
rect 44983 6554 45039 6556
rect 44743 6502 44789 6554
rect 44789 6502 44799 6554
rect 44823 6502 44853 6554
rect 44853 6502 44865 6554
rect 44865 6502 44879 6554
rect 44903 6502 44917 6554
rect 44917 6502 44929 6554
rect 44929 6502 44959 6554
rect 44983 6502 44993 6554
rect 44993 6502 45039 6554
rect 44743 6500 44799 6502
rect 44823 6500 44879 6502
rect 44903 6500 44959 6502
rect 44983 6500 45039 6502
rect 45006 5616 45062 5672
rect 44743 5466 44799 5468
rect 44823 5466 44879 5468
rect 44903 5466 44959 5468
rect 44983 5466 45039 5468
rect 44743 5414 44789 5466
rect 44789 5414 44799 5466
rect 44823 5414 44853 5466
rect 44853 5414 44865 5466
rect 44865 5414 44879 5466
rect 44903 5414 44917 5466
rect 44917 5414 44929 5466
rect 44929 5414 44959 5466
rect 44983 5414 44993 5466
rect 44993 5414 45039 5466
rect 44743 5412 44799 5414
rect 44823 5412 44879 5414
rect 44903 5412 44959 5414
rect 44983 5412 45039 5414
rect 44743 4378 44799 4380
rect 44823 4378 44879 4380
rect 44903 4378 44959 4380
rect 44983 4378 45039 4380
rect 44743 4326 44789 4378
rect 44789 4326 44799 4378
rect 44823 4326 44853 4378
rect 44853 4326 44865 4378
rect 44865 4326 44879 4378
rect 44903 4326 44917 4378
rect 44917 4326 44929 4378
rect 44929 4326 44959 4378
rect 44983 4326 44993 4378
rect 44993 4326 45039 4378
rect 44743 4324 44799 4326
rect 44823 4324 44879 4326
rect 44903 4324 44959 4326
rect 44983 4324 45039 4326
rect 33796 2202 33852 2204
rect 33876 2202 33932 2204
rect 33956 2202 34012 2204
rect 34036 2202 34092 2204
rect 33796 2150 33842 2202
rect 33842 2150 33852 2202
rect 33876 2150 33906 2202
rect 33906 2150 33918 2202
rect 33918 2150 33932 2202
rect 33956 2150 33970 2202
rect 33970 2150 33982 2202
rect 33982 2150 34012 2202
rect 34036 2150 34046 2202
rect 34046 2150 34092 2202
rect 33796 2148 33852 2150
rect 33876 2148 33932 2150
rect 33956 2148 34012 2150
rect 34036 2148 34092 2150
rect 44270 1944 44326 2000
rect 44743 3290 44799 3292
rect 44823 3290 44879 3292
rect 44903 3290 44959 3292
rect 44983 3290 45039 3292
rect 44743 3238 44789 3290
rect 44789 3238 44799 3290
rect 44823 3238 44853 3290
rect 44853 3238 44865 3290
rect 44865 3238 44879 3290
rect 44903 3238 44917 3290
rect 44917 3238 44929 3290
rect 44929 3238 44959 3290
rect 44983 3238 44993 3290
rect 44993 3238 45039 3290
rect 44743 3236 44799 3238
rect 44823 3236 44879 3238
rect 44903 3236 44959 3238
rect 44983 3236 45039 3238
rect 44743 2202 44799 2204
rect 44823 2202 44879 2204
rect 44903 2202 44959 2204
rect 44983 2202 45039 2204
rect 44743 2150 44789 2202
rect 44789 2150 44799 2202
rect 44823 2150 44853 2202
rect 44853 2150 44865 2202
rect 44865 2150 44879 2202
rect 44903 2150 44917 2202
rect 44917 2150 44929 2202
rect 44929 2150 44959 2202
rect 44983 2150 44993 2202
rect 44993 2150 45039 2202
rect 44743 2148 44799 2150
rect 44823 2148 44879 2150
rect 44903 2148 44959 2150
rect 44983 2148 45039 2150
rect 44638 720 44694 776
<< metal3 >>
rect 45001 19138 45067 19141
rect 45200 19138 46000 19228
rect 45001 19136 46000 19138
rect 45001 19080 45006 19136
rect 45062 19080 46000 19136
rect 45001 19078 46000 19080
rect 45001 19075 45067 19078
rect 45200 18988 46000 19078
rect 0 18458 800 18548
rect 1025 18458 1091 18461
rect 0 18456 1091 18458
rect 0 18400 1030 18456
rect 1086 18400 1091 18456
rect 0 18398 1091 18400
rect 0 18308 800 18398
rect 1025 18395 1091 18398
rect 44265 17778 44331 17781
rect 45200 17778 46000 17868
rect 44265 17776 46000 17778
rect 44265 17720 44270 17776
rect 44326 17720 46000 17776
rect 44265 17718 46000 17720
rect 44265 17715 44331 17718
rect 45200 17628 46000 17718
rect 11892 17440 12208 17441
rect 11892 17376 11898 17440
rect 11962 17376 11978 17440
rect 12042 17376 12058 17440
rect 12122 17376 12138 17440
rect 12202 17376 12208 17440
rect 11892 17375 12208 17376
rect 22839 17440 23155 17441
rect 22839 17376 22845 17440
rect 22909 17376 22925 17440
rect 22989 17376 23005 17440
rect 23069 17376 23085 17440
rect 23149 17376 23155 17440
rect 22839 17375 23155 17376
rect 33786 17440 34102 17441
rect 33786 17376 33792 17440
rect 33856 17376 33872 17440
rect 33936 17376 33952 17440
rect 34016 17376 34032 17440
rect 34096 17376 34102 17440
rect 33786 17375 34102 17376
rect 44733 17440 45049 17441
rect 44733 17376 44739 17440
rect 44803 17376 44819 17440
rect 44883 17376 44899 17440
rect 44963 17376 44979 17440
rect 45043 17376 45049 17440
rect 44733 17375 45049 17376
rect 0 17098 800 17188
rect 933 17098 999 17101
rect 0 17096 999 17098
rect 0 17040 938 17096
rect 994 17040 999 17096
rect 0 17038 999 17040
rect 0 16948 800 17038
rect 933 17035 999 17038
rect 6419 16896 6735 16897
rect 6419 16832 6425 16896
rect 6489 16832 6505 16896
rect 6569 16832 6585 16896
rect 6649 16832 6665 16896
rect 6729 16832 6735 16896
rect 6419 16831 6735 16832
rect 17366 16896 17682 16897
rect 17366 16832 17372 16896
rect 17436 16832 17452 16896
rect 17516 16832 17532 16896
rect 17596 16832 17612 16896
rect 17676 16832 17682 16896
rect 17366 16831 17682 16832
rect 28313 16896 28629 16897
rect 28313 16832 28319 16896
rect 28383 16832 28399 16896
rect 28463 16832 28479 16896
rect 28543 16832 28559 16896
rect 28623 16832 28629 16896
rect 28313 16831 28629 16832
rect 39260 16896 39576 16897
rect 39260 16832 39266 16896
rect 39330 16832 39346 16896
rect 39410 16832 39426 16896
rect 39490 16832 39506 16896
rect 39570 16832 39576 16896
rect 39260 16831 39576 16832
rect 11892 16352 12208 16353
rect 11892 16288 11898 16352
rect 11962 16288 11978 16352
rect 12042 16288 12058 16352
rect 12122 16288 12138 16352
rect 12202 16288 12208 16352
rect 11892 16287 12208 16288
rect 22839 16352 23155 16353
rect 22839 16288 22845 16352
rect 22909 16288 22925 16352
rect 22989 16288 23005 16352
rect 23069 16288 23085 16352
rect 23149 16288 23155 16352
rect 22839 16287 23155 16288
rect 33786 16352 34102 16353
rect 33786 16288 33792 16352
rect 33856 16288 33872 16352
rect 33936 16288 33952 16352
rect 34016 16288 34032 16352
rect 34096 16288 34102 16352
rect 33786 16287 34102 16288
rect 44733 16352 45049 16353
rect 44733 16288 44739 16352
rect 44803 16288 44819 16352
rect 44883 16288 44899 16352
rect 44963 16288 44979 16352
rect 45043 16288 45049 16352
rect 44733 16287 45049 16288
rect 6419 15808 6735 15809
rect 6419 15744 6425 15808
rect 6489 15744 6505 15808
rect 6569 15744 6585 15808
rect 6649 15744 6665 15808
rect 6729 15744 6735 15808
rect 6419 15743 6735 15744
rect 17366 15808 17682 15809
rect 17366 15744 17372 15808
rect 17436 15744 17452 15808
rect 17516 15744 17532 15808
rect 17596 15744 17612 15808
rect 17676 15744 17682 15808
rect 17366 15743 17682 15744
rect 28313 15808 28629 15809
rect 28313 15744 28319 15808
rect 28383 15744 28399 15808
rect 28463 15744 28479 15808
rect 28543 15744 28559 15808
rect 28623 15744 28629 15808
rect 28313 15743 28629 15744
rect 39260 15808 39576 15809
rect 39260 15744 39266 15808
rect 39330 15744 39346 15808
rect 39410 15744 39426 15808
rect 39490 15744 39506 15808
rect 39570 15744 39576 15808
rect 39260 15743 39576 15744
rect 44357 15738 44423 15741
rect 45200 15738 46000 15828
rect 44357 15736 46000 15738
rect 44357 15680 44362 15736
rect 44418 15680 46000 15736
rect 44357 15678 46000 15680
rect 44357 15675 44423 15678
rect 45200 15588 46000 15678
rect 11892 15264 12208 15265
rect 11892 15200 11898 15264
rect 11962 15200 11978 15264
rect 12042 15200 12058 15264
rect 12122 15200 12138 15264
rect 12202 15200 12208 15264
rect 11892 15199 12208 15200
rect 22839 15264 23155 15265
rect 22839 15200 22845 15264
rect 22909 15200 22925 15264
rect 22989 15200 23005 15264
rect 23069 15200 23085 15264
rect 23149 15200 23155 15264
rect 22839 15199 23155 15200
rect 33786 15264 34102 15265
rect 33786 15200 33792 15264
rect 33856 15200 33872 15264
rect 33936 15200 33952 15264
rect 34016 15200 34032 15264
rect 34096 15200 34102 15264
rect 33786 15199 34102 15200
rect 44733 15264 45049 15265
rect 44733 15200 44739 15264
rect 44803 15200 44819 15264
rect 44883 15200 44899 15264
rect 44963 15200 44979 15264
rect 45043 15200 45049 15264
rect 44733 15199 45049 15200
rect 0 15058 800 15148
rect 933 15058 999 15061
rect 0 15056 999 15058
rect 0 15000 938 15056
rect 994 15000 999 15056
rect 0 14998 999 15000
rect 0 14908 800 14998
rect 933 14995 999 14998
rect 32581 14922 32647 14925
rect 33961 14922 34027 14925
rect 32581 14920 34027 14922
rect 32581 14864 32586 14920
rect 32642 14864 33966 14920
rect 34022 14864 34027 14920
rect 32581 14862 34027 14864
rect 32581 14859 32647 14862
rect 33961 14859 34027 14862
rect 6419 14720 6735 14721
rect 6419 14656 6425 14720
rect 6489 14656 6505 14720
rect 6569 14656 6585 14720
rect 6649 14656 6665 14720
rect 6729 14656 6735 14720
rect 6419 14655 6735 14656
rect 17366 14720 17682 14721
rect 17366 14656 17372 14720
rect 17436 14656 17452 14720
rect 17516 14656 17532 14720
rect 17596 14656 17612 14720
rect 17676 14656 17682 14720
rect 17366 14655 17682 14656
rect 28313 14720 28629 14721
rect 28313 14656 28319 14720
rect 28383 14656 28399 14720
rect 28463 14656 28479 14720
rect 28543 14656 28559 14720
rect 28623 14656 28629 14720
rect 28313 14655 28629 14656
rect 39260 14720 39576 14721
rect 39260 14656 39266 14720
rect 39330 14656 39346 14720
rect 39410 14656 39426 14720
rect 39490 14656 39506 14720
rect 39570 14656 39576 14720
rect 39260 14655 39576 14656
rect 16297 14514 16363 14517
rect 42977 14514 43043 14517
rect 16297 14512 43043 14514
rect 16297 14456 16302 14512
rect 16358 14456 42982 14512
rect 43038 14456 43043 14512
rect 16297 14454 43043 14456
rect 16297 14451 16363 14454
rect 42977 14451 43043 14454
rect 44265 14378 44331 14381
rect 45200 14378 46000 14468
rect 44265 14376 46000 14378
rect 44265 14320 44270 14376
rect 44326 14320 46000 14376
rect 44265 14318 46000 14320
rect 44265 14315 44331 14318
rect 45200 14228 46000 14318
rect 11892 14176 12208 14177
rect 11892 14112 11898 14176
rect 11962 14112 11978 14176
rect 12042 14112 12058 14176
rect 12122 14112 12138 14176
rect 12202 14112 12208 14176
rect 11892 14111 12208 14112
rect 22839 14176 23155 14177
rect 22839 14112 22845 14176
rect 22909 14112 22925 14176
rect 22989 14112 23005 14176
rect 23069 14112 23085 14176
rect 23149 14112 23155 14176
rect 22839 14111 23155 14112
rect 33786 14176 34102 14177
rect 33786 14112 33792 14176
rect 33856 14112 33872 14176
rect 33936 14112 33952 14176
rect 34016 14112 34032 14176
rect 34096 14112 34102 14176
rect 33786 14111 34102 14112
rect 44733 14176 45049 14177
rect 44733 14112 44739 14176
rect 44803 14112 44819 14176
rect 44883 14112 44899 14176
rect 44963 14112 44979 14176
rect 45043 14112 45049 14176
rect 44733 14111 45049 14112
rect 0 13698 800 13788
rect 933 13698 999 13701
rect 0 13696 999 13698
rect 0 13640 938 13696
rect 994 13640 999 13696
rect 0 13638 999 13640
rect 0 13548 800 13638
rect 933 13635 999 13638
rect 6419 13632 6735 13633
rect 6419 13568 6425 13632
rect 6489 13568 6505 13632
rect 6569 13568 6585 13632
rect 6649 13568 6665 13632
rect 6729 13568 6735 13632
rect 6419 13567 6735 13568
rect 17366 13632 17682 13633
rect 17366 13568 17372 13632
rect 17436 13568 17452 13632
rect 17516 13568 17532 13632
rect 17596 13568 17612 13632
rect 17676 13568 17682 13632
rect 17366 13567 17682 13568
rect 28313 13632 28629 13633
rect 28313 13568 28319 13632
rect 28383 13568 28399 13632
rect 28463 13568 28479 13632
rect 28543 13568 28559 13632
rect 28623 13568 28629 13632
rect 28313 13567 28629 13568
rect 39260 13632 39576 13633
rect 39260 13568 39266 13632
rect 39330 13568 39346 13632
rect 39410 13568 39426 13632
rect 39490 13568 39506 13632
rect 39570 13568 39576 13632
rect 39260 13567 39576 13568
rect 32489 13290 32555 13293
rect 39389 13290 39455 13293
rect 32489 13288 39455 13290
rect 32489 13232 32494 13288
rect 32550 13232 39394 13288
rect 39450 13232 39455 13288
rect 32489 13230 39455 13232
rect 32489 13227 32555 13230
rect 39389 13227 39455 13230
rect 11892 13088 12208 13089
rect 11892 13024 11898 13088
rect 11962 13024 11978 13088
rect 12042 13024 12058 13088
rect 12122 13024 12138 13088
rect 12202 13024 12208 13088
rect 11892 13023 12208 13024
rect 22839 13088 23155 13089
rect 22839 13024 22845 13088
rect 22909 13024 22925 13088
rect 22989 13024 23005 13088
rect 23069 13024 23085 13088
rect 23149 13024 23155 13088
rect 22839 13023 23155 13024
rect 33786 13088 34102 13089
rect 33786 13024 33792 13088
rect 33856 13024 33872 13088
rect 33936 13024 33952 13088
rect 34016 13024 34032 13088
rect 34096 13024 34102 13088
rect 33786 13023 34102 13024
rect 44733 13088 45049 13089
rect 44733 13024 44739 13088
rect 44803 13024 44819 13088
rect 44883 13024 44899 13088
rect 44963 13024 44979 13088
rect 45043 13024 45049 13088
rect 44733 13023 45049 13024
rect 3141 12882 3207 12885
rect 24761 12882 24827 12885
rect 3141 12880 24827 12882
rect 3141 12824 3146 12880
rect 3202 12824 24766 12880
rect 24822 12824 24827 12880
rect 3141 12822 24827 12824
rect 3141 12819 3207 12822
rect 24761 12819 24827 12822
rect 31569 12882 31635 12885
rect 33501 12882 33567 12885
rect 31569 12880 33567 12882
rect 31569 12824 31574 12880
rect 31630 12824 33506 12880
rect 33562 12824 33567 12880
rect 31569 12822 33567 12824
rect 31569 12819 31635 12822
rect 33501 12819 33567 12822
rect 32581 12746 32647 12749
rect 41873 12746 41939 12749
rect 32581 12744 41939 12746
rect 32581 12688 32586 12744
rect 32642 12688 41878 12744
rect 41934 12688 41939 12744
rect 32581 12686 41939 12688
rect 32581 12683 32647 12686
rect 41873 12683 41939 12686
rect 6419 12544 6735 12545
rect 6419 12480 6425 12544
rect 6489 12480 6505 12544
rect 6569 12480 6585 12544
rect 6649 12480 6665 12544
rect 6729 12480 6735 12544
rect 6419 12479 6735 12480
rect 17366 12544 17682 12545
rect 17366 12480 17372 12544
rect 17436 12480 17452 12544
rect 17516 12480 17532 12544
rect 17596 12480 17612 12544
rect 17676 12480 17682 12544
rect 17366 12479 17682 12480
rect 28313 12544 28629 12545
rect 28313 12480 28319 12544
rect 28383 12480 28399 12544
rect 28463 12480 28479 12544
rect 28543 12480 28559 12544
rect 28623 12480 28629 12544
rect 28313 12479 28629 12480
rect 39260 12544 39576 12545
rect 39260 12480 39266 12544
rect 39330 12480 39346 12544
rect 39410 12480 39426 12544
rect 39490 12480 39506 12544
rect 39570 12480 39576 12544
rect 39260 12479 39576 12480
rect 45001 12338 45067 12341
rect 45200 12338 46000 12428
rect 45001 12336 46000 12338
rect 45001 12280 45006 12336
rect 45062 12280 46000 12336
rect 45001 12278 46000 12280
rect 45001 12275 45067 12278
rect 45200 12188 46000 12278
rect 11892 12000 12208 12001
rect 11892 11936 11898 12000
rect 11962 11936 11978 12000
rect 12042 11936 12058 12000
rect 12122 11936 12138 12000
rect 12202 11936 12208 12000
rect 11892 11935 12208 11936
rect 22839 12000 23155 12001
rect 22839 11936 22845 12000
rect 22909 11936 22925 12000
rect 22989 11936 23005 12000
rect 23069 11936 23085 12000
rect 23149 11936 23155 12000
rect 22839 11935 23155 11936
rect 33786 12000 34102 12001
rect 33786 11936 33792 12000
rect 33856 11936 33872 12000
rect 33936 11936 33952 12000
rect 34016 11936 34032 12000
rect 34096 11936 34102 12000
rect 33786 11935 34102 11936
rect 44733 12000 45049 12001
rect 44733 11936 44739 12000
rect 44803 11936 44819 12000
rect 44883 11936 44899 12000
rect 44963 11936 44979 12000
rect 45043 11936 45049 12000
rect 44733 11935 45049 11936
rect 4061 11930 4127 11933
rect 4061 11928 4170 11930
rect 4061 11872 4066 11928
rect 4122 11872 4170 11928
rect 4061 11867 4170 11872
rect 4110 11794 4170 11867
rect 39205 11794 39271 11797
rect 4110 11792 39271 11794
rect 0 11658 800 11748
rect 4110 11736 39210 11792
rect 39266 11736 39271 11792
rect 4110 11734 39271 11736
rect 39205 11731 39271 11734
rect 4061 11658 4127 11661
rect 0 11656 4127 11658
rect 0 11600 4066 11656
rect 4122 11600 4127 11656
rect 0 11598 4127 11600
rect 0 11508 800 11598
rect 4061 11595 4127 11598
rect 6419 11456 6735 11457
rect 6419 11392 6425 11456
rect 6489 11392 6505 11456
rect 6569 11392 6585 11456
rect 6649 11392 6665 11456
rect 6729 11392 6735 11456
rect 6419 11391 6735 11392
rect 17366 11456 17682 11457
rect 17366 11392 17372 11456
rect 17436 11392 17452 11456
rect 17516 11392 17532 11456
rect 17596 11392 17612 11456
rect 17676 11392 17682 11456
rect 17366 11391 17682 11392
rect 28313 11456 28629 11457
rect 28313 11392 28319 11456
rect 28383 11392 28399 11456
rect 28463 11392 28479 11456
rect 28543 11392 28559 11456
rect 28623 11392 28629 11456
rect 28313 11391 28629 11392
rect 39260 11456 39576 11457
rect 39260 11392 39266 11456
rect 39330 11392 39346 11456
rect 39410 11392 39426 11456
rect 39490 11392 39506 11456
rect 39570 11392 39576 11456
rect 39260 11391 39576 11392
rect 45001 11114 45067 11117
rect 45001 11112 45202 11114
rect 45001 11056 45006 11112
rect 45062 11068 45202 11112
rect 45062 11056 46000 11068
rect 45001 11054 46000 11056
rect 45001 11051 45067 11054
rect 45142 10918 46000 11054
rect 11892 10912 12208 10913
rect 11892 10848 11898 10912
rect 11962 10848 11978 10912
rect 12042 10848 12058 10912
rect 12122 10848 12138 10912
rect 12202 10848 12208 10912
rect 11892 10847 12208 10848
rect 22839 10912 23155 10913
rect 22839 10848 22845 10912
rect 22909 10848 22925 10912
rect 22989 10848 23005 10912
rect 23069 10848 23085 10912
rect 23149 10848 23155 10912
rect 22839 10847 23155 10848
rect 33786 10912 34102 10913
rect 33786 10848 33792 10912
rect 33856 10848 33872 10912
rect 33936 10848 33952 10912
rect 34016 10848 34032 10912
rect 34096 10848 34102 10912
rect 33786 10847 34102 10848
rect 44733 10912 45049 10913
rect 44733 10848 44739 10912
rect 44803 10848 44819 10912
rect 44883 10848 44899 10912
rect 44963 10848 44979 10912
rect 45043 10848 45049 10912
rect 44733 10847 45049 10848
rect 45200 10828 46000 10918
rect 0 10298 800 10388
rect 6419 10368 6735 10369
rect 6419 10304 6425 10368
rect 6489 10304 6505 10368
rect 6569 10304 6585 10368
rect 6649 10304 6665 10368
rect 6729 10304 6735 10368
rect 6419 10303 6735 10304
rect 17366 10368 17682 10369
rect 17366 10304 17372 10368
rect 17436 10304 17452 10368
rect 17516 10304 17532 10368
rect 17596 10304 17612 10368
rect 17676 10304 17682 10368
rect 17366 10303 17682 10304
rect 28313 10368 28629 10369
rect 28313 10304 28319 10368
rect 28383 10304 28399 10368
rect 28463 10304 28479 10368
rect 28543 10304 28559 10368
rect 28623 10304 28629 10368
rect 28313 10303 28629 10304
rect 39260 10368 39576 10369
rect 39260 10304 39266 10368
rect 39330 10304 39346 10368
rect 39410 10304 39426 10368
rect 39490 10304 39506 10368
rect 39570 10304 39576 10368
rect 39260 10303 39576 10304
rect 933 10298 999 10301
rect 0 10296 999 10298
rect 0 10240 938 10296
rect 994 10240 999 10296
rect 0 10238 999 10240
rect 0 10148 800 10238
rect 933 10235 999 10238
rect 12801 10026 12867 10029
rect 29821 10026 29887 10029
rect 12801 10024 29887 10026
rect 12801 9968 12806 10024
rect 12862 9968 29826 10024
rect 29882 9968 29887 10024
rect 12801 9966 29887 9968
rect 12801 9963 12867 9966
rect 29821 9963 29887 9966
rect 11892 9824 12208 9825
rect 11892 9760 11898 9824
rect 11962 9760 11978 9824
rect 12042 9760 12058 9824
rect 12122 9760 12138 9824
rect 12202 9760 12208 9824
rect 11892 9759 12208 9760
rect 22839 9824 23155 9825
rect 22839 9760 22845 9824
rect 22909 9760 22925 9824
rect 22989 9760 23005 9824
rect 23069 9760 23085 9824
rect 23149 9760 23155 9824
rect 22839 9759 23155 9760
rect 33786 9824 34102 9825
rect 33786 9760 33792 9824
rect 33856 9760 33872 9824
rect 33936 9760 33952 9824
rect 34016 9760 34032 9824
rect 34096 9760 34102 9824
rect 33786 9759 34102 9760
rect 44733 9824 45049 9825
rect 44733 9760 44739 9824
rect 44803 9760 44819 9824
rect 44883 9760 44899 9824
rect 44963 9760 44979 9824
rect 45043 9760 45049 9824
rect 44733 9759 45049 9760
rect 6419 9280 6735 9281
rect 6419 9216 6425 9280
rect 6489 9216 6505 9280
rect 6569 9216 6585 9280
rect 6649 9216 6665 9280
rect 6729 9216 6735 9280
rect 6419 9215 6735 9216
rect 17366 9280 17682 9281
rect 17366 9216 17372 9280
rect 17436 9216 17452 9280
rect 17516 9216 17532 9280
rect 17596 9216 17612 9280
rect 17676 9216 17682 9280
rect 17366 9215 17682 9216
rect 28313 9280 28629 9281
rect 28313 9216 28319 9280
rect 28383 9216 28399 9280
rect 28463 9216 28479 9280
rect 28543 9216 28559 9280
rect 28623 9216 28629 9280
rect 28313 9215 28629 9216
rect 39260 9280 39576 9281
rect 39260 9216 39266 9280
rect 39330 9216 39346 9280
rect 39410 9216 39426 9280
rect 39490 9216 39506 9280
rect 39570 9216 39576 9280
rect 39260 9215 39576 9216
rect 27705 8938 27771 8941
rect 44173 8938 44239 8941
rect 27705 8936 44239 8938
rect 27705 8880 27710 8936
rect 27766 8880 44178 8936
rect 44234 8880 44239 8936
rect 27705 8878 44239 8880
rect 27705 8875 27771 8878
rect 44173 8875 44239 8878
rect 44357 8938 44423 8941
rect 45200 8938 46000 9028
rect 44357 8936 46000 8938
rect 44357 8880 44362 8936
rect 44418 8880 46000 8936
rect 44357 8878 46000 8880
rect 44357 8875 44423 8878
rect 45200 8788 46000 8878
rect 11892 8736 12208 8737
rect 11892 8672 11898 8736
rect 11962 8672 11978 8736
rect 12042 8672 12058 8736
rect 12122 8672 12138 8736
rect 12202 8672 12208 8736
rect 11892 8671 12208 8672
rect 22839 8736 23155 8737
rect 22839 8672 22845 8736
rect 22909 8672 22925 8736
rect 22989 8672 23005 8736
rect 23069 8672 23085 8736
rect 23149 8672 23155 8736
rect 22839 8671 23155 8672
rect 33786 8736 34102 8737
rect 33786 8672 33792 8736
rect 33856 8672 33872 8736
rect 33936 8672 33952 8736
rect 34016 8672 34032 8736
rect 34096 8672 34102 8736
rect 33786 8671 34102 8672
rect 44733 8736 45049 8737
rect 44733 8672 44739 8736
rect 44803 8672 44819 8736
rect 44883 8672 44899 8736
rect 44963 8672 44979 8736
rect 45043 8672 45049 8736
rect 44733 8671 45049 8672
rect 0 8258 800 8348
rect 933 8258 999 8261
rect 0 8256 999 8258
rect 0 8200 938 8256
rect 994 8200 999 8256
rect 0 8198 999 8200
rect 0 8108 800 8198
rect 933 8195 999 8198
rect 6419 8192 6735 8193
rect 6419 8128 6425 8192
rect 6489 8128 6505 8192
rect 6569 8128 6585 8192
rect 6649 8128 6665 8192
rect 6729 8128 6735 8192
rect 6419 8127 6735 8128
rect 17366 8192 17682 8193
rect 17366 8128 17372 8192
rect 17436 8128 17452 8192
rect 17516 8128 17532 8192
rect 17596 8128 17612 8192
rect 17676 8128 17682 8192
rect 17366 8127 17682 8128
rect 28313 8192 28629 8193
rect 28313 8128 28319 8192
rect 28383 8128 28399 8192
rect 28463 8128 28479 8192
rect 28543 8128 28559 8192
rect 28623 8128 28629 8192
rect 28313 8127 28629 8128
rect 39260 8192 39576 8193
rect 39260 8128 39266 8192
rect 39330 8128 39346 8192
rect 39410 8128 39426 8192
rect 39490 8128 39506 8192
rect 39570 8128 39576 8192
rect 39260 8127 39576 8128
rect 14825 7986 14891 7989
rect 27613 7986 27679 7989
rect 14825 7984 27679 7986
rect 14825 7928 14830 7984
rect 14886 7928 27618 7984
rect 27674 7928 27679 7984
rect 14825 7926 27679 7928
rect 14825 7923 14891 7926
rect 27613 7923 27679 7926
rect 11892 7648 12208 7649
rect 11892 7584 11898 7648
rect 11962 7584 11978 7648
rect 12042 7584 12058 7648
rect 12122 7584 12138 7648
rect 12202 7584 12208 7648
rect 11892 7583 12208 7584
rect 22839 7648 23155 7649
rect 22839 7584 22845 7648
rect 22909 7584 22925 7648
rect 22989 7584 23005 7648
rect 23069 7584 23085 7648
rect 23149 7584 23155 7648
rect 22839 7583 23155 7584
rect 33786 7648 34102 7649
rect 33786 7584 33792 7648
rect 33856 7584 33872 7648
rect 33936 7584 33952 7648
rect 34016 7584 34032 7648
rect 34096 7584 34102 7648
rect 33786 7583 34102 7584
rect 44733 7648 45049 7649
rect 44733 7584 44739 7648
rect 44803 7584 44819 7648
rect 44883 7584 44899 7648
rect 44963 7584 44979 7648
rect 45043 7584 45049 7648
rect 44733 7583 45049 7584
rect 45200 7578 46000 7668
rect 44357 7442 44423 7445
rect 45142 7442 46000 7578
rect 44357 7440 46000 7442
rect 44357 7384 44362 7440
rect 44418 7428 46000 7440
rect 44418 7384 45202 7428
rect 44357 7382 45202 7384
rect 44357 7379 44423 7382
rect 6419 7104 6735 7105
rect 6419 7040 6425 7104
rect 6489 7040 6505 7104
rect 6569 7040 6585 7104
rect 6649 7040 6665 7104
rect 6729 7040 6735 7104
rect 6419 7039 6735 7040
rect 17366 7104 17682 7105
rect 17366 7040 17372 7104
rect 17436 7040 17452 7104
rect 17516 7040 17532 7104
rect 17596 7040 17612 7104
rect 17676 7040 17682 7104
rect 17366 7039 17682 7040
rect 28313 7104 28629 7105
rect 28313 7040 28319 7104
rect 28383 7040 28399 7104
rect 28463 7040 28479 7104
rect 28543 7040 28559 7104
rect 28623 7040 28629 7104
rect 28313 7039 28629 7040
rect 39260 7104 39576 7105
rect 39260 7040 39266 7104
rect 39330 7040 39346 7104
rect 39410 7040 39426 7104
rect 39490 7040 39506 7104
rect 39570 7040 39576 7104
rect 39260 7039 39576 7040
rect 0 6898 800 6988
rect 933 6898 999 6901
rect 0 6896 999 6898
rect 0 6840 938 6896
rect 994 6840 999 6896
rect 0 6838 999 6840
rect 0 6748 800 6838
rect 933 6835 999 6838
rect 11892 6560 12208 6561
rect 11892 6496 11898 6560
rect 11962 6496 11978 6560
rect 12042 6496 12058 6560
rect 12122 6496 12138 6560
rect 12202 6496 12208 6560
rect 11892 6495 12208 6496
rect 22839 6560 23155 6561
rect 22839 6496 22845 6560
rect 22909 6496 22925 6560
rect 22989 6496 23005 6560
rect 23069 6496 23085 6560
rect 23149 6496 23155 6560
rect 22839 6495 23155 6496
rect 33786 6560 34102 6561
rect 33786 6496 33792 6560
rect 33856 6496 33872 6560
rect 33936 6496 33952 6560
rect 34016 6496 34032 6560
rect 34096 6496 34102 6560
rect 33786 6495 34102 6496
rect 44733 6560 45049 6561
rect 44733 6496 44739 6560
rect 44803 6496 44819 6560
rect 44883 6496 44899 6560
rect 44963 6496 44979 6560
rect 45043 6496 45049 6560
rect 44733 6495 45049 6496
rect 12065 6354 12131 6357
rect 17769 6354 17835 6357
rect 30189 6354 30255 6357
rect 12065 6352 30255 6354
rect 12065 6296 12070 6352
rect 12126 6296 17774 6352
rect 17830 6296 30194 6352
rect 30250 6296 30255 6352
rect 12065 6294 30255 6296
rect 12065 6291 12131 6294
rect 17769 6291 17835 6294
rect 30189 6291 30255 6294
rect 32949 6354 33015 6357
rect 34237 6354 34303 6357
rect 32949 6352 34303 6354
rect 32949 6296 32954 6352
rect 33010 6296 34242 6352
rect 34298 6296 34303 6352
rect 32949 6294 34303 6296
rect 32949 6291 33015 6294
rect 34237 6291 34303 6294
rect 13629 6218 13695 6221
rect 25313 6218 25379 6221
rect 13629 6216 25379 6218
rect 13629 6160 13634 6216
rect 13690 6160 25318 6216
rect 25374 6160 25379 6216
rect 13629 6158 25379 6160
rect 13629 6155 13695 6158
rect 25313 6155 25379 6158
rect 6419 6016 6735 6017
rect 6419 5952 6425 6016
rect 6489 5952 6505 6016
rect 6569 5952 6585 6016
rect 6649 5952 6665 6016
rect 6729 5952 6735 6016
rect 6419 5951 6735 5952
rect 17366 6016 17682 6017
rect 17366 5952 17372 6016
rect 17436 5952 17452 6016
rect 17516 5952 17532 6016
rect 17596 5952 17612 6016
rect 17676 5952 17682 6016
rect 17366 5951 17682 5952
rect 28313 6016 28629 6017
rect 28313 5952 28319 6016
rect 28383 5952 28399 6016
rect 28463 5952 28479 6016
rect 28543 5952 28559 6016
rect 28623 5952 28629 6016
rect 28313 5951 28629 5952
rect 39260 6016 39576 6017
rect 39260 5952 39266 6016
rect 39330 5952 39346 6016
rect 39410 5952 39426 6016
rect 39490 5952 39506 6016
rect 39570 5952 39576 6016
rect 39260 5951 39576 5952
rect 45001 5674 45067 5677
rect 45001 5672 45202 5674
rect 45001 5616 45006 5672
rect 45062 5628 45202 5672
rect 45062 5616 46000 5628
rect 45001 5614 46000 5616
rect 45001 5611 45067 5614
rect 45142 5478 46000 5614
rect 11892 5472 12208 5473
rect 11892 5408 11898 5472
rect 11962 5408 11978 5472
rect 12042 5408 12058 5472
rect 12122 5408 12138 5472
rect 12202 5408 12208 5472
rect 11892 5407 12208 5408
rect 22839 5472 23155 5473
rect 22839 5408 22845 5472
rect 22909 5408 22925 5472
rect 22989 5408 23005 5472
rect 23069 5408 23085 5472
rect 23149 5408 23155 5472
rect 22839 5407 23155 5408
rect 33786 5472 34102 5473
rect 33786 5408 33792 5472
rect 33856 5408 33872 5472
rect 33936 5408 33952 5472
rect 34016 5408 34032 5472
rect 34096 5408 34102 5472
rect 33786 5407 34102 5408
rect 44733 5472 45049 5473
rect 44733 5408 44739 5472
rect 44803 5408 44819 5472
rect 44883 5408 44899 5472
rect 44963 5408 44979 5472
rect 45043 5408 45049 5472
rect 44733 5407 45049 5408
rect 45200 5388 46000 5478
rect 0 4858 800 4948
rect 6419 4928 6735 4929
rect 6419 4864 6425 4928
rect 6489 4864 6505 4928
rect 6569 4864 6585 4928
rect 6649 4864 6665 4928
rect 6729 4864 6735 4928
rect 6419 4863 6735 4864
rect 17366 4928 17682 4929
rect 17366 4864 17372 4928
rect 17436 4864 17452 4928
rect 17516 4864 17532 4928
rect 17596 4864 17612 4928
rect 17676 4864 17682 4928
rect 17366 4863 17682 4864
rect 28313 4928 28629 4929
rect 28313 4864 28319 4928
rect 28383 4864 28399 4928
rect 28463 4864 28479 4928
rect 28543 4864 28559 4928
rect 28623 4864 28629 4928
rect 28313 4863 28629 4864
rect 39260 4928 39576 4929
rect 39260 4864 39266 4928
rect 39330 4864 39346 4928
rect 39410 4864 39426 4928
rect 39490 4864 39506 4928
rect 39570 4864 39576 4928
rect 39260 4863 39576 4864
rect 933 4858 999 4861
rect 0 4856 999 4858
rect 0 4800 938 4856
rect 994 4800 999 4856
rect 0 4798 999 4800
rect 0 4708 800 4798
rect 933 4795 999 4798
rect 32121 4586 32187 4589
rect 33869 4586 33935 4589
rect 32121 4584 33935 4586
rect 32121 4528 32126 4584
rect 32182 4528 33874 4584
rect 33930 4528 33935 4584
rect 32121 4526 33935 4528
rect 32121 4523 32187 4526
rect 33869 4523 33935 4526
rect 11892 4384 12208 4385
rect 11892 4320 11898 4384
rect 11962 4320 11978 4384
rect 12042 4320 12058 4384
rect 12122 4320 12138 4384
rect 12202 4320 12208 4384
rect 11892 4319 12208 4320
rect 22839 4384 23155 4385
rect 22839 4320 22845 4384
rect 22909 4320 22925 4384
rect 22989 4320 23005 4384
rect 23069 4320 23085 4384
rect 23149 4320 23155 4384
rect 22839 4319 23155 4320
rect 33786 4384 34102 4385
rect 33786 4320 33792 4384
rect 33856 4320 33872 4384
rect 33936 4320 33952 4384
rect 34016 4320 34032 4384
rect 34096 4320 34102 4384
rect 33786 4319 34102 4320
rect 44733 4384 45049 4385
rect 44733 4320 44739 4384
rect 44803 4320 44819 4384
rect 44883 4320 44899 4384
rect 44963 4320 44979 4384
rect 45043 4320 45049 4384
rect 44733 4319 45049 4320
rect 44265 4178 44331 4181
rect 45200 4178 46000 4268
rect 44265 4176 46000 4178
rect 44265 4120 44270 4176
rect 44326 4120 46000 4176
rect 44265 4118 46000 4120
rect 44265 4115 44331 4118
rect 45200 4028 46000 4118
rect 6419 3840 6735 3841
rect 6419 3776 6425 3840
rect 6489 3776 6505 3840
rect 6569 3776 6585 3840
rect 6649 3776 6665 3840
rect 6729 3776 6735 3840
rect 6419 3775 6735 3776
rect 17366 3840 17682 3841
rect 17366 3776 17372 3840
rect 17436 3776 17452 3840
rect 17516 3776 17532 3840
rect 17596 3776 17612 3840
rect 17676 3776 17682 3840
rect 17366 3775 17682 3776
rect 28313 3840 28629 3841
rect 28313 3776 28319 3840
rect 28383 3776 28399 3840
rect 28463 3776 28479 3840
rect 28543 3776 28559 3840
rect 28623 3776 28629 3840
rect 28313 3775 28629 3776
rect 39260 3840 39576 3841
rect 39260 3776 39266 3840
rect 39330 3776 39346 3840
rect 39410 3776 39426 3840
rect 39490 3776 39506 3840
rect 39570 3776 39576 3840
rect 39260 3775 39576 3776
rect 0 3498 800 3588
rect 933 3498 999 3501
rect 0 3496 999 3498
rect 0 3440 938 3496
rect 994 3440 999 3496
rect 0 3438 999 3440
rect 0 3348 800 3438
rect 933 3435 999 3438
rect 11892 3296 12208 3297
rect 11892 3232 11898 3296
rect 11962 3232 11978 3296
rect 12042 3232 12058 3296
rect 12122 3232 12138 3296
rect 12202 3232 12208 3296
rect 11892 3231 12208 3232
rect 22839 3296 23155 3297
rect 22839 3232 22845 3296
rect 22909 3232 22925 3296
rect 22989 3232 23005 3296
rect 23069 3232 23085 3296
rect 23149 3232 23155 3296
rect 22839 3231 23155 3232
rect 33786 3296 34102 3297
rect 33786 3232 33792 3296
rect 33856 3232 33872 3296
rect 33936 3232 33952 3296
rect 34016 3232 34032 3296
rect 34096 3232 34102 3296
rect 33786 3231 34102 3232
rect 44733 3296 45049 3297
rect 44733 3232 44739 3296
rect 44803 3232 44819 3296
rect 44883 3232 44899 3296
rect 44963 3232 44979 3296
rect 45043 3232 45049 3296
rect 44733 3231 45049 3232
rect 6419 2752 6735 2753
rect 6419 2688 6425 2752
rect 6489 2688 6505 2752
rect 6569 2688 6585 2752
rect 6649 2688 6665 2752
rect 6729 2688 6735 2752
rect 6419 2687 6735 2688
rect 17366 2752 17682 2753
rect 17366 2688 17372 2752
rect 17436 2688 17452 2752
rect 17516 2688 17532 2752
rect 17596 2688 17612 2752
rect 17676 2688 17682 2752
rect 17366 2687 17682 2688
rect 28313 2752 28629 2753
rect 28313 2688 28319 2752
rect 28383 2688 28399 2752
rect 28463 2688 28479 2752
rect 28543 2688 28559 2752
rect 28623 2688 28629 2752
rect 28313 2687 28629 2688
rect 39260 2752 39576 2753
rect 39260 2688 39266 2752
rect 39330 2688 39346 2752
rect 39410 2688 39426 2752
rect 39490 2688 39506 2752
rect 39570 2688 39576 2752
rect 39260 2687 39576 2688
rect 11892 2208 12208 2209
rect 11892 2144 11898 2208
rect 11962 2144 11978 2208
rect 12042 2144 12058 2208
rect 12122 2144 12138 2208
rect 12202 2144 12208 2208
rect 11892 2143 12208 2144
rect 22839 2208 23155 2209
rect 22839 2144 22845 2208
rect 22909 2144 22925 2208
rect 22989 2144 23005 2208
rect 23069 2144 23085 2208
rect 23149 2144 23155 2208
rect 22839 2143 23155 2144
rect 33786 2208 34102 2209
rect 33786 2144 33792 2208
rect 33856 2144 33872 2208
rect 33936 2144 33952 2208
rect 34016 2144 34032 2208
rect 34096 2144 34102 2208
rect 33786 2143 34102 2144
rect 44733 2208 45049 2209
rect 44733 2144 44739 2208
rect 44803 2144 44819 2208
rect 44883 2144 44899 2208
rect 44963 2144 44979 2208
rect 45043 2144 45049 2208
rect 44733 2143 45049 2144
rect 45200 2138 46000 2228
rect 44265 2002 44331 2005
rect 45142 2002 46000 2138
rect 44265 2000 46000 2002
rect 44265 1944 44270 2000
rect 44326 1988 46000 2000
rect 44326 1944 45202 1988
rect 44265 1942 45202 1944
rect 44265 1939 44331 1942
rect 0 1458 800 1548
rect 933 1458 999 1461
rect 0 1456 999 1458
rect 0 1400 938 1456
rect 994 1400 999 1456
rect 0 1398 999 1400
rect 0 1308 800 1398
rect 933 1395 999 1398
rect 44633 778 44699 781
rect 45200 778 46000 868
rect 44633 776 46000 778
rect 44633 720 44638 776
rect 44694 720 46000 776
rect 44633 718 46000 720
rect 44633 715 44699 718
rect 45200 628 46000 718
<< via3 >>
rect 11898 17436 11962 17440
rect 11898 17380 11902 17436
rect 11902 17380 11958 17436
rect 11958 17380 11962 17436
rect 11898 17376 11962 17380
rect 11978 17436 12042 17440
rect 11978 17380 11982 17436
rect 11982 17380 12038 17436
rect 12038 17380 12042 17436
rect 11978 17376 12042 17380
rect 12058 17436 12122 17440
rect 12058 17380 12062 17436
rect 12062 17380 12118 17436
rect 12118 17380 12122 17436
rect 12058 17376 12122 17380
rect 12138 17436 12202 17440
rect 12138 17380 12142 17436
rect 12142 17380 12198 17436
rect 12198 17380 12202 17436
rect 12138 17376 12202 17380
rect 22845 17436 22909 17440
rect 22845 17380 22849 17436
rect 22849 17380 22905 17436
rect 22905 17380 22909 17436
rect 22845 17376 22909 17380
rect 22925 17436 22989 17440
rect 22925 17380 22929 17436
rect 22929 17380 22985 17436
rect 22985 17380 22989 17436
rect 22925 17376 22989 17380
rect 23005 17436 23069 17440
rect 23005 17380 23009 17436
rect 23009 17380 23065 17436
rect 23065 17380 23069 17436
rect 23005 17376 23069 17380
rect 23085 17436 23149 17440
rect 23085 17380 23089 17436
rect 23089 17380 23145 17436
rect 23145 17380 23149 17436
rect 23085 17376 23149 17380
rect 33792 17436 33856 17440
rect 33792 17380 33796 17436
rect 33796 17380 33852 17436
rect 33852 17380 33856 17436
rect 33792 17376 33856 17380
rect 33872 17436 33936 17440
rect 33872 17380 33876 17436
rect 33876 17380 33932 17436
rect 33932 17380 33936 17436
rect 33872 17376 33936 17380
rect 33952 17436 34016 17440
rect 33952 17380 33956 17436
rect 33956 17380 34012 17436
rect 34012 17380 34016 17436
rect 33952 17376 34016 17380
rect 34032 17436 34096 17440
rect 34032 17380 34036 17436
rect 34036 17380 34092 17436
rect 34092 17380 34096 17436
rect 34032 17376 34096 17380
rect 44739 17436 44803 17440
rect 44739 17380 44743 17436
rect 44743 17380 44799 17436
rect 44799 17380 44803 17436
rect 44739 17376 44803 17380
rect 44819 17436 44883 17440
rect 44819 17380 44823 17436
rect 44823 17380 44879 17436
rect 44879 17380 44883 17436
rect 44819 17376 44883 17380
rect 44899 17436 44963 17440
rect 44899 17380 44903 17436
rect 44903 17380 44959 17436
rect 44959 17380 44963 17436
rect 44899 17376 44963 17380
rect 44979 17436 45043 17440
rect 44979 17380 44983 17436
rect 44983 17380 45039 17436
rect 45039 17380 45043 17436
rect 44979 17376 45043 17380
rect 6425 16892 6489 16896
rect 6425 16836 6429 16892
rect 6429 16836 6485 16892
rect 6485 16836 6489 16892
rect 6425 16832 6489 16836
rect 6505 16892 6569 16896
rect 6505 16836 6509 16892
rect 6509 16836 6565 16892
rect 6565 16836 6569 16892
rect 6505 16832 6569 16836
rect 6585 16892 6649 16896
rect 6585 16836 6589 16892
rect 6589 16836 6645 16892
rect 6645 16836 6649 16892
rect 6585 16832 6649 16836
rect 6665 16892 6729 16896
rect 6665 16836 6669 16892
rect 6669 16836 6725 16892
rect 6725 16836 6729 16892
rect 6665 16832 6729 16836
rect 17372 16892 17436 16896
rect 17372 16836 17376 16892
rect 17376 16836 17432 16892
rect 17432 16836 17436 16892
rect 17372 16832 17436 16836
rect 17452 16892 17516 16896
rect 17452 16836 17456 16892
rect 17456 16836 17512 16892
rect 17512 16836 17516 16892
rect 17452 16832 17516 16836
rect 17532 16892 17596 16896
rect 17532 16836 17536 16892
rect 17536 16836 17592 16892
rect 17592 16836 17596 16892
rect 17532 16832 17596 16836
rect 17612 16892 17676 16896
rect 17612 16836 17616 16892
rect 17616 16836 17672 16892
rect 17672 16836 17676 16892
rect 17612 16832 17676 16836
rect 28319 16892 28383 16896
rect 28319 16836 28323 16892
rect 28323 16836 28379 16892
rect 28379 16836 28383 16892
rect 28319 16832 28383 16836
rect 28399 16892 28463 16896
rect 28399 16836 28403 16892
rect 28403 16836 28459 16892
rect 28459 16836 28463 16892
rect 28399 16832 28463 16836
rect 28479 16892 28543 16896
rect 28479 16836 28483 16892
rect 28483 16836 28539 16892
rect 28539 16836 28543 16892
rect 28479 16832 28543 16836
rect 28559 16892 28623 16896
rect 28559 16836 28563 16892
rect 28563 16836 28619 16892
rect 28619 16836 28623 16892
rect 28559 16832 28623 16836
rect 39266 16892 39330 16896
rect 39266 16836 39270 16892
rect 39270 16836 39326 16892
rect 39326 16836 39330 16892
rect 39266 16832 39330 16836
rect 39346 16892 39410 16896
rect 39346 16836 39350 16892
rect 39350 16836 39406 16892
rect 39406 16836 39410 16892
rect 39346 16832 39410 16836
rect 39426 16892 39490 16896
rect 39426 16836 39430 16892
rect 39430 16836 39486 16892
rect 39486 16836 39490 16892
rect 39426 16832 39490 16836
rect 39506 16892 39570 16896
rect 39506 16836 39510 16892
rect 39510 16836 39566 16892
rect 39566 16836 39570 16892
rect 39506 16832 39570 16836
rect 11898 16348 11962 16352
rect 11898 16292 11902 16348
rect 11902 16292 11958 16348
rect 11958 16292 11962 16348
rect 11898 16288 11962 16292
rect 11978 16348 12042 16352
rect 11978 16292 11982 16348
rect 11982 16292 12038 16348
rect 12038 16292 12042 16348
rect 11978 16288 12042 16292
rect 12058 16348 12122 16352
rect 12058 16292 12062 16348
rect 12062 16292 12118 16348
rect 12118 16292 12122 16348
rect 12058 16288 12122 16292
rect 12138 16348 12202 16352
rect 12138 16292 12142 16348
rect 12142 16292 12198 16348
rect 12198 16292 12202 16348
rect 12138 16288 12202 16292
rect 22845 16348 22909 16352
rect 22845 16292 22849 16348
rect 22849 16292 22905 16348
rect 22905 16292 22909 16348
rect 22845 16288 22909 16292
rect 22925 16348 22989 16352
rect 22925 16292 22929 16348
rect 22929 16292 22985 16348
rect 22985 16292 22989 16348
rect 22925 16288 22989 16292
rect 23005 16348 23069 16352
rect 23005 16292 23009 16348
rect 23009 16292 23065 16348
rect 23065 16292 23069 16348
rect 23005 16288 23069 16292
rect 23085 16348 23149 16352
rect 23085 16292 23089 16348
rect 23089 16292 23145 16348
rect 23145 16292 23149 16348
rect 23085 16288 23149 16292
rect 33792 16348 33856 16352
rect 33792 16292 33796 16348
rect 33796 16292 33852 16348
rect 33852 16292 33856 16348
rect 33792 16288 33856 16292
rect 33872 16348 33936 16352
rect 33872 16292 33876 16348
rect 33876 16292 33932 16348
rect 33932 16292 33936 16348
rect 33872 16288 33936 16292
rect 33952 16348 34016 16352
rect 33952 16292 33956 16348
rect 33956 16292 34012 16348
rect 34012 16292 34016 16348
rect 33952 16288 34016 16292
rect 34032 16348 34096 16352
rect 34032 16292 34036 16348
rect 34036 16292 34092 16348
rect 34092 16292 34096 16348
rect 34032 16288 34096 16292
rect 44739 16348 44803 16352
rect 44739 16292 44743 16348
rect 44743 16292 44799 16348
rect 44799 16292 44803 16348
rect 44739 16288 44803 16292
rect 44819 16348 44883 16352
rect 44819 16292 44823 16348
rect 44823 16292 44879 16348
rect 44879 16292 44883 16348
rect 44819 16288 44883 16292
rect 44899 16348 44963 16352
rect 44899 16292 44903 16348
rect 44903 16292 44959 16348
rect 44959 16292 44963 16348
rect 44899 16288 44963 16292
rect 44979 16348 45043 16352
rect 44979 16292 44983 16348
rect 44983 16292 45039 16348
rect 45039 16292 45043 16348
rect 44979 16288 45043 16292
rect 6425 15804 6489 15808
rect 6425 15748 6429 15804
rect 6429 15748 6485 15804
rect 6485 15748 6489 15804
rect 6425 15744 6489 15748
rect 6505 15804 6569 15808
rect 6505 15748 6509 15804
rect 6509 15748 6565 15804
rect 6565 15748 6569 15804
rect 6505 15744 6569 15748
rect 6585 15804 6649 15808
rect 6585 15748 6589 15804
rect 6589 15748 6645 15804
rect 6645 15748 6649 15804
rect 6585 15744 6649 15748
rect 6665 15804 6729 15808
rect 6665 15748 6669 15804
rect 6669 15748 6725 15804
rect 6725 15748 6729 15804
rect 6665 15744 6729 15748
rect 17372 15804 17436 15808
rect 17372 15748 17376 15804
rect 17376 15748 17432 15804
rect 17432 15748 17436 15804
rect 17372 15744 17436 15748
rect 17452 15804 17516 15808
rect 17452 15748 17456 15804
rect 17456 15748 17512 15804
rect 17512 15748 17516 15804
rect 17452 15744 17516 15748
rect 17532 15804 17596 15808
rect 17532 15748 17536 15804
rect 17536 15748 17592 15804
rect 17592 15748 17596 15804
rect 17532 15744 17596 15748
rect 17612 15804 17676 15808
rect 17612 15748 17616 15804
rect 17616 15748 17672 15804
rect 17672 15748 17676 15804
rect 17612 15744 17676 15748
rect 28319 15804 28383 15808
rect 28319 15748 28323 15804
rect 28323 15748 28379 15804
rect 28379 15748 28383 15804
rect 28319 15744 28383 15748
rect 28399 15804 28463 15808
rect 28399 15748 28403 15804
rect 28403 15748 28459 15804
rect 28459 15748 28463 15804
rect 28399 15744 28463 15748
rect 28479 15804 28543 15808
rect 28479 15748 28483 15804
rect 28483 15748 28539 15804
rect 28539 15748 28543 15804
rect 28479 15744 28543 15748
rect 28559 15804 28623 15808
rect 28559 15748 28563 15804
rect 28563 15748 28619 15804
rect 28619 15748 28623 15804
rect 28559 15744 28623 15748
rect 39266 15804 39330 15808
rect 39266 15748 39270 15804
rect 39270 15748 39326 15804
rect 39326 15748 39330 15804
rect 39266 15744 39330 15748
rect 39346 15804 39410 15808
rect 39346 15748 39350 15804
rect 39350 15748 39406 15804
rect 39406 15748 39410 15804
rect 39346 15744 39410 15748
rect 39426 15804 39490 15808
rect 39426 15748 39430 15804
rect 39430 15748 39486 15804
rect 39486 15748 39490 15804
rect 39426 15744 39490 15748
rect 39506 15804 39570 15808
rect 39506 15748 39510 15804
rect 39510 15748 39566 15804
rect 39566 15748 39570 15804
rect 39506 15744 39570 15748
rect 11898 15260 11962 15264
rect 11898 15204 11902 15260
rect 11902 15204 11958 15260
rect 11958 15204 11962 15260
rect 11898 15200 11962 15204
rect 11978 15260 12042 15264
rect 11978 15204 11982 15260
rect 11982 15204 12038 15260
rect 12038 15204 12042 15260
rect 11978 15200 12042 15204
rect 12058 15260 12122 15264
rect 12058 15204 12062 15260
rect 12062 15204 12118 15260
rect 12118 15204 12122 15260
rect 12058 15200 12122 15204
rect 12138 15260 12202 15264
rect 12138 15204 12142 15260
rect 12142 15204 12198 15260
rect 12198 15204 12202 15260
rect 12138 15200 12202 15204
rect 22845 15260 22909 15264
rect 22845 15204 22849 15260
rect 22849 15204 22905 15260
rect 22905 15204 22909 15260
rect 22845 15200 22909 15204
rect 22925 15260 22989 15264
rect 22925 15204 22929 15260
rect 22929 15204 22985 15260
rect 22985 15204 22989 15260
rect 22925 15200 22989 15204
rect 23005 15260 23069 15264
rect 23005 15204 23009 15260
rect 23009 15204 23065 15260
rect 23065 15204 23069 15260
rect 23005 15200 23069 15204
rect 23085 15260 23149 15264
rect 23085 15204 23089 15260
rect 23089 15204 23145 15260
rect 23145 15204 23149 15260
rect 23085 15200 23149 15204
rect 33792 15260 33856 15264
rect 33792 15204 33796 15260
rect 33796 15204 33852 15260
rect 33852 15204 33856 15260
rect 33792 15200 33856 15204
rect 33872 15260 33936 15264
rect 33872 15204 33876 15260
rect 33876 15204 33932 15260
rect 33932 15204 33936 15260
rect 33872 15200 33936 15204
rect 33952 15260 34016 15264
rect 33952 15204 33956 15260
rect 33956 15204 34012 15260
rect 34012 15204 34016 15260
rect 33952 15200 34016 15204
rect 34032 15260 34096 15264
rect 34032 15204 34036 15260
rect 34036 15204 34092 15260
rect 34092 15204 34096 15260
rect 34032 15200 34096 15204
rect 44739 15260 44803 15264
rect 44739 15204 44743 15260
rect 44743 15204 44799 15260
rect 44799 15204 44803 15260
rect 44739 15200 44803 15204
rect 44819 15260 44883 15264
rect 44819 15204 44823 15260
rect 44823 15204 44879 15260
rect 44879 15204 44883 15260
rect 44819 15200 44883 15204
rect 44899 15260 44963 15264
rect 44899 15204 44903 15260
rect 44903 15204 44959 15260
rect 44959 15204 44963 15260
rect 44899 15200 44963 15204
rect 44979 15260 45043 15264
rect 44979 15204 44983 15260
rect 44983 15204 45039 15260
rect 45039 15204 45043 15260
rect 44979 15200 45043 15204
rect 6425 14716 6489 14720
rect 6425 14660 6429 14716
rect 6429 14660 6485 14716
rect 6485 14660 6489 14716
rect 6425 14656 6489 14660
rect 6505 14716 6569 14720
rect 6505 14660 6509 14716
rect 6509 14660 6565 14716
rect 6565 14660 6569 14716
rect 6505 14656 6569 14660
rect 6585 14716 6649 14720
rect 6585 14660 6589 14716
rect 6589 14660 6645 14716
rect 6645 14660 6649 14716
rect 6585 14656 6649 14660
rect 6665 14716 6729 14720
rect 6665 14660 6669 14716
rect 6669 14660 6725 14716
rect 6725 14660 6729 14716
rect 6665 14656 6729 14660
rect 17372 14716 17436 14720
rect 17372 14660 17376 14716
rect 17376 14660 17432 14716
rect 17432 14660 17436 14716
rect 17372 14656 17436 14660
rect 17452 14716 17516 14720
rect 17452 14660 17456 14716
rect 17456 14660 17512 14716
rect 17512 14660 17516 14716
rect 17452 14656 17516 14660
rect 17532 14716 17596 14720
rect 17532 14660 17536 14716
rect 17536 14660 17592 14716
rect 17592 14660 17596 14716
rect 17532 14656 17596 14660
rect 17612 14716 17676 14720
rect 17612 14660 17616 14716
rect 17616 14660 17672 14716
rect 17672 14660 17676 14716
rect 17612 14656 17676 14660
rect 28319 14716 28383 14720
rect 28319 14660 28323 14716
rect 28323 14660 28379 14716
rect 28379 14660 28383 14716
rect 28319 14656 28383 14660
rect 28399 14716 28463 14720
rect 28399 14660 28403 14716
rect 28403 14660 28459 14716
rect 28459 14660 28463 14716
rect 28399 14656 28463 14660
rect 28479 14716 28543 14720
rect 28479 14660 28483 14716
rect 28483 14660 28539 14716
rect 28539 14660 28543 14716
rect 28479 14656 28543 14660
rect 28559 14716 28623 14720
rect 28559 14660 28563 14716
rect 28563 14660 28619 14716
rect 28619 14660 28623 14716
rect 28559 14656 28623 14660
rect 39266 14716 39330 14720
rect 39266 14660 39270 14716
rect 39270 14660 39326 14716
rect 39326 14660 39330 14716
rect 39266 14656 39330 14660
rect 39346 14716 39410 14720
rect 39346 14660 39350 14716
rect 39350 14660 39406 14716
rect 39406 14660 39410 14716
rect 39346 14656 39410 14660
rect 39426 14716 39490 14720
rect 39426 14660 39430 14716
rect 39430 14660 39486 14716
rect 39486 14660 39490 14716
rect 39426 14656 39490 14660
rect 39506 14716 39570 14720
rect 39506 14660 39510 14716
rect 39510 14660 39566 14716
rect 39566 14660 39570 14716
rect 39506 14656 39570 14660
rect 11898 14172 11962 14176
rect 11898 14116 11902 14172
rect 11902 14116 11958 14172
rect 11958 14116 11962 14172
rect 11898 14112 11962 14116
rect 11978 14172 12042 14176
rect 11978 14116 11982 14172
rect 11982 14116 12038 14172
rect 12038 14116 12042 14172
rect 11978 14112 12042 14116
rect 12058 14172 12122 14176
rect 12058 14116 12062 14172
rect 12062 14116 12118 14172
rect 12118 14116 12122 14172
rect 12058 14112 12122 14116
rect 12138 14172 12202 14176
rect 12138 14116 12142 14172
rect 12142 14116 12198 14172
rect 12198 14116 12202 14172
rect 12138 14112 12202 14116
rect 22845 14172 22909 14176
rect 22845 14116 22849 14172
rect 22849 14116 22905 14172
rect 22905 14116 22909 14172
rect 22845 14112 22909 14116
rect 22925 14172 22989 14176
rect 22925 14116 22929 14172
rect 22929 14116 22985 14172
rect 22985 14116 22989 14172
rect 22925 14112 22989 14116
rect 23005 14172 23069 14176
rect 23005 14116 23009 14172
rect 23009 14116 23065 14172
rect 23065 14116 23069 14172
rect 23005 14112 23069 14116
rect 23085 14172 23149 14176
rect 23085 14116 23089 14172
rect 23089 14116 23145 14172
rect 23145 14116 23149 14172
rect 23085 14112 23149 14116
rect 33792 14172 33856 14176
rect 33792 14116 33796 14172
rect 33796 14116 33852 14172
rect 33852 14116 33856 14172
rect 33792 14112 33856 14116
rect 33872 14172 33936 14176
rect 33872 14116 33876 14172
rect 33876 14116 33932 14172
rect 33932 14116 33936 14172
rect 33872 14112 33936 14116
rect 33952 14172 34016 14176
rect 33952 14116 33956 14172
rect 33956 14116 34012 14172
rect 34012 14116 34016 14172
rect 33952 14112 34016 14116
rect 34032 14172 34096 14176
rect 34032 14116 34036 14172
rect 34036 14116 34092 14172
rect 34092 14116 34096 14172
rect 34032 14112 34096 14116
rect 44739 14172 44803 14176
rect 44739 14116 44743 14172
rect 44743 14116 44799 14172
rect 44799 14116 44803 14172
rect 44739 14112 44803 14116
rect 44819 14172 44883 14176
rect 44819 14116 44823 14172
rect 44823 14116 44879 14172
rect 44879 14116 44883 14172
rect 44819 14112 44883 14116
rect 44899 14172 44963 14176
rect 44899 14116 44903 14172
rect 44903 14116 44959 14172
rect 44959 14116 44963 14172
rect 44899 14112 44963 14116
rect 44979 14172 45043 14176
rect 44979 14116 44983 14172
rect 44983 14116 45039 14172
rect 45039 14116 45043 14172
rect 44979 14112 45043 14116
rect 6425 13628 6489 13632
rect 6425 13572 6429 13628
rect 6429 13572 6485 13628
rect 6485 13572 6489 13628
rect 6425 13568 6489 13572
rect 6505 13628 6569 13632
rect 6505 13572 6509 13628
rect 6509 13572 6565 13628
rect 6565 13572 6569 13628
rect 6505 13568 6569 13572
rect 6585 13628 6649 13632
rect 6585 13572 6589 13628
rect 6589 13572 6645 13628
rect 6645 13572 6649 13628
rect 6585 13568 6649 13572
rect 6665 13628 6729 13632
rect 6665 13572 6669 13628
rect 6669 13572 6725 13628
rect 6725 13572 6729 13628
rect 6665 13568 6729 13572
rect 17372 13628 17436 13632
rect 17372 13572 17376 13628
rect 17376 13572 17432 13628
rect 17432 13572 17436 13628
rect 17372 13568 17436 13572
rect 17452 13628 17516 13632
rect 17452 13572 17456 13628
rect 17456 13572 17512 13628
rect 17512 13572 17516 13628
rect 17452 13568 17516 13572
rect 17532 13628 17596 13632
rect 17532 13572 17536 13628
rect 17536 13572 17592 13628
rect 17592 13572 17596 13628
rect 17532 13568 17596 13572
rect 17612 13628 17676 13632
rect 17612 13572 17616 13628
rect 17616 13572 17672 13628
rect 17672 13572 17676 13628
rect 17612 13568 17676 13572
rect 28319 13628 28383 13632
rect 28319 13572 28323 13628
rect 28323 13572 28379 13628
rect 28379 13572 28383 13628
rect 28319 13568 28383 13572
rect 28399 13628 28463 13632
rect 28399 13572 28403 13628
rect 28403 13572 28459 13628
rect 28459 13572 28463 13628
rect 28399 13568 28463 13572
rect 28479 13628 28543 13632
rect 28479 13572 28483 13628
rect 28483 13572 28539 13628
rect 28539 13572 28543 13628
rect 28479 13568 28543 13572
rect 28559 13628 28623 13632
rect 28559 13572 28563 13628
rect 28563 13572 28619 13628
rect 28619 13572 28623 13628
rect 28559 13568 28623 13572
rect 39266 13628 39330 13632
rect 39266 13572 39270 13628
rect 39270 13572 39326 13628
rect 39326 13572 39330 13628
rect 39266 13568 39330 13572
rect 39346 13628 39410 13632
rect 39346 13572 39350 13628
rect 39350 13572 39406 13628
rect 39406 13572 39410 13628
rect 39346 13568 39410 13572
rect 39426 13628 39490 13632
rect 39426 13572 39430 13628
rect 39430 13572 39486 13628
rect 39486 13572 39490 13628
rect 39426 13568 39490 13572
rect 39506 13628 39570 13632
rect 39506 13572 39510 13628
rect 39510 13572 39566 13628
rect 39566 13572 39570 13628
rect 39506 13568 39570 13572
rect 11898 13084 11962 13088
rect 11898 13028 11902 13084
rect 11902 13028 11958 13084
rect 11958 13028 11962 13084
rect 11898 13024 11962 13028
rect 11978 13084 12042 13088
rect 11978 13028 11982 13084
rect 11982 13028 12038 13084
rect 12038 13028 12042 13084
rect 11978 13024 12042 13028
rect 12058 13084 12122 13088
rect 12058 13028 12062 13084
rect 12062 13028 12118 13084
rect 12118 13028 12122 13084
rect 12058 13024 12122 13028
rect 12138 13084 12202 13088
rect 12138 13028 12142 13084
rect 12142 13028 12198 13084
rect 12198 13028 12202 13084
rect 12138 13024 12202 13028
rect 22845 13084 22909 13088
rect 22845 13028 22849 13084
rect 22849 13028 22905 13084
rect 22905 13028 22909 13084
rect 22845 13024 22909 13028
rect 22925 13084 22989 13088
rect 22925 13028 22929 13084
rect 22929 13028 22985 13084
rect 22985 13028 22989 13084
rect 22925 13024 22989 13028
rect 23005 13084 23069 13088
rect 23005 13028 23009 13084
rect 23009 13028 23065 13084
rect 23065 13028 23069 13084
rect 23005 13024 23069 13028
rect 23085 13084 23149 13088
rect 23085 13028 23089 13084
rect 23089 13028 23145 13084
rect 23145 13028 23149 13084
rect 23085 13024 23149 13028
rect 33792 13084 33856 13088
rect 33792 13028 33796 13084
rect 33796 13028 33852 13084
rect 33852 13028 33856 13084
rect 33792 13024 33856 13028
rect 33872 13084 33936 13088
rect 33872 13028 33876 13084
rect 33876 13028 33932 13084
rect 33932 13028 33936 13084
rect 33872 13024 33936 13028
rect 33952 13084 34016 13088
rect 33952 13028 33956 13084
rect 33956 13028 34012 13084
rect 34012 13028 34016 13084
rect 33952 13024 34016 13028
rect 34032 13084 34096 13088
rect 34032 13028 34036 13084
rect 34036 13028 34092 13084
rect 34092 13028 34096 13084
rect 34032 13024 34096 13028
rect 44739 13084 44803 13088
rect 44739 13028 44743 13084
rect 44743 13028 44799 13084
rect 44799 13028 44803 13084
rect 44739 13024 44803 13028
rect 44819 13084 44883 13088
rect 44819 13028 44823 13084
rect 44823 13028 44879 13084
rect 44879 13028 44883 13084
rect 44819 13024 44883 13028
rect 44899 13084 44963 13088
rect 44899 13028 44903 13084
rect 44903 13028 44959 13084
rect 44959 13028 44963 13084
rect 44899 13024 44963 13028
rect 44979 13084 45043 13088
rect 44979 13028 44983 13084
rect 44983 13028 45039 13084
rect 45039 13028 45043 13084
rect 44979 13024 45043 13028
rect 6425 12540 6489 12544
rect 6425 12484 6429 12540
rect 6429 12484 6485 12540
rect 6485 12484 6489 12540
rect 6425 12480 6489 12484
rect 6505 12540 6569 12544
rect 6505 12484 6509 12540
rect 6509 12484 6565 12540
rect 6565 12484 6569 12540
rect 6505 12480 6569 12484
rect 6585 12540 6649 12544
rect 6585 12484 6589 12540
rect 6589 12484 6645 12540
rect 6645 12484 6649 12540
rect 6585 12480 6649 12484
rect 6665 12540 6729 12544
rect 6665 12484 6669 12540
rect 6669 12484 6725 12540
rect 6725 12484 6729 12540
rect 6665 12480 6729 12484
rect 17372 12540 17436 12544
rect 17372 12484 17376 12540
rect 17376 12484 17432 12540
rect 17432 12484 17436 12540
rect 17372 12480 17436 12484
rect 17452 12540 17516 12544
rect 17452 12484 17456 12540
rect 17456 12484 17512 12540
rect 17512 12484 17516 12540
rect 17452 12480 17516 12484
rect 17532 12540 17596 12544
rect 17532 12484 17536 12540
rect 17536 12484 17592 12540
rect 17592 12484 17596 12540
rect 17532 12480 17596 12484
rect 17612 12540 17676 12544
rect 17612 12484 17616 12540
rect 17616 12484 17672 12540
rect 17672 12484 17676 12540
rect 17612 12480 17676 12484
rect 28319 12540 28383 12544
rect 28319 12484 28323 12540
rect 28323 12484 28379 12540
rect 28379 12484 28383 12540
rect 28319 12480 28383 12484
rect 28399 12540 28463 12544
rect 28399 12484 28403 12540
rect 28403 12484 28459 12540
rect 28459 12484 28463 12540
rect 28399 12480 28463 12484
rect 28479 12540 28543 12544
rect 28479 12484 28483 12540
rect 28483 12484 28539 12540
rect 28539 12484 28543 12540
rect 28479 12480 28543 12484
rect 28559 12540 28623 12544
rect 28559 12484 28563 12540
rect 28563 12484 28619 12540
rect 28619 12484 28623 12540
rect 28559 12480 28623 12484
rect 39266 12540 39330 12544
rect 39266 12484 39270 12540
rect 39270 12484 39326 12540
rect 39326 12484 39330 12540
rect 39266 12480 39330 12484
rect 39346 12540 39410 12544
rect 39346 12484 39350 12540
rect 39350 12484 39406 12540
rect 39406 12484 39410 12540
rect 39346 12480 39410 12484
rect 39426 12540 39490 12544
rect 39426 12484 39430 12540
rect 39430 12484 39486 12540
rect 39486 12484 39490 12540
rect 39426 12480 39490 12484
rect 39506 12540 39570 12544
rect 39506 12484 39510 12540
rect 39510 12484 39566 12540
rect 39566 12484 39570 12540
rect 39506 12480 39570 12484
rect 11898 11996 11962 12000
rect 11898 11940 11902 11996
rect 11902 11940 11958 11996
rect 11958 11940 11962 11996
rect 11898 11936 11962 11940
rect 11978 11996 12042 12000
rect 11978 11940 11982 11996
rect 11982 11940 12038 11996
rect 12038 11940 12042 11996
rect 11978 11936 12042 11940
rect 12058 11996 12122 12000
rect 12058 11940 12062 11996
rect 12062 11940 12118 11996
rect 12118 11940 12122 11996
rect 12058 11936 12122 11940
rect 12138 11996 12202 12000
rect 12138 11940 12142 11996
rect 12142 11940 12198 11996
rect 12198 11940 12202 11996
rect 12138 11936 12202 11940
rect 22845 11996 22909 12000
rect 22845 11940 22849 11996
rect 22849 11940 22905 11996
rect 22905 11940 22909 11996
rect 22845 11936 22909 11940
rect 22925 11996 22989 12000
rect 22925 11940 22929 11996
rect 22929 11940 22985 11996
rect 22985 11940 22989 11996
rect 22925 11936 22989 11940
rect 23005 11996 23069 12000
rect 23005 11940 23009 11996
rect 23009 11940 23065 11996
rect 23065 11940 23069 11996
rect 23005 11936 23069 11940
rect 23085 11996 23149 12000
rect 23085 11940 23089 11996
rect 23089 11940 23145 11996
rect 23145 11940 23149 11996
rect 23085 11936 23149 11940
rect 33792 11996 33856 12000
rect 33792 11940 33796 11996
rect 33796 11940 33852 11996
rect 33852 11940 33856 11996
rect 33792 11936 33856 11940
rect 33872 11996 33936 12000
rect 33872 11940 33876 11996
rect 33876 11940 33932 11996
rect 33932 11940 33936 11996
rect 33872 11936 33936 11940
rect 33952 11996 34016 12000
rect 33952 11940 33956 11996
rect 33956 11940 34012 11996
rect 34012 11940 34016 11996
rect 33952 11936 34016 11940
rect 34032 11996 34096 12000
rect 34032 11940 34036 11996
rect 34036 11940 34092 11996
rect 34092 11940 34096 11996
rect 34032 11936 34096 11940
rect 44739 11996 44803 12000
rect 44739 11940 44743 11996
rect 44743 11940 44799 11996
rect 44799 11940 44803 11996
rect 44739 11936 44803 11940
rect 44819 11996 44883 12000
rect 44819 11940 44823 11996
rect 44823 11940 44879 11996
rect 44879 11940 44883 11996
rect 44819 11936 44883 11940
rect 44899 11996 44963 12000
rect 44899 11940 44903 11996
rect 44903 11940 44959 11996
rect 44959 11940 44963 11996
rect 44899 11936 44963 11940
rect 44979 11996 45043 12000
rect 44979 11940 44983 11996
rect 44983 11940 45039 11996
rect 45039 11940 45043 11996
rect 44979 11936 45043 11940
rect 6425 11452 6489 11456
rect 6425 11396 6429 11452
rect 6429 11396 6485 11452
rect 6485 11396 6489 11452
rect 6425 11392 6489 11396
rect 6505 11452 6569 11456
rect 6505 11396 6509 11452
rect 6509 11396 6565 11452
rect 6565 11396 6569 11452
rect 6505 11392 6569 11396
rect 6585 11452 6649 11456
rect 6585 11396 6589 11452
rect 6589 11396 6645 11452
rect 6645 11396 6649 11452
rect 6585 11392 6649 11396
rect 6665 11452 6729 11456
rect 6665 11396 6669 11452
rect 6669 11396 6725 11452
rect 6725 11396 6729 11452
rect 6665 11392 6729 11396
rect 17372 11452 17436 11456
rect 17372 11396 17376 11452
rect 17376 11396 17432 11452
rect 17432 11396 17436 11452
rect 17372 11392 17436 11396
rect 17452 11452 17516 11456
rect 17452 11396 17456 11452
rect 17456 11396 17512 11452
rect 17512 11396 17516 11452
rect 17452 11392 17516 11396
rect 17532 11452 17596 11456
rect 17532 11396 17536 11452
rect 17536 11396 17592 11452
rect 17592 11396 17596 11452
rect 17532 11392 17596 11396
rect 17612 11452 17676 11456
rect 17612 11396 17616 11452
rect 17616 11396 17672 11452
rect 17672 11396 17676 11452
rect 17612 11392 17676 11396
rect 28319 11452 28383 11456
rect 28319 11396 28323 11452
rect 28323 11396 28379 11452
rect 28379 11396 28383 11452
rect 28319 11392 28383 11396
rect 28399 11452 28463 11456
rect 28399 11396 28403 11452
rect 28403 11396 28459 11452
rect 28459 11396 28463 11452
rect 28399 11392 28463 11396
rect 28479 11452 28543 11456
rect 28479 11396 28483 11452
rect 28483 11396 28539 11452
rect 28539 11396 28543 11452
rect 28479 11392 28543 11396
rect 28559 11452 28623 11456
rect 28559 11396 28563 11452
rect 28563 11396 28619 11452
rect 28619 11396 28623 11452
rect 28559 11392 28623 11396
rect 39266 11452 39330 11456
rect 39266 11396 39270 11452
rect 39270 11396 39326 11452
rect 39326 11396 39330 11452
rect 39266 11392 39330 11396
rect 39346 11452 39410 11456
rect 39346 11396 39350 11452
rect 39350 11396 39406 11452
rect 39406 11396 39410 11452
rect 39346 11392 39410 11396
rect 39426 11452 39490 11456
rect 39426 11396 39430 11452
rect 39430 11396 39486 11452
rect 39486 11396 39490 11452
rect 39426 11392 39490 11396
rect 39506 11452 39570 11456
rect 39506 11396 39510 11452
rect 39510 11396 39566 11452
rect 39566 11396 39570 11452
rect 39506 11392 39570 11396
rect 11898 10908 11962 10912
rect 11898 10852 11902 10908
rect 11902 10852 11958 10908
rect 11958 10852 11962 10908
rect 11898 10848 11962 10852
rect 11978 10908 12042 10912
rect 11978 10852 11982 10908
rect 11982 10852 12038 10908
rect 12038 10852 12042 10908
rect 11978 10848 12042 10852
rect 12058 10908 12122 10912
rect 12058 10852 12062 10908
rect 12062 10852 12118 10908
rect 12118 10852 12122 10908
rect 12058 10848 12122 10852
rect 12138 10908 12202 10912
rect 12138 10852 12142 10908
rect 12142 10852 12198 10908
rect 12198 10852 12202 10908
rect 12138 10848 12202 10852
rect 22845 10908 22909 10912
rect 22845 10852 22849 10908
rect 22849 10852 22905 10908
rect 22905 10852 22909 10908
rect 22845 10848 22909 10852
rect 22925 10908 22989 10912
rect 22925 10852 22929 10908
rect 22929 10852 22985 10908
rect 22985 10852 22989 10908
rect 22925 10848 22989 10852
rect 23005 10908 23069 10912
rect 23005 10852 23009 10908
rect 23009 10852 23065 10908
rect 23065 10852 23069 10908
rect 23005 10848 23069 10852
rect 23085 10908 23149 10912
rect 23085 10852 23089 10908
rect 23089 10852 23145 10908
rect 23145 10852 23149 10908
rect 23085 10848 23149 10852
rect 33792 10908 33856 10912
rect 33792 10852 33796 10908
rect 33796 10852 33852 10908
rect 33852 10852 33856 10908
rect 33792 10848 33856 10852
rect 33872 10908 33936 10912
rect 33872 10852 33876 10908
rect 33876 10852 33932 10908
rect 33932 10852 33936 10908
rect 33872 10848 33936 10852
rect 33952 10908 34016 10912
rect 33952 10852 33956 10908
rect 33956 10852 34012 10908
rect 34012 10852 34016 10908
rect 33952 10848 34016 10852
rect 34032 10908 34096 10912
rect 34032 10852 34036 10908
rect 34036 10852 34092 10908
rect 34092 10852 34096 10908
rect 34032 10848 34096 10852
rect 44739 10908 44803 10912
rect 44739 10852 44743 10908
rect 44743 10852 44799 10908
rect 44799 10852 44803 10908
rect 44739 10848 44803 10852
rect 44819 10908 44883 10912
rect 44819 10852 44823 10908
rect 44823 10852 44879 10908
rect 44879 10852 44883 10908
rect 44819 10848 44883 10852
rect 44899 10908 44963 10912
rect 44899 10852 44903 10908
rect 44903 10852 44959 10908
rect 44959 10852 44963 10908
rect 44899 10848 44963 10852
rect 44979 10908 45043 10912
rect 44979 10852 44983 10908
rect 44983 10852 45039 10908
rect 45039 10852 45043 10908
rect 44979 10848 45043 10852
rect 6425 10364 6489 10368
rect 6425 10308 6429 10364
rect 6429 10308 6485 10364
rect 6485 10308 6489 10364
rect 6425 10304 6489 10308
rect 6505 10364 6569 10368
rect 6505 10308 6509 10364
rect 6509 10308 6565 10364
rect 6565 10308 6569 10364
rect 6505 10304 6569 10308
rect 6585 10364 6649 10368
rect 6585 10308 6589 10364
rect 6589 10308 6645 10364
rect 6645 10308 6649 10364
rect 6585 10304 6649 10308
rect 6665 10364 6729 10368
rect 6665 10308 6669 10364
rect 6669 10308 6725 10364
rect 6725 10308 6729 10364
rect 6665 10304 6729 10308
rect 17372 10364 17436 10368
rect 17372 10308 17376 10364
rect 17376 10308 17432 10364
rect 17432 10308 17436 10364
rect 17372 10304 17436 10308
rect 17452 10364 17516 10368
rect 17452 10308 17456 10364
rect 17456 10308 17512 10364
rect 17512 10308 17516 10364
rect 17452 10304 17516 10308
rect 17532 10364 17596 10368
rect 17532 10308 17536 10364
rect 17536 10308 17592 10364
rect 17592 10308 17596 10364
rect 17532 10304 17596 10308
rect 17612 10364 17676 10368
rect 17612 10308 17616 10364
rect 17616 10308 17672 10364
rect 17672 10308 17676 10364
rect 17612 10304 17676 10308
rect 28319 10364 28383 10368
rect 28319 10308 28323 10364
rect 28323 10308 28379 10364
rect 28379 10308 28383 10364
rect 28319 10304 28383 10308
rect 28399 10364 28463 10368
rect 28399 10308 28403 10364
rect 28403 10308 28459 10364
rect 28459 10308 28463 10364
rect 28399 10304 28463 10308
rect 28479 10364 28543 10368
rect 28479 10308 28483 10364
rect 28483 10308 28539 10364
rect 28539 10308 28543 10364
rect 28479 10304 28543 10308
rect 28559 10364 28623 10368
rect 28559 10308 28563 10364
rect 28563 10308 28619 10364
rect 28619 10308 28623 10364
rect 28559 10304 28623 10308
rect 39266 10364 39330 10368
rect 39266 10308 39270 10364
rect 39270 10308 39326 10364
rect 39326 10308 39330 10364
rect 39266 10304 39330 10308
rect 39346 10364 39410 10368
rect 39346 10308 39350 10364
rect 39350 10308 39406 10364
rect 39406 10308 39410 10364
rect 39346 10304 39410 10308
rect 39426 10364 39490 10368
rect 39426 10308 39430 10364
rect 39430 10308 39486 10364
rect 39486 10308 39490 10364
rect 39426 10304 39490 10308
rect 39506 10364 39570 10368
rect 39506 10308 39510 10364
rect 39510 10308 39566 10364
rect 39566 10308 39570 10364
rect 39506 10304 39570 10308
rect 11898 9820 11962 9824
rect 11898 9764 11902 9820
rect 11902 9764 11958 9820
rect 11958 9764 11962 9820
rect 11898 9760 11962 9764
rect 11978 9820 12042 9824
rect 11978 9764 11982 9820
rect 11982 9764 12038 9820
rect 12038 9764 12042 9820
rect 11978 9760 12042 9764
rect 12058 9820 12122 9824
rect 12058 9764 12062 9820
rect 12062 9764 12118 9820
rect 12118 9764 12122 9820
rect 12058 9760 12122 9764
rect 12138 9820 12202 9824
rect 12138 9764 12142 9820
rect 12142 9764 12198 9820
rect 12198 9764 12202 9820
rect 12138 9760 12202 9764
rect 22845 9820 22909 9824
rect 22845 9764 22849 9820
rect 22849 9764 22905 9820
rect 22905 9764 22909 9820
rect 22845 9760 22909 9764
rect 22925 9820 22989 9824
rect 22925 9764 22929 9820
rect 22929 9764 22985 9820
rect 22985 9764 22989 9820
rect 22925 9760 22989 9764
rect 23005 9820 23069 9824
rect 23005 9764 23009 9820
rect 23009 9764 23065 9820
rect 23065 9764 23069 9820
rect 23005 9760 23069 9764
rect 23085 9820 23149 9824
rect 23085 9764 23089 9820
rect 23089 9764 23145 9820
rect 23145 9764 23149 9820
rect 23085 9760 23149 9764
rect 33792 9820 33856 9824
rect 33792 9764 33796 9820
rect 33796 9764 33852 9820
rect 33852 9764 33856 9820
rect 33792 9760 33856 9764
rect 33872 9820 33936 9824
rect 33872 9764 33876 9820
rect 33876 9764 33932 9820
rect 33932 9764 33936 9820
rect 33872 9760 33936 9764
rect 33952 9820 34016 9824
rect 33952 9764 33956 9820
rect 33956 9764 34012 9820
rect 34012 9764 34016 9820
rect 33952 9760 34016 9764
rect 34032 9820 34096 9824
rect 34032 9764 34036 9820
rect 34036 9764 34092 9820
rect 34092 9764 34096 9820
rect 34032 9760 34096 9764
rect 44739 9820 44803 9824
rect 44739 9764 44743 9820
rect 44743 9764 44799 9820
rect 44799 9764 44803 9820
rect 44739 9760 44803 9764
rect 44819 9820 44883 9824
rect 44819 9764 44823 9820
rect 44823 9764 44879 9820
rect 44879 9764 44883 9820
rect 44819 9760 44883 9764
rect 44899 9820 44963 9824
rect 44899 9764 44903 9820
rect 44903 9764 44959 9820
rect 44959 9764 44963 9820
rect 44899 9760 44963 9764
rect 44979 9820 45043 9824
rect 44979 9764 44983 9820
rect 44983 9764 45039 9820
rect 45039 9764 45043 9820
rect 44979 9760 45043 9764
rect 6425 9276 6489 9280
rect 6425 9220 6429 9276
rect 6429 9220 6485 9276
rect 6485 9220 6489 9276
rect 6425 9216 6489 9220
rect 6505 9276 6569 9280
rect 6505 9220 6509 9276
rect 6509 9220 6565 9276
rect 6565 9220 6569 9276
rect 6505 9216 6569 9220
rect 6585 9276 6649 9280
rect 6585 9220 6589 9276
rect 6589 9220 6645 9276
rect 6645 9220 6649 9276
rect 6585 9216 6649 9220
rect 6665 9276 6729 9280
rect 6665 9220 6669 9276
rect 6669 9220 6725 9276
rect 6725 9220 6729 9276
rect 6665 9216 6729 9220
rect 17372 9276 17436 9280
rect 17372 9220 17376 9276
rect 17376 9220 17432 9276
rect 17432 9220 17436 9276
rect 17372 9216 17436 9220
rect 17452 9276 17516 9280
rect 17452 9220 17456 9276
rect 17456 9220 17512 9276
rect 17512 9220 17516 9276
rect 17452 9216 17516 9220
rect 17532 9276 17596 9280
rect 17532 9220 17536 9276
rect 17536 9220 17592 9276
rect 17592 9220 17596 9276
rect 17532 9216 17596 9220
rect 17612 9276 17676 9280
rect 17612 9220 17616 9276
rect 17616 9220 17672 9276
rect 17672 9220 17676 9276
rect 17612 9216 17676 9220
rect 28319 9276 28383 9280
rect 28319 9220 28323 9276
rect 28323 9220 28379 9276
rect 28379 9220 28383 9276
rect 28319 9216 28383 9220
rect 28399 9276 28463 9280
rect 28399 9220 28403 9276
rect 28403 9220 28459 9276
rect 28459 9220 28463 9276
rect 28399 9216 28463 9220
rect 28479 9276 28543 9280
rect 28479 9220 28483 9276
rect 28483 9220 28539 9276
rect 28539 9220 28543 9276
rect 28479 9216 28543 9220
rect 28559 9276 28623 9280
rect 28559 9220 28563 9276
rect 28563 9220 28619 9276
rect 28619 9220 28623 9276
rect 28559 9216 28623 9220
rect 39266 9276 39330 9280
rect 39266 9220 39270 9276
rect 39270 9220 39326 9276
rect 39326 9220 39330 9276
rect 39266 9216 39330 9220
rect 39346 9276 39410 9280
rect 39346 9220 39350 9276
rect 39350 9220 39406 9276
rect 39406 9220 39410 9276
rect 39346 9216 39410 9220
rect 39426 9276 39490 9280
rect 39426 9220 39430 9276
rect 39430 9220 39486 9276
rect 39486 9220 39490 9276
rect 39426 9216 39490 9220
rect 39506 9276 39570 9280
rect 39506 9220 39510 9276
rect 39510 9220 39566 9276
rect 39566 9220 39570 9276
rect 39506 9216 39570 9220
rect 11898 8732 11962 8736
rect 11898 8676 11902 8732
rect 11902 8676 11958 8732
rect 11958 8676 11962 8732
rect 11898 8672 11962 8676
rect 11978 8732 12042 8736
rect 11978 8676 11982 8732
rect 11982 8676 12038 8732
rect 12038 8676 12042 8732
rect 11978 8672 12042 8676
rect 12058 8732 12122 8736
rect 12058 8676 12062 8732
rect 12062 8676 12118 8732
rect 12118 8676 12122 8732
rect 12058 8672 12122 8676
rect 12138 8732 12202 8736
rect 12138 8676 12142 8732
rect 12142 8676 12198 8732
rect 12198 8676 12202 8732
rect 12138 8672 12202 8676
rect 22845 8732 22909 8736
rect 22845 8676 22849 8732
rect 22849 8676 22905 8732
rect 22905 8676 22909 8732
rect 22845 8672 22909 8676
rect 22925 8732 22989 8736
rect 22925 8676 22929 8732
rect 22929 8676 22985 8732
rect 22985 8676 22989 8732
rect 22925 8672 22989 8676
rect 23005 8732 23069 8736
rect 23005 8676 23009 8732
rect 23009 8676 23065 8732
rect 23065 8676 23069 8732
rect 23005 8672 23069 8676
rect 23085 8732 23149 8736
rect 23085 8676 23089 8732
rect 23089 8676 23145 8732
rect 23145 8676 23149 8732
rect 23085 8672 23149 8676
rect 33792 8732 33856 8736
rect 33792 8676 33796 8732
rect 33796 8676 33852 8732
rect 33852 8676 33856 8732
rect 33792 8672 33856 8676
rect 33872 8732 33936 8736
rect 33872 8676 33876 8732
rect 33876 8676 33932 8732
rect 33932 8676 33936 8732
rect 33872 8672 33936 8676
rect 33952 8732 34016 8736
rect 33952 8676 33956 8732
rect 33956 8676 34012 8732
rect 34012 8676 34016 8732
rect 33952 8672 34016 8676
rect 34032 8732 34096 8736
rect 34032 8676 34036 8732
rect 34036 8676 34092 8732
rect 34092 8676 34096 8732
rect 34032 8672 34096 8676
rect 44739 8732 44803 8736
rect 44739 8676 44743 8732
rect 44743 8676 44799 8732
rect 44799 8676 44803 8732
rect 44739 8672 44803 8676
rect 44819 8732 44883 8736
rect 44819 8676 44823 8732
rect 44823 8676 44879 8732
rect 44879 8676 44883 8732
rect 44819 8672 44883 8676
rect 44899 8732 44963 8736
rect 44899 8676 44903 8732
rect 44903 8676 44959 8732
rect 44959 8676 44963 8732
rect 44899 8672 44963 8676
rect 44979 8732 45043 8736
rect 44979 8676 44983 8732
rect 44983 8676 45039 8732
rect 45039 8676 45043 8732
rect 44979 8672 45043 8676
rect 6425 8188 6489 8192
rect 6425 8132 6429 8188
rect 6429 8132 6485 8188
rect 6485 8132 6489 8188
rect 6425 8128 6489 8132
rect 6505 8188 6569 8192
rect 6505 8132 6509 8188
rect 6509 8132 6565 8188
rect 6565 8132 6569 8188
rect 6505 8128 6569 8132
rect 6585 8188 6649 8192
rect 6585 8132 6589 8188
rect 6589 8132 6645 8188
rect 6645 8132 6649 8188
rect 6585 8128 6649 8132
rect 6665 8188 6729 8192
rect 6665 8132 6669 8188
rect 6669 8132 6725 8188
rect 6725 8132 6729 8188
rect 6665 8128 6729 8132
rect 17372 8188 17436 8192
rect 17372 8132 17376 8188
rect 17376 8132 17432 8188
rect 17432 8132 17436 8188
rect 17372 8128 17436 8132
rect 17452 8188 17516 8192
rect 17452 8132 17456 8188
rect 17456 8132 17512 8188
rect 17512 8132 17516 8188
rect 17452 8128 17516 8132
rect 17532 8188 17596 8192
rect 17532 8132 17536 8188
rect 17536 8132 17592 8188
rect 17592 8132 17596 8188
rect 17532 8128 17596 8132
rect 17612 8188 17676 8192
rect 17612 8132 17616 8188
rect 17616 8132 17672 8188
rect 17672 8132 17676 8188
rect 17612 8128 17676 8132
rect 28319 8188 28383 8192
rect 28319 8132 28323 8188
rect 28323 8132 28379 8188
rect 28379 8132 28383 8188
rect 28319 8128 28383 8132
rect 28399 8188 28463 8192
rect 28399 8132 28403 8188
rect 28403 8132 28459 8188
rect 28459 8132 28463 8188
rect 28399 8128 28463 8132
rect 28479 8188 28543 8192
rect 28479 8132 28483 8188
rect 28483 8132 28539 8188
rect 28539 8132 28543 8188
rect 28479 8128 28543 8132
rect 28559 8188 28623 8192
rect 28559 8132 28563 8188
rect 28563 8132 28619 8188
rect 28619 8132 28623 8188
rect 28559 8128 28623 8132
rect 39266 8188 39330 8192
rect 39266 8132 39270 8188
rect 39270 8132 39326 8188
rect 39326 8132 39330 8188
rect 39266 8128 39330 8132
rect 39346 8188 39410 8192
rect 39346 8132 39350 8188
rect 39350 8132 39406 8188
rect 39406 8132 39410 8188
rect 39346 8128 39410 8132
rect 39426 8188 39490 8192
rect 39426 8132 39430 8188
rect 39430 8132 39486 8188
rect 39486 8132 39490 8188
rect 39426 8128 39490 8132
rect 39506 8188 39570 8192
rect 39506 8132 39510 8188
rect 39510 8132 39566 8188
rect 39566 8132 39570 8188
rect 39506 8128 39570 8132
rect 11898 7644 11962 7648
rect 11898 7588 11902 7644
rect 11902 7588 11958 7644
rect 11958 7588 11962 7644
rect 11898 7584 11962 7588
rect 11978 7644 12042 7648
rect 11978 7588 11982 7644
rect 11982 7588 12038 7644
rect 12038 7588 12042 7644
rect 11978 7584 12042 7588
rect 12058 7644 12122 7648
rect 12058 7588 12062 7644
rect 12062 7588 12118 7644
rect 12118 7588 12122 7644
rect 12058 7584 12122 7588
rect 12138 7644 12202 7648
rect 12138 7588 12142 7644
rect 12142 7588 12198 7644
rect 12198 7588 12202 7644
rect 12138 7584 12202 7588
rect 22845 7644 22909 7648
rect 22845 7588 22849 7644
rect 22849 7588 22905 7644
rect 22905 7588 22909 7644
rect 22845 7584 22909 7588
rect 22925 7644 22989 7648
rect 22925 7588 22929 7644
rect 22929 7588 22985 7644
rect 22985 7588 22989 7644
rect 22925 7584 22989 7588
rect 23005 7644 23069 7648
rect 23005 7588 23009 7644
rect 23009 7588 23065 7644
rect 23065 7588 23069 7644
rect 23005 7584 23069 7588
rect 23085 7644 23149 7648
rect 23085 7588 23089 7644
rect 23089 7588 23145 7644
rect 23145 7588 23149 7644
rect 23085 7584 23149 7588
rect 33792 7644 33856 7648
rect 33792 7588 33796 7644
rect 33796 7588 33852 7644
rect 33852 7588 33856 7644
rect 33792 7584 33856 7588
rect 33872 7644 33936 7648
rect 33872 7588 33876 7644
rect 33876 7588 33932 7644
rect 33932 7588 33936 7644
rect 33872 7584 33936 7588
rect 33952 7644 34016 7648
rect 33952 7588 33956 7644
rect 33956 7588 34012 7644
rect 34012 7588 34016 7644
rect 33952 7584 34016 7588
rect 34032 7644 34096 7648
rect 34032 7588 34036 7644
rect 34036 7588 34092 7644
rect 34092 7588 34096 7644
rect 34032 7584 34096 7588
rect 44739 7644 44803 7648
rect 44739 7588 44743 7644
rect 44743 7588 44799 7644
rect 44799 7588 44803 7644
rect 44739 7584 44803 7588
rect 44819 7644 44883 7648
rect 44819 7588 44823 7644
rect 44823 7588 44879 7644
rect 44879 7588 44883 7644
rect 44819 7584 44883 7588
rect 44899 7644 44963 7648
rect 44899 7588 44903 7644
rect 44903 7588 44959 7644
rect 44959 7588 44963 7644
rect 44899 7584 44963 7588
rect 44979 7644 45043 7648
rect 44979 7588 44983 7644
rect 44983 7588 45039 7644
rect 45039 7588 45043 7644
rect 44979 7584 45043 7588
rect 6425 7100 6489 7104
rect 6425 7044 6429 7100
rect 6429 7044 6485 7100
rect 6485 7044 6489 7100
rect 6425 7040 6489 7044
rect 6505 7100 6569 7104
rect 6505 7044 6509 7100
rect 6509 7044 6565 7100
rect 6565 7044 6569 7100
rect 6505 7040 6569 7044
rect 6585 7100 6649 7104
rect 6585 7044 6589 7100
rect 6589 7044 6645 7100
rect 6645 7044 6649 7100
rect 6585 7040 6649 7044
rect 6665 7100 6729 7104
rect 6665 7044 6669 7100
rect 6669 7044 6725 7100
rect 6725 7044 6729 7100
rect 6665 7040 6729 7044
rect 17372 7100 17436 7104
rect 17372 7044 17376 7100
rect 17376 7044 17432 7100
rect 17432 7044 17436 7100
rect 17372 7040 17436 7044
rect 17452 7100 17516 7104
rect 17452 7044 17456 7100
rect 17456 7044 17512 7100
rect 17512 7044 17516 7100
rect 17452 7040 17516 7044
rect 17532 7100 17596 7104
rect 17532 7044 17536 7100
rect 17536 7044 17592 7100
rect 17592 7044 17596 7100
rect 17532 7040 17596 7044
rect 17612 7100 17676 7104
rect 17612 7044 17616 7100
rect 17616 7044 17672 7100
rect 17672 7044 17676 7100
rect 17612 7040 17676 7044
rect 28319 7100 28383 7104
rect 28319 7044 28323 7100
rect 28323 7044 28379 7100
rect 28379 7044 28383 7100
rect 28319 7040 28383 7044
rect 28399 7100 28463 7104
rect 28399 7044 28403 7100
rect 28403 7044 28459 7100
rect 28459 7044 28463 7100
rect 28399 7040 28463 7044
rect 28479 7100 28543 7104
rect 28479 7044 28483 7100
rect 28483 7044 28539 7100
rect 28539 7044 28543 7100
rect 28479 7040 28543 7044
rect 28559 7100 28623 7104
rect 28559 7044 28563 7100
rect 28563 7044 28619 7100
rect 28619 7044 28623 7100
rect 28559 7040 28623 7044
rect 39266 7100 39330 7104
rect 39266 7044 39270 7100
rect 39270 7044 39326 7100
rect 39326 7044 39330 7100
rect 39266 7040 39330 7044
rect 39346 7100 39410 7104
rect 39346 7044 39350 7100
rect 39350 7044 39406 7100
rect 39406 7044 39410 7100
rect 39346 7040 39410 7044
rect 39426 7100 39490 7104
rect 39426 7044 39430 7100
rect 39430 7044 39486 7100
rect 39486 7044 39490 7100
rect 39426 7040 39490 7044
rect 39506 7100 39570 7104
rect 39506 7044 39510 7100
rect 39510 7044 39566 7100
rect 39566 7044 39570 7100
rect 39506 7040 39570 7044
rect 11898 6556 11962 6560
rect 11898 6500 11902 6556
rect 11902 6500 11958 6556
rect 11958 6500 11962 6556
rect 11898 6496 11962 6500
rect 11978 6556 12042 6560
rect 11978 6500 11982 6556
rect 11982 6500 12038 6556
rect 12038 6500 12042 6556
rect 11978 6496 12042 6500
rect 12058 6556 12122 6560
rect 12058 6500 12062 6556
rect 12062 6500 12118 6556
rect 12118 6500 12122 6556
rect 12058 6496 12122 6500
rect 12138 6556 12202 6560
rect 12138 6500 12142 6556
rect 12142 6500 12198 6556
rect 12198 6500 12202 6556
rect 12138 6496 12202 6500
rect 22845 6556 22909 6560
rect 22845 6500 22849 6556
rect 22849 6500 22905 6556
rect 22905 6500 22909 6556
rect 22845 6496 22909 6500
rect 22925 6556 22989 6560
rect 22925 6500 22929 6556
rect 22929 6500 22985 6556
rect 22985 6500 22989 6556
rect 22925 6496 22989 6500
rect 23005 6556 23069 6560
rect 23005 6500 23009 6556
rect 23009 6500 23065 6556
rect 23065 6500 23069 6556
rect 23005 6496 23069 6500
rect 23085 6556 23149 6560
rect 23085 6500 23089 6556
rect 23089 6500 23145 6556
rect 23145 6500 23149 6556
rect 23085 6496 23149 6500
rect 33792 6556 33856 6560
rect 33792 6500 33796 6556
rect 33796 6500 33852 6556
rect 33852 6500 33856 6556
rect 33792 6496 33856 6500
rect 33872 6556 33936 6560
rect 33872 6500 33876 6556
rect 33876 6500 33932 6556
rect 33932 6500 33936 6556
rect 33872 6496 33936 6500
rect 33952 6556 34016 6560
rect 33952 6500 33956 6556
rect 33956 6500 34012 6556
rect 34012 6500 34016 6556
rect 33952 6496 34016 6500
rect 34032 6556 34096 6560
rect 34032 6500 34036 6556
rect 34036 6500 34092 6556
rect 34092 6500 34096 6556
rect 34032 6496 34096 6500
rect 44739 6556 44803 6560
rect 44739 6500 44743 6556
rect 44743 6500 44799 6556
rect 44799 6500 44803 6556
rect 44739 6496 44803 6500
rect 44819 6556 44883 6560
rect 44819 6500 44823 6556
rect 44823 6500 44879 6556
rect 44879 6500 44883 6556
rect 44819 6496 44883 6500
rect 44899 6556 44963 6560
rect 44899 6500 44903 6556
rect 44903 6500 44959 6556
rect 44959 6500 44963 6556
rect 44899 6496 44963 6500
rect 44979 6556 45043 6560
rect 44979 6500 44983 6556
rect 44983 6500 45039 6556
rect 45039 6500 45043 6556
rect 44979 6496 45043 6500
rect 6425 6012 6489 6016
rect 6425 5956 6429 6012
rect 6429 5956 6485 6012
rect 6485 5956 6489 6012
rect 6425 5952 6489 5956
rect 6505 6012 6569 6016
rect 6505 5956 6509 6012
rect 6509 5956 6565 6012
rect 6565 5956 6569 6012
rect 6505 5952 6569 5956
rect 6585 6012 6649 6016
rect 6585 5956 6589 6012
rect 6589 5956 6645 6012
rect 6645 5956 6649 6012
rect 6585 5952 6649 5956
rect 6665 6012 6729 6016
rect 6665 5956 6669 6012
rect 6669 5956 6725 6012
rect 6725 5956 6729 6012
rect 6665 5952 6729 5956
rect 17372 6012 17436 6016
rect 17372 5956 17376 6012
rect 17376 5956 17432 6012
rect 17432 5956 17436 6012
rect 17372 5952 17436 5956
rect 17452 6012 17516 6016
rect 17452 5956 17456 6012
rect 17456 5956 17512 6012
rect 17512 5956 17516 6012
rect 17452 5952 17516 5956
rect 17532 6012 17596 6016
rect 17532 5956 17536 6012
rect 17536 5956 17592 6012
rect 17592 5956 17596 6012
rect 17532 5952 17596 5956
rect 17612 6012 17676 6016
rect 17612 5956 17616 6012
rect 17616 5956 17672 6012
rect 17672 5956 17676 6012
rect 17612 5952 17676 5956
rect 28319 6012 28383 6016
rect 28319 5956 28323 6012
rect 28323 5956 28379 6012
rect 28379 5956 28383 6012
rect 28319 5952 28383 5956
rect 28399 6012 28463 6016
rect 28399 5956 28403 6012
rect 28403 5956 28459 6012
rect 28459 5956 28463 6012
rect 28399 5952 28463 5956
rect 28479 6012 28543 6016
rect 28479 5956 28483 6012
rect 28483 5956 28539 6012
rect 28539 5956 28543 6012
rect 28479 5952 28543 5956
rect 28559 6012 28623 6016
rect 28559 5956 28563 6012
rect 28563 5956 28619 6012
rect 28619 5956 28623 6012
rect 28559 5952 28623 5956
rect 39266 6012 39330 6016
rect 39266 5956 39270 6012
rect 39270 5956 39326 6012
rect 39326 5956 39330 6012
rect 39266 5952 39330 5956
rect 39346 6012 39410 6016
rect 39346 5956 39350 6012
rect 39350 5956 39406 6012
rect 39406 5956 39410 6012
rect 39346 5952 39410 5956
rect 39426 6012 39490 6016
rect 39426 5956 39430 6012
rect 39430 5956 39486 6012
rect 39486 5956 39490 6012
rect 39426 5952 39490 5956
rect 39506 6012 39570 6016
rect 39506 5956 39510 6012
rect 39510 5956 39566 6012
rect 39566 5956 39570 6012
rect 39506 5952 39570 5956
rect 11898 5468 11962 5472
rect 11898 5412 11902 5468
rect 11902 5412 11958 5468
rect 11958 5412 11962 5468
rect 11898 5408 11962 5412
rect 11978 5468 12042 5472
rect 11978 5412 11982 5468
rect 11982 5412 12038 5468
rect 12038 5412 12042 5468
rect 11978 5408 12042 5412
rect 12058 5468 12122 5472
rect 12058 5412 12062 5468
rect 12062 5412 12118 5468
rect 12118 5412 12122 5468
rect 12058 5408 12122 5412
rect 12138 5468 12202 5472
rect 12138 5412 12142 5468
rect 12142 5412 12198 5468
rect 12198 5412 12202 5468
rect 12138 5408 12202 5412
rect 22845 5468 22909 5472
rect 22845 5412 22849 5468
rect 22849 5412 22905 5468
rect 22905 5412 22909 5468
rect 22845 5408 22909 5412
rect 22925 5468 22989 5472
rect 22925 5412 22929 5468
rect 22929 5412 22985 5468
rect 22985 5412 22989 5468
rect 22925 5408 22989 5412
rect 23005 5468 23069 5472
rect 23005 5412 23009 5468
rect 23009 5412 23065 5468
rect 23065 5412 23069 5468
rect 23005 5408 23069 5412
rect 23085 5468 23149 5472
rect 23085 5412 23089 5468
rect 23089 5412 23145 5468
rect 23145 5412 23149 5468
rect 23085 5408 23149 5412
rect 33792 5468 33856 5472
rect 33792 5412 33796 5468
rect 33796 5412 33852 5468
rect 33852 5412 33856 5468
rect 33792 5408 33856 5412
rect 33872 5468 33936 5472
rect 33872 5412 33876 5468
rect 33876 5412 33932 5468
rect 33932 5412 33936 5468
rect 33872 5408 33936 5412
rect 33952 5468 34016 5472
rect 33952 5412 33956 5468
rect 33956 5412 34012 5468
rect 34012 5412 34016 5468
rect 33952 5408 34016 5412
rect 34032 5468 34096 5472
rect 34032 5412 34036 5468
rect 34036 5412 34092 5468
rect 34092 5412 34096 5468
rect 34032 5408 34096 5412
rect 44739 5468 44803 5472
rect 44739 5412 44743 5468
rect 44743 5412 44799 5468
rect 44799 5412 44803 5468
rect 44739 5408 44803 5412
rect 44819 5468 44883 5472
rect 44819 5412 44823 5468
rect 44823 5412 44879 5468
rect 44879 5412 44883 5468
rect 44819 5408 44883 5412
rect 44899 5468 44963 5472
rect 44899 5412 44903 5468
rect 44903 5412 44959 5468
rect 44959 5412 44963 5468
rect 44899 5408 44963 5412
rect 44979 5468 45043 5472
rect 44979 5412 44983 5468
rect 44983 5412 45039 5468
rect 45039 5412 45043 5468
rect 44979 5408 45043 5412
rect 6425 4924 6489 4928
rect 6425 4868 6429 4924
rect 6429 4868 6485 4924
rect 6485 4868 6489 4924
rect 6425 4864 6489 4868
rect 6505 4924 6569 4928
rect 6505 4868 6509 4924
rect 6509 4868 6565 4924
rect 6565 4868 6569 4924
rect 6505 4864 6569 4868
rect 6585 4924 6649 4928
rect 6585 4868 6589 4924
rect 6589 4868 6645 4924
rect 6645 4868 6649 4924
rect 6585 4864 6649 4868
rect 6665 4924 6729 4928
rect 6665 4868 6669 4924
rect 6669 4868 6725 4924
rect 6725 4868 6729 4924
rect 6665 4864 6729 4868
rect 17372 4924 17436 4928
rect 17372 4868 17376 4924
rect 17376 4868 17432 4924
rect 17432 4868 17436 4924
rect 17372 4864 17436 4868
rect 17452 4924 17516 4928
rect 17452 4868 17456 4924
rect 17456 4868 17512 4924
rect 17512 4868 17516 4924
rect 17452 4864 17516 4868
rect 17532 4924 17596 4928
rect 17532 4868 17536 4924
rect 17536 4868 17592 4924
rect 17592 4868 17596 4924
rect 17532 4864 17596 4868
rect 17612 4924 17676 4928
rect 17612 4868 17616 4924
rect 17616 4868 17672 4924
rect 17672 4868 17676 4924
rect 17612 4864 17676 4868
rect 28319 4924 28383 4928
rect 28319 4868 28323 4924
rect 28323 4868 28379 4924
rect 28379 4868 28383 4924
rect 28319 4864 28383 4868
rect 28399 4924 28463 4928
rect 28399 4868 28403 4924
rect 28403 4868 28459 4924
rect 28459 4868 28463 4924
rect 28399 4864 28463 4868
rect 28479 4924 28543 4928
rect 28479 4868 28483 4924
rect 28483 4868 28539 4924
rect 28539 4868 28543 4924
rect 28479 4864 28543 4868
rect 28559 4924 28623 4928
rect 28559 4868 28563 4924
rect 28563 4868 28619 4924
rect 28619 4868 28623 4924
rect 28559 4864 28623 4868
rect 39266 4924 39330 4928
rect 39266 4868 39270 4924
rect 39270 4868 39326 4924
rect 39326 4868 39330 4924
rect 39266 4864 39330 4868
rect 39346 4924 39410 4928
rect 39346 4868 39350 4924
rect 39350 4868 39406 4924
rect 39406 4868 39410 4924
rect 39346 4864 39410 4868
rect 39426 4924 39490 4928
rect 39426 4868 39430 4924
rect 39430 4868 39486 4924
rect 39486 4868 39490 4924
rect 39426 4864 39490 4868
rect 39506 4924 39570 4928
rect 39506 4868 39510 4924
rect 39510 4868 39566 4924
rect 39566 4868 39570 4924
rect 39506 4864 39570 4868
rect 11898 4380 11962 4384
rect 11898 4324 11902 4380
rect 11902 4324 11958 4380
rect 11958 4324 11962 4380
rect 11898 4320 11962 4324
rect 11978 4380 12042 4384
rect 11978 4324 11982 4380
rect 11982 4324 12038 4380
rect 12038 4324 12042 4380
rect 11978 4320 12042 4324
rect 12058 4380 12122 4384
rect 12058 4324 12062 4380
rect 12062 4324 12118 4380
rect 12118 4324 12122 4380
rect 12058 4320 12122 4324
rect 12138 4380 12202 4384
rect 12138 4324 12142 4380
rect 12142 4324 12198 4380
rect 12198 4324 12202 4380
rect 12138 4320 12202 4324
rect 22845 4380 22909 4384
rect 22845 4324 22849 4380
rect 22849 4324 22905 4380
rect 22905 4324 22909 4380
rect 22845 4320 22909 4324
rect 22925 4380 22989 4384
rect 22925 4324 22929 4380
rect 22929 4324 22985 4380
rect 22985 4324 22989 4380
rect 22925 4320 22989 4324
rect 23005 4380 23069 4384
rect 23005 4324 23009 4380
rect 23009 4324 23065 4380
rect 23065 4324 23069 4380
rect 23005 4320 23069 4324
rect 23085 4380 23149 4384
rect 23085 4324 23089 4380
rect 23089 4324 23145 4380
rect 23145 4324 23149 4380
rect 23085 4320 23149 4324
rect 33792 4380 33856 4384
rect 33792 4324 33796 4380
rect 33796 4324 33852 4380
rect 33852 4324 33856 4380
rect 33792 4320 33856 4324
rect 33872 4380 33936 4384
rect 33872 4324 33876 4380
rect 33876 4324 33932 4380
rect 33932 4324 33936 4380
rect 33872 4320 33936 4324
rect 33952 4380 34016 4384
rect 33952 4324 33956 4380
rect 33956 4324 34012 4380
rect 34012 4324 34016 4380
rect 33952 4320 34016 4324
rect 34032 4380 34096 4384
rect 34032 4324 34036 4380
rect 34036 4324 34092 4380
rect 34092 4324 34096 4380
rect 34032 4320 34096 4324
rect 44739 4380 44803 4384
rect 44739 4324 44743 4380
rect 44743 4324 44799 4380
rect 44799 4324 44803 4380
rect 44739 4320 44803 4324
rect 44819 4380 44883 4384
rect 44819 4324 44823 4380
rect 44823 4324 44879 4380
rect 44879 4324 44883 4380
rect 44819 4320 44883 4324
rect 44899 4380 44963 4384
rect 44899 4324 44903 4380
rect 44903 4324 44959 4380
rect 44959 4324 44963 4380
rect 44899 4320 44963 4324
rect 44979 4380 45043 4384
rect 44979 4324 44983 4380
rect 44983 4324 45039 4380
rect 45039 4324 45043 4380
rect 44979 4320 45043 4324
rect 6425 3836 6489 3840
rect 6425 3780 6429 3836
rect 6429 3780 6485 3836
rect 6485 3780 6489 3836
rect 6425 3776 6489 3780
rect 6505 3836 6569 3840
rect 6505 3780 6509 3836
rect 6509 3780 6565 3836
rect 6565 3780 6569 3836
rect 6505 3776 6569 3780
rect 6585 3836 6649 3840
rect 6585 3780 6589 3836
rect 6589 3780 6645 3836
rect 6645 3780 6649 3836
rect 6585 3776 6649 3780
rect 6665 3836 6729 3840
rect 6665 3780 6669 3836
rect 6669 3780 6725 3836
rect 6725 3780 6729 3836
rect 6665 3776 6729 3780
rect 17372 3836 17436 3840
rect 17372 3780 17376 3836
rect 17376 3780 17432 3836
rect 17432 3780 17436 3836
rect 17372 3776 17436 3780
rect 17452 3836 17516 3840
rect 17452 3780 17456 3836
rect 17456 3780 17512 3836
rect 17512 3780 17516 3836
rect 17452 3776 17516 3780
rect 17532 3836 17596 3840
rect 17532 3780 17536 3836
rect 17536 3780 17592 3836
rect 17592 3780 17596 3836
rect 17532 3776 17596 3780
rect 17612 3836 17676 3840
rect 17612 3780 17616 3836
rect 17616 3780 17672 3836
rect 17672 3780 17676 3836
rect 17612 3776 17676 3780
rect 28319 3836 28383 3840
rect 28319 3780 28323 3836
rect 28323 3780 28379 3836
rect 28379 3780 28383 3836
rect 28319 3776 28383 3780
rect 28399 3836 28463 3840
rect 28399 3780 28403 3836
rect 28403 3780 28459 3836
rect 28459 3780 28463 3836
rect 28399 3776 28463 3780
rect 28479 3836 28543 3840
rect 28479 3780 28483 3836
rect 28483 3780 28539 3836
rect 28539 3780 28543 3836
rect 28479 3776 28543 3780
rect 28559 3836 28623 3840
rect 28559 3780 28563 3836
rect 28563 3780 28619 3836
rect 28619 3780 28623 3836
rect 28559 3776 28623 3780
rect 39266 3836 39330 3840
rect 39266 3780 39270 3836
rect 39270 3780 39326 3836
rect 39326 3780 39330 3836
rect 39266 3776 39330 3780
rect 39346 3836 39410 3840
rect 39346 3780 39350 3836
rect 39350 3780 39406 3836
rect 39406 3780 39410 3836
rect 39346 3776 39410 3780
rect 39426 3836 39490 3840
rect 39426 3780 39430 3836
rect 39430 3780 39486 3836
rect 39486 3780 39490 3836
rect 39426 3776 39490 3780
rect 39506 3836 39570 3840
rect 39506 3780 39510 3836
rect 39510 3780 39566 3836
rect 39566 3780 39570 3836
rect 39506 3776 39570 3780
rect 11898 3292 11962 3296
rect 11898 3236 11902 3292
rect 11902 3236 11958 3292
rect 11958 3236 11962 3292
rect 11898 3232 11962 3236
rect 11978 3292 12042 3296
rect 11978 3236 11982 3292
rect 11982 3236 12038 3292
rect 12038 3236 12042 3292
rect 11978 3232 12042 3236
rect 12058 3292 12122 3296
rect 12058 3236 12062 3292
rect 12062 3236 12118 3292
rect 12118 3236 12122 3292
rect 12058 3232 12122 3236
rect 12138 3292 12202 3296
rect 12138 3236 12142 3292
rect 12142 3236 12198 3292
rect 12198 3236 12202 3292
rect 12138 3232 12202 3236
rect 22845 3292 22909 3296
rect 22845 3236 22849 3292
rect 22849 3236 22905 3292
rect 22905 3236 22909 3292
rect 22845 3232 22909 3236
rect 22925 3292 22989 3296
rect 22925 3236 22929 3292
rect 22929 3236 22985 3292
rect 22985 3236 22989 3292
rect 22925 3232 22989 3236
rect 23005 3292 23069 3296
rect 23005 3236 23009 3292
rect 23009 3236 23065 3292
rect 23065 3236 23069 3292
rect 23005 3232 23069 3236
rect 23085 3292 23149 3296
rect 23085 3236 23089 3292
rect 23089 3236 23145 3292
rect 23145 3236 23149 3292
rect 23085 3232 23149 3236
rect 33792 3292 33856 3296
rect 33792 3236 33796 3292
rect 33796 3236 33852 3292
rect 33852 3236 33856 3292
rect 33792 3232 33856 3236
rect 33872 3292 33936 3296
rect 33872 3236 33876 3292
rect 33876 3236 33932 3292
rect 33932 3236 33936 3292
rect 33872 3232 33936 3236
rect 33952 3292 34016 3296
rect 33952 3236 33956 3292
rect 33956 3236 34012 3292
rect 34012 3236 34016 3292
rect 33952 3232 34016 3236
rect 34032 3292 34096 3296
rect 34032 3236 34036 3292
rect 34036 3236 34092 3292
rect 34092 3236 34096 3292
rect 34032 3232 34096 3236
rect 44739 3292 44803 3296
rect 44739 3236 44743 3292
rect 44743 3236 44799 3292
rect 44799 3236 44803 3292
rect 44739 3232 44803 3236
rect 44819 3292 44883 3296
rect 44819 3236 44823 3292
rect 44823 3236 44879 3292
rect 44879 3236 44883 3292
rect 44819 3232 44883 3236
rect 44899 3292 44963 3296
rect 44899 3236 44903 3292
rect 44903 3236 44959 3292
rect 44959 3236 44963 3292
rect 44899 3232 44963 3236
rect 44979 3292 45043 3296
rect 44979 3236 44983 3292
rect 44983 3236 45039 3292
rect 45039 3236 45043 3292
rect 44979 3232 45043 3236
rect 6425 2748 6489 2752
rect 6425 2692 6429 2748
rect 6429 2692 6485 2748
rect 6485 2692 6489 2748
rect 6425 2688 6489 2692
rect 6505 2748 6569 2752
rect 6505 2692 6509 2748
rect 6509 2692 6565 2748
rect 6565 2692 6569 2748
rect 6505 2688 6569 2692
rect 6585 2748 6649 2752
rect 6585 2692 6589 2748
rect 6589 2692 6645 2748
rect 6645 2692 6649 2748
rect 6585 2688 6649 2692
rect 6665 2748 6729 2752
rect 6665 2692 6669 2748
rect 6669 2692 6725 2748
rect 6725 2692 6729 2748
rect 6665 2688 6729 2692
rect 17372 2748 17436 2752
rect 17372 2692 17376 2748
rect 17376 2692 17432 2748
rect 17432 2692 17436 2748
rect 17372 2688 17436 2692
rect 17452 2748 17516 2752
rect 17452 2692 17456 2748
rect 17456 2692 17512 2748
rect 17512 2692 17516 2748
rect 17452 2688 17516 2692
rect 17532 2748 17596 2752
rect 17532 2692 17536 2748
rect 17536 2692 17592 2748
rect 17592 2692 17596 2748
rect 17532 2688 17596 2692
rect 17612 2748 17676 2752
rect 17612 2692 17616 2748
rect 17616 2692 17672 2748
rect 17672 2692 17676 2748
rect 17612 2688 17676 2692
rect 28319 2748 28383 2752
rect 28319 2692 28323 2748
rect 28323 2692 28379 2748
rect 28379 2692 28383 2748
rect 28319 2688 28383 2692
rect 28399 2748 28463 2752
rect 28399 2692 28403 2748
rect 28403 2692 28459 2748
rect 28459 2692 28463 2748
rect 28399 2688 28463 2692
rect 28479 2748 28543 2752
rect 28479 2692 28483 2748
rect 28483 2692 28539 2748
rect 28539 2692 28543 2748
rect 28479 2688 28543 2692
rect 28559 2748 28623 2752
rect 28559 2692 28563 2748
rect 28563 2692 28619 2748
rect 28619 2692 28623 2748
rect 28559 2688 28623 2692
rect 39266 2748 39330 2752
rect 39266 2692 39270 2748
rect 39270 2692 39326 2748
rect 39326 2692 39330 2748
rect 39266 2688 39330 2692
rect 39346 2748 39410 2752
rect 39346 2692 39350 2748
rect 39350 2692 39406 2748
rect 39406 2692 39410 2748
rect 39346 2688 39410 2692
rect 39426 2748 39490 2752
rect 39426 2692 39430 2748
rect 39430 2692 39486 2748
rect 39486 2692 39490 2748
rect 39426 2688 39490 2692
rect 39506 2748 39570 2752
rect 39506 2692 39510 2748
rect 39510 2692 39566 2748
rect 39566 2692 39570 2748
rect 39506 2688 39570 2692
rect 11898 2204 11962 2208
rect 11898 2148 11902 2204
rect 11902 2148 11958 2204
rect 11958 2148 11962 2204
rect 11898 2144 11962 2148
rect 11978 2204 12042 2208
rect 11978 2148 11982 2204
rect 11982 2148 12038 2204
rect 12038 2148 12042 2204
rect 11978 2144 12042 2148
rect 12058 2204 12122 2208
rect 12058 2148 12062 2204
rect 12062 2148 12118 2204
rect 12118 2148 12122 2204
rect 12058 2144 12122 2148
rect 12138 2204 12202 2208
rect 12138 2148 12142 2204
rect 12142 2148 12198 2204
rect 12198 2148 12202 2204
rect 12138 2144 12202 2148
rect 22845 2204 22909 2208
rect 22845 2148 22849 2204
rect 22849 2148 22905 2204
rect 22905 2148 22909 2204
rect 22845 2144 22909 2148
rect 22925 2204 22989 2208
rect 22925 2148 22929 2204
rect 22929 2148 22985 2204
rect 22985 2148 22989 2204
rect 22925 2144 22989 2148
rect 23005 2204 23069 2208
rect 23005 2148 23009 2204
rect 23009 2148 23065 2204
rect 23065 2148 23069 2204
rect 23005 2144 23069 2148
rect 23085 2204 23149 2208
rect 23085 2148 23089 2204
rect 23089 2148 23145 2204
rect 23145 2148 23149 2204
rect 23085 2144 23149 2148
rect 33792 2204 33856 2208
rect 33792 2148 33796 2204
rect 33796 2148 33852 2204
rect 33852 2148 33856 2204
rect 33792 2144 33856 2148
rect 33872 2204 33936 2208
rect 33872 2148 33876 2204
rect 33876 2148 33932 2204
rect 33932 2148 33936 2204
rect 33872 2144 33936 2148
rect 33952 2204 34016 2208
rect 33952 2148 33956 2204
rect 33956 2148 34012 2204
rect 34012 2148 34016 2204
rect 33952 2144 34016 2148
rect 34032 2204 34096 2208
rect 34032 2148 34036 2204
rect 34036 2148 34092 2204
rect 34092 2148 34096 2204
rect 34032 2144 34096 2148
rect 44739 2204 44803 2208
rect 44739 2148 44743 2204
rect 44743 2148 44799 2204
rect 44799 2148 44803 2204
rect 44739 2144 44803 2148
rect 44819 2204 44883 2208
rect 44819 2148 44823 2204
rect 44823 2148 44879 2204
rect 44879 2148 44883 2204
rect 44819 2144 44883 2148
rect 44899 2204 44963 2208
rect 44899 2148 44903 2204
rect 44903 2148 44959 2204
rect 44959 2148 44963 2204
rect 44899 2144 44963 2148
rect 44979 2204 45043 2208
rect 44979 2148 44983 2204
rect 44983 2148 45039 2204
rect 45039 2148 45043 2204
rect 44979 2144 45043 2148
<< metal4 >>
rect 6417 16896 6737 17456
rect 6417 16832 6425 16896
rect 6489 16832 6505 16896
rect 6569 16832 6585 16896
rect 6649 16832 6665 16896
rect 6729 16832 6737 16896
rect 6417 15808 6737 16832
rect 6417 15744 6425 15808
rect 6489 15744 6505 15808
rect 6569 15744 6585 15808
rect 6649 15744 6665 15808
rect 6729 15744 6737 15808
rect 6417 14720 6737 15744
rect 6417 14656 6425 14720
rect 6489 14656 6505 14720
rect 6569 14656 6585 14720
rect 6649 14656 6665 14720
rect 6729 14656 6737 14720
rect 6417 13632 6737 14656
rect 6417 13568 6425 13632
rect 6489 13568 6505 13632
rect 6569 13568 6585 13632
rect 6649 13568 6665 13632
rect 6729 13568 6737 13632
rect 6417 12544 6737 13568
rect 6417 12480 6425 12544
rect 6489 12480 6505 12544
rect 6569 12480 6585 12544
rect 6649 12480 6665 12544
rect 6729 12480 6737 12544
rect 6417 11456 6737 12480
rect 6417 11392 6425 11456
rect 6489 11392 6505 11456
rect 6569 11392 6585 11456
rect 6649 11392 6665 11456
rect 6729 11392 6737 11456
rect 6417 10368 6737 11392
rect 6417 10304 6425 10368
rect 6489 10304 6505 10368
rect 6569 10304 6585 10368
rect 6649 10304 6665 10368
rect 6729 10304 6737 10368
rect 6417 9280 6737 10304
rect 6417 9216 6425 9280
rect 6489 9216 6505 9280
rect 6569 9216 6585 9280
rect 6649 9216 6665 9280
rect 6729 9216 6737 9280
rect 6417 8192 6737 9216
rect 6417 8128 6425 8192
rect 6489 8128 6505 8192
rect 6569 8128 6585 8192
rect 6649 8128 6665 8192
rect 6729 8128 6737 8192
rect 6417 7104 6737 8128
rect 6417 7040 6425 7104
rect 6489 7040 6505 7104
rect 6569 7040 6585 7104
rect 6649 7040 6665 7104
rect 6729 7040 6737 7104
rect 6417 6016 6737 7040
rect 6417 5952 6425 6016
rect 6489 5952 6505 6016
rect 6569 5952 6585 6016
rect 6649 5952 6665 6016
rect 6729 5952 6737 6016
rect 6417 4928 6737 5952
rect 6417 4864 6425 4928
rect 6489 4864 6505 4928
rect 6569 4864 6585 4928
rect 6649 4864 6665 4928
rect 6729 4864 6737 4928
rect 6417 3840 6737 4864
rect 6417 3776 6425 3840
rect 6489 3776 6505 3840
rect 6569 3776 6585 3840
rect 6649 3776 6665 3840
rect 6729 3776 6737 3840
rect 6417 2752 6737 3776
rect 6417 2688 6425 2752
rect 6489 2688 6505 2752
rect 6569 2688 6585 2752
rect 6649 2688 6665 2752
rect 6729 2688 6737 2752
rect 6417 2128 6737 2688
rect 11890 17440 12210 17456
rect 11890 17376 11898 17440
rect 11962 17376 11978 17440
rect 12042 17376 12058 17440
rect 12122 17376 12138 17440
rect 12202 17376 12210 17440
rect 11890 16352 12210 17376
rect 11890 16288 11898 16352
rect 11962 16288 11978 16352
rect 12042 16288 12058 16352
rect 12122 16288 12138 16352
rect 12202 16288 12210 16352
rect 11890 15264 12210 16288
rect 11890 15200 11898 15264
rect 11962 15200 11978 15264
rect 12042 15200 12058 15264
rect 12122 15200 12138 15264
rect 12202 15200 12210 15264
rect 11890 14176 12210 15200
rect 11890 14112 11898 14176
rect 11962 14112 11978 14176
rect 12042 14112 12058 14176
rect 12122 14112 12138 14176
rect 12202 14112 12210 14176
rect 11890 13088 12210 14112
rect 11890 13024 11898 13088
rect 11962 13024 11978 13088
rect 12042 13024 12058 13088
rect 12122 13024 12138 13088
rect 12202 13024 12210 13088
rect 11890 12000 12210 13024
rect 11890 11936 11898 12000
rect 11962 11936 11978 12000
rect 12042 11936 12058 12000
rect 12122 11936 12138 12000
rect 12202 11936 12210 12000
rect 11890 10912 12210 11936
rect 11890 10848 11898 10912
rect 11962 10848 11978 10912
rect 12042 10848 12058 10912
rect 12122 10848 12138 10912
rect 12202 10848 12210 10912
rect 11890 9824 12210 10848
rect 11890 9760 11898 9824
rect 11962 9760 11978 9824
rect 12042 9760 12058 9824
rect 12122 9760 12138 9824
rect 12202 9760 12210 9824
rect 11890 8736 12210 9760
rect 11890 8672 11898 8736
rect 11962 8672 11978 8736
rect 12042 8672 12058 8736
rect 12122 8672 12138 8736
rect 12202 8672 12210 8736
rect 11890 7648 12210 8672
rect 11890 7584 11898 7648
rect 11962 7584 11978 7648
rect 12042 7584 12058 7648
rect 12122 7584 12138 7648
rect 12202 7584 12210 7648
rect 11890 6560 12210 7584
rect 11890 6496 11898 6560
rect 11962 6496 11978 6560
rect 12042 6496 12058 6560
rect 12122 6496 12138 6560
rect 12202 6496 12210 6560
rect 11890 5472 12210 6496
rect 11890 5408 11898 5472
rect 11962 5408 11978 5472
rect 12042 5408 12058 5472
rect 12122 5408 12138 5472
rect 12202 5408 12210 5472
rect 11890 4384 12210 5408
rect 11890 4320 11898 4384
rect 11962 4320 11978 4384
rect 12042 4320 12058 4384
rect 12122 4320 12138 4384
rect 12202 4320 12210 4384
rect 11890 3296 12210 4320
rect 11890 3232 11898 3296
rect 11962 3232 11978 3296
rect 12042 3232 12058 3296
rect 12122 3232 12138 3296
rect 12202 3232 12210 3296
rect 11890 2208 12210 3232
rect 11890 2144 11898 2208
rect 11962 2144 11978 2208
rect 12042 2144 12058 2208
rect 12122 2144 12138 2208
rect 12202 2144 12210 2208
rect 11890 2128 12210 2144
rect 17364 16896 17684 17456
rect 17364 16832 17372 16896
rect 17436 16832 17452 16896
rect 17516 16832 17532 16896
rect 17596 16832 17612 16896
rect 17676 16832 17684 16896
rect 17364 15808 17684 16832
rect 17364 15744 17372 15808
rect 17436 15744 17452 15808
rect 17516 15744 17532 15808
rect 17596 15744 17612 15808
rect 17676 15744 17684 15808
rect 17364 14720 17684 15744
rect 17364 14656 17372 14720
rect 17436 14656 17452 14720
rect 17516 14656 17532 14720
rect 17596 14656 17612 14720
rect 17676 14656 17684 14720
rect 17364 13632 17684 14656
rect 17364 13568 17372 13632
rect 17436 13568 17452 13632
rect 17516 13568 17532 13632
rect 17596 13568 17612 13632
rect 17676 13568 17684 13632
rect 17364 12544 17684 13568
rect 17364 12480 17372 12544
rect 17436 12480 17452 12544
rect 17516 12480 17532 12544
rect 17596 12480 17612 12544
rect 17676 12480 17684 12544
rect 17364 11456 17684 12480
rect 17364 11392 17372 11456
rect 17436 11392 17452 11456
rect 17516 11392 17532 11456
rect 17596 11392 17612 11456
rect 17676 11392 17684 11456
rect 17364 10368 17684 11392
rect 17364 10304 17372 10368
rect 17436 10304 17452 10368
rect 17516 10304 17532 10368
rect 17596 10304 17612 10368
rect 17676 10304 17684 10368
rect 17364 9280 17684 10304
rect 17364 9216 17372 9280
rect 17436 9216 17452 9280
rect 17516 9216 17532 9280
rect 17596 9216 17612 9280
rect 17676 9216 17684 9280
rect 17364 8192 17684 9216
rect 17364 8128 17372 8192
rect 17436 8128 17452 8192
rect 17516 8128 17532 8192
rect 17596 8128 17612 8192
rect 17676 8128 17684 8192
rect 17364 7104 17684 8128
rect 17364 7040 17372 7104
rect 17436 7040 17452 7104
rect 17516 7040 17532 7104
rect 17596 7040 17612 7104
rect 17676 7040 17684 7104
rect 17364 6016 17684 7040
rect 17364 5952 17372 6016
rect 17436 5952 17452 6016
rect 17516 5952 17532 6016
rect 17596 5952 17612 6016
rect 17676 5952 17684 6016
rect 17364 4928 17684 5952
rect 17364 4864 17372 4928
rect 17436 4864 17452 4928
rect 17516 4864 17532 4928
rect 17596 4864 17612 4928
rect 17676 4864 17684 4928
rect 17364 3840 17684 4864
rect 17364 3776 17372 3840
rect 17436 3776 17452 3840
rect 17516 3776 17532 3840
rect 17596 3776 17612 3840
rect 17676 3776 17684 3840
rect 17364 2752 17684 3776
rect 17364 2688 17372 2752
rect 17436 2688 17452 2752
rect 17516 2688 17532 2752
rect 17596 2688 17612 2752
rect 17676 2688 17684 2752
rect 17364 2128 17684 2688
rect 22837 17440 23157 17456
rect 22837 17376 22845 17440
rect 22909 17376 22925 17440
rect 22989 17376 23005 17440
rect 23069 17376 23085 17440
rect 23149 17376 23157 17440
rect 22837 16352 23157 17376
rect 22837 16288 22845 16352
rect 22909 16288 22925 16352
rect 22989 16288 23005 16352
rect 23069 16288 23085 16352
rect 23149 16288 23157 16352
rect 22837 15264 23157 16288
rect 22837 15200 22845 15264
rect 22909 15200 22925 15264
rect 22989 15200 23005 15264
rect 23069 15200 23085 15264
rect 23149 15200 23157 15264
rect 22837 14176 23157 15200
rect 22837 14112 22845 14176
rect 22909 14112 22925 14176
rect 22989 14112 23005 14176
rect 23069 14112 23085 14176
rect 23149 14112 23157 14176
rect 22837 13088 23157 14112
rect 22837 13024 22845 13088
rect 22909 13024 22925 13088
rect 22989 13024 23005 13088
rect 23069 13024 23085 13088
rect 23149 13024 23157 13088
rect 22837 12000 23157 13024
rect 22837 11936 22845 12000
rect 22909 11936 22925 12000
rect 22989 11936 23005 12000
rect 23069 11936 23085 12000
rect 23149 11936 23157 12000
rect 22837 10912 23157 11936
rect 22837 10848 22845 10912
rect 22909 10848 22925 10912
rect 22989 10848 23005 10912
rect 23069 10848 23085 10912
rect 23149 10848 23157 10912
rect 22837 9824 23157 10848
rect 22837 9760 22845 9824
rect 22909 9760 22925 9824
rect 22989 9760 23005 9824
rect 23069 9760 23085 9824
rect 23149 9760 23157 9824
rect 22837 8736 23157 9760
rect 22837 8672 22845 8736
rect 22909 8672 22925 8736
rect 22989 8672 23005 8736
rect 23069 8672 23085 8736
rect 23149 8672 23157 8736
rect 22837 7648 23157 8672
rect 22837 7584 22845 7648
rect 22909 7584 22925 7648
rect 22989 7584 23005 7648
rect 23069 7584 23085 7648
rect 23149 7584 23157 7648
rect 22837 6560 23157 7584
rect 22837 6496 22845 6560
rect 22909 6496 22925 6560
rect 22989 6496 23005 6560
rect 23069 6496 23085 6560
rect 23149 6496 23157 6560
rect 22837 5472 23157 6496
rect 22837 5408 22845 5472
rect 22909 5408 22925 5472
rect 22989 5408 23005 5472
rect 23069 5408 23085 5472
rect 23149 5408 23157 5472
rect 22837 4384 23157 5408
rect 22837 4320 22845 4384
rect 22909 4320 22925 4384
rect 22989 4320 23005 4384
rect 23069 4320 23085 4384
rect 23149 4320 23157 4384
rect 22837 3296 23157 4320
rect 22837 3232 22845 3296
rect 22909 3232 22925 3296
rect 22989 3232 23005 3296
rect 23069 3232 23085 3296
rect 23149 3232 23157 3296
rect 22837 2208 23157 3232
rect 22837 2144 22845 2208
rect 22909 2144 22925 2208
rect 22989 2144 23005 2208
rect 23069 2144 23085 2208
rect 23149 2144 23157 2208
rect 22837 2128 23157 2144
rect 28311 16896 28631 17456
rect 28311 16832 28319 16896
rect 28383 16832 28399 16896
rect 28463 16832 28479 16896
rect 28543 16832 28559 16896
rect 28623 16832 28631 16896
rect 28311 15808 28631 16832
rect 28311 15744 28319 15808
rect 28383 15744 28399 15808
rect 28463 15744 28479 15808
rect 28543 15744 28559 15808
rect 28623 15744 28631 15808
rect 28311 14720 28631 15744
rect 28311 14656 28319 14720
rect 28383 14656 28399 14720
rect 28463 14656 28479 14720
rect 28543 14656 28559 14720
rect 28623 14656 28631 14720
rect 28311 13632 28631 14656
rect 28311 13568 28319 13632
rect 28383 13568 28399 13632
rect 28463 13568 28479 13632
rect 28543 13568 28559 13632
rect 28623 13568 28631 13632
rect 28311 12544 28631 13568
rect 28311 12480 28319 12544
rect 28383 12480 28399 12544
rect 28463 12480 28479 12544
rect 28543 12480 28559 12544
rect 28623 12480 28631 12544
rect 28311 11456 28631 12480
rect 28311 11392 28319 11456
rect 28383 11392 28399 11456
rect 28463 11392 28479 11456
rect 28543 11392 28559 11456
rect 28623 11392 28631 11456
rect 28311 10368 28631 11392
rect 28311 10304 28319 10368
rect 28383 10304 28399 10368
rect 28463 10304 28479 10368
rect 28543 10304 28559 10368
rect 28623 10304 28631 10368
rect 28311 9280 28631 10304
rect 28311 9216 28319 9280
rect 28383 9216 28399 9280
rect 28463 9216 28479 9280
rect 28543 9216 28559 9280
rect 28623 9216 28631 9280
rect 28311 8192 28631 9216
rect 28311 8128 28319 8192
rect 28383 8128 28399 8192
rect 28463 8128 28479 8192
rect 28543 8128 28559 8192
rect 28623 8128 28631 8192
rect 28311 7104 28631 8128
rect 28311 7040 28319 7104
rect 28383 7040 28399 7104
rect 28463 7040 28479 7104
rect 28543 7040 28559 7104
rect 28623 7040 28631 7104
rect 28311 6016 28631 7040
rect 28311 5952 28319 6016
rect 28383 5952 28399 6016
rect 28463 5952 28479 6016
rect 28543 5952 28559 6016
rect 28623 5952 28631 6016
rect 28311 4928 28631 5952
rect 28311 4864 28319 4928
rect 28383 4864 28399 4928
rect 28463 4864 28479 4928
rect 28543 4864 28559 4928
rect 28623 4864 28631 4928
rect 28311 3840 28631 4864
rect 28311 3776 28319 3840
rect 28383 3776 28399 3840
rect 28463 3776 28479 3840
rect 28543 3776 28559 3840
rect 28623 3776 28631 3840
rect 28311 2752 28631 3776
rect 28311 2688 28319 2752
rect 28383 2688 28399 2752
rect 28463 2688 28479 2752
rect 28543 2688 28559 2752
rect 28623 2688 28631 2752
rect 28311 2128 28631 2688
rect 33784 17440 34104 17456
rect 33784 17376 33792 17440
rect 33856 17376 33872 17440
rect 33936 17376 33952 17440
rect 34016 17376 34032 17440
rect 34096 17376 34104 17440
rect 33784 16352 34104 17376
rect 33784 16288 33792 16352
rect 33856 16288 33872 16352
rect 33936 16288 33952 16352
rect 34016 16288 34032 16352
rect 34096 16288 34104 16352
rect 33784 15264 34104 16288
rect 33784 15200 33792 15264
rect 33856 15200 33872 15264
rect 33936 15200 33952 15264
rect 34016 15200 34032 15264
rect 34096 15200 34104 15264
rect 33784 14176 34104 15200
rect 33784 14112 33792 14176
rect 33856 14112 33872 14176
rect 33936 14112 33952 14176
rect 34016 14112 34032 14176
rect 34096 14112 34104 14176
rect 33784 13088 34104 14112
rect 33784 13024 33792 13088
rect 33856 13024 33872 13088
rect 33936 13024 33952 13088
rect 34016 13024 34032 13088
rect 34096 13024 34104 13088
rect 33784 12000 34104 13024
rect 33784 11936 33792 12000
rect 33856 11936 33872 12000
rect 33936 11936 33952 12000
rect 34016 11936 34032 12000
rect 34096 11936 34104 12000
rect 33784 10912 34104 11936
rect 33784 10848 33792 10912
rect 33856 10848 33872 10912
rect 33936 10848 33952 10912
rect 34016 10848 34032 10912
rect 34096 10848 34104 10912
rect 33784 9824 34104 10848
rect 33784 9760 33792 9824
rect 33856 9760 33872 9824
rect 33936 9760 33952 9824
rect 34016 9760 34032 9824
rect 34096 9760 34104 9824
rect 33784 8736 34104 9760
rect 33784 8672 33792 8736
rect 33856 8672 33872 8736
rect 33936 8672 33952 8736
rect 34016 8672 34032 8736
rect 34096 8672 34104 8736
rect 33784 7648 34104 8672
rect 33784 7584 33792 7648
rect 33856 7584 33872 7648
rect 33936 7584 33952 7648
rect 34016 7584 34032 7648
rect 34096 7584 34104 7648
rect 33784 6560 34104 7584
rect 33784 6496 33792 6560
rect 33856 6496 33872 6560
rect 33936 6496 33952 6560
rect 34016 6496 34032 6560
rect 34096 6496 34104 6560
rect 33784 5472 34104 6496
rect 33784 5408 33792 5472
rect 33856 5408 33872 5472
rect 33936 5408 33952 5472
rect 34016 5408 34032 5472
rect 34096 5408 34104 5472
rect 33784 4384 34104 5408
rect 33784 4320 33792 4384
rect 33856 4320 33872 4384
rect 33936 4320 33952 4384
rect 34016 4320 34032 4384
rect 34096 4320 34104 4384
rect 33784 3296 34104 4320
rect 33784 3232 33792 3296
rect 33856 3232 33872 3296
rect 33936 3232 33952 3296
rect 34016 3232 34032 3296
rect 34096 3232 34104 3296
rect 33784 2208 34104 3232
rect 33784 2144 33792 2208
rect 33856 2144 33872 2208
rect 33936 2144 33952 2208
rect 34016 2144 34032 2208
rect 34096 2144 34104 2208
rect 33784 2128 34104 2144
rect 39258 16896 39578 17456
rect 39258 16832 39266 16896
rect 39330 16832 39346 16896
rect 39410 16832 39426 16896
rect 39490 16832 39506 16896
rect 39570 16832 39578 16896
rect 39258 15808 39578 16832
rect 39258 15744 39266 15808
rect 39330 15744 39346 15808
rect 39410 15744 39426 15808
rect 39490 15744 39506 15808
rect 39570 15744 39578 15808
rect 39258 14720 39578 15744
rect 39258 14656 39266 14720
rect 39330 14656 39346 14720
rect 39410 14656 39426 14720
rect 39490 14656 39506 14720
rect 39570 14656 39578 14720
rect 39258 13632 39578 14656
rect 39258 13568 39266 13632
rect 39330 13568 39346 13632
rect 39410 13568 39426 13632
rect 39490 13568 39506 13632
rect 39570 13568 39578 13632
rect 39258 12544 39578 13568
rect 39258 12480 39266 12544
rect 39330 12480 39346 12544
rect 39410 12480 39426 12544
rect 39490 12480 39506 12544
rect 39570 12480 39578 12544
rect 39258 11456 39578 12480
rect 39258 11392 39266 11456
rect 39330 11392 39346 11456
rect 39410 11392 39426 11456
rect 39490 11392 39506 11456
rect 39570 11392 39578 11456
rect 39258 10368 39578 11392
rect 39258 10304 39266 10368
rect 39330 10304 39346 10368
rect 39410 10304 39426 10368
rect 39490 10304 39506 10368
rect 39570 10304 39578 10368
rect 39258 9280 39578 10304
rect 39258 9216 39266 9280
rect 39330 9216 39346 9280
rect 39410 9216 39426 9280
rect 39490 9216 39506 9280
rect 39570 9216 39578 9280
rect 39258 8192 39578 9216
rect 39258 8128 39266 8192
rect 39330 8128 39346 8192
rect 39410 8128 39426 8192
rect 39490 8128 39506 8192
rect 39570 8128 39578 8192
rect 39258 7104 39578 8128
rect 39258 7040 39266 7104
rect 39330 7040 39346 7104
rect 39410 7040 39426 7104
rect 39490 7040 39506 7104
rect 39570 7040 39578 7104
rect 39258 6016 39578 7040
rect 39258 5952 39266 6016
rect 39330 5952 39346 6016
rect 39410 5952 39426 6016
rect 39490 5952 39506 6016
rect 39570 5952 39578 6016
rect 39258 4928 39578 5952
rect 39258 4864 39266 4928
rect 39330 4864 39346 4928
rect 39410 4864 39426 4928
rect 39490 4864 39506 4928
rect 39570 4864 39578 4928
rect 39258 3840 39578 4864
rect 39258 3776 39266 3840
rect 39330 3776 39346 3840
rect 39410 3776 39426 3840
rect 39490 3776 39506 3840
rect 39570 3776 39578 3840
rect 39258 2752 39578 3776
rect 39258 2688 39266 2752
rect 39330 2688 39346 2752
rect 39410 2688 39426 2752
rect 39490 2688 39506 2752
rect 39570 2688 39578 2752
rect 39258 2128 39578 2688
rect 44731 17440 45051 17456
rect 44731 17376 44739 17440
rect 44803 17376 44819 17440
rect 44883 17376 44899 17440
rect 44963 17376 44979 17440
rect 45043 17376 45051 17440
rect 44731 16352 45051 17376
rect 44731 16288 44739 16352
rect 44803 16288 44819 16352
rect 44883 16288 44899 16352
rect 44963 16288 44979 16352
rect 45043 16288 45051 16352
rect 44731 15264 45051 16288
rect 44731 15200 44739 15264
rect 44803 15200 44819 15264
rect 44883 15200 44899 15264
rect 44963 15200 44979 15264
rect 45043 15200 45051 15264
rect 44731 14176 45051 15200
rect 44731 14112 44739 14176
rect 44803 14112 44819 14176
rect 44883 14112 44899 14176
rect 44963 14112 44979 14176
rect 45043 14112 45051 14176
rect 44731 13088 45051 14112
rect 44731 13024 44739 13088
rect 44803 13024 44819 13088
rect 44883 13024 44899 13088
rect 44963 13024 44979 13088
rect 45043 13024 45051 13088
rect 44731 12000 45051 13024
rect 44731 11936 44739 12000
rect 44803 11936 44819 12000
rect 44883 11936 44899 12000
rect 44963 11936 44979 12000
rect 45043 11936 45051 12000
rect 44731 10912 45051 11936
rect 44731 10848 44739 10912
rect 44803 10848 44819 10912
rect 44883 10848 44899 10912
rect 44963 10848 44979 10912
rect 45043 10848 45051 10912
rect 44731 9824 45051 10848
rect 44731 9760 44739 9824
rect 44803 9760 44819 9824
rect 44883 9760 44899 9824
rect 44963 9760 44979 9824
rect 45043 9760 45051 9824
rect 44731 8736 45051 9760
rect 44731 8672 44739 8736
rect 44803 8672 44819 8736
rect 44883 8672 44899 8736
rect 44963 8672 44979 8736
rect 45043 8672 45051 8736
rect 44731 7648 45051 8672
rect 44731 7584 44739 7648
rect 44803 7584 44819 7648
rect 44883 7584 44899 7648
rect 44963 7584 44979 7648
rect 45043 7584 45051 7648
rect 44731 6560 45051 7584
rect 44731 6496 44739 6560
rect 44803 6496 44819 6560
rect 44883 6496 44899 6560
rect 44963 6496 44979 6560
rect 45043 6496 45051 6560
rect 44731 5472 45051 6496
rect 44731 5408 44739 5472
rect 44803 5408 44819 5472
rect 44883 5408 44899 5472
rect 44963 5408 44979 5472
rect 45043 5408 45051 5472
rect 44731 4384 45051 5408
rect 44731 4320 44739 4384
rect 44803 4320 44819 4384
rect 44883 4320 44899 4384
rect 44963 4320 44979 4384
rect 45043 4320 45051 4384
rect 44731 3296 45051 4320
rect 44731 3232 44739 3296
rect 44803 3232 44819 3296
rect 44883 3232 44899 3296
rect 44963 3232 44979 3296
rect 45043 3232 45051 3296
rect 44731 2208 45051 3232
rect 44731 2144 44739 2208
rect 44803 2144 44819 2208
rect 44883 2144 44899 2208
rect 44963 2144 44979 2208
rect 45043 2144 45051 2208
rect 44731 2128 45051 2144
use sky130_fd_sc_hd__diode_2  ANTENNA_1 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 43424 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1676037725
transform -1 0 34040 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp 1676037725
transform -1 0 31924 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 1380 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 1840 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 2484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29
timestamp 1676037725
transform 1 0 3772 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34
timestamp 1676037725
transform 1 0 4232 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41
timestamp 1676037725
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_57
timestamp 1676037725
transform 1 0 6348 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_63 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 6900 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_71
timestamp 1676037725
transform 1 0 7636 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_76
timestamp 1676037725
transform 1 0 8096 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_85
timestamp 1676037725
transform 1 0 8924 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_93
timestamp 1676037725
transform 1 0 9660 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98
timestamp 1676037725
transform 1 0 10120 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_110
timestamp 1676037725
transform 1 0 11224 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_113
timestamp 1676037725
transform 1 0 11500 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_118
timestamp 1676037725
transform 1 0 11960 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_126
timestamp 1676037725
transform 1 0 12696 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_138
timestamp 1676037725
transform 1 0 13800 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_141
timestamp 1676037725
transform 1 0 14076 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_153
timestamp 1676037725
transform 1 0 15180 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_159
timestamp 1676037725
transform 1 0 15732 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_167
timestamp 1676037725
transform 1 0 16468 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_169
timestamp 1676037725
transform 1 0 16652 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_174
timestamp 1676037725
transform 1 0 17112 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_188
timestamp 1676037725
transform 1 0 18400 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_197
timestamp 1676037725
transform 1 0 19228 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_202
timestamp 1676037725
transform 1 0 19688 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_210
timestamp 1676037725
transform 1 0 20424 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_216
timestamp 1676037725
transform 1 0 20976 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_225
timestamp 1676037725
transform 1 0 21804 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_233
timestamp 1676037725
transform 1 0 22540 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_238
timestamp 1676037725
transform 1 0 23000 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_250
timestamp 1676037725
transform 1 0 24104 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_253
timestamp 1676037725
transform 1 0 24380 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_258
timestamp 1676037725
transform 1 0 24840 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_266
timestamp 1676037725
transform 1 0 25576 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_272
timestamp 1676037725
transform 1 0 26128 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_281
timestamp 1676037725
transform 1 0 26956 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_287
timestamp 1676037725
transform 1 0 27508 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_299
timestamp 1676037725
transform 1 0 28612 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_307
timestamp 1676037725
transform 1 0 29348 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_309
timestamp 1676037725
transform 1 0 29532 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_314
timestamp 1676037725
transform 1 0 29992 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_321
timestamp 1676037725
transform 1 0 30636 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_333
timestamp 1676037725
transform 1 0 31740 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_337
timestamp 1676037725
transform 1 0 32108 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_349
timestamp 1676037725
transform 1 0 33212 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_361
timestamp 1676037725
transform 1 0 34316 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_365
timestamp 1676037725
transform 1 0 34684 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_373
timestamp 1676037725
transform 1 0 35420 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_378
timestamp 1676037725
transform 1 0 35880 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_390
timestamp 1676037725
transform 1 0 36984 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_393
timestamp 1676037725
transform 1 0 37260 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_398
timestamp 1676037725
transform 1 0 37720 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_406
timestamp 1676037725
transform 1 0 38456 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_412
timestamp 1676037725
transform 1 0 39008 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_421
timestamp 1676037725
transform 1 0 39836 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_426
timestamp 1676037725
transform 1 0 40296 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_438
timestamp 1676037725
transform 1 0 41400 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_446
timestamp 1676037725
transform 1 0 42136 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_449
timestamp 1676037725
transform 1 0 42412 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_455
timestamp 1676037725
transform 1 0 42964 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_459
timestamp 1676037725
transform 1 0 43332 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_463
timestamp 1676037725
transform 1 0 43700 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_471
timestamp 1676037725
transform 1 0 44436 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_3
timestamp 1676037725
transform 1 0 1380 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_8
timestamp 1676037725
transform 1 0 1840 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_20
timestamp 1676037725
transform 1 0 2944 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_32
timestamp 1676037725
transform 1 0 4048 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_44
timestamp 1676037725
transform 1 0 5152 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_57
timestamp 1676037725
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_69
timestamp 1676037725
transform 1 0 7452 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_73
timestamp 1676037725
transform 1 0 7820 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_85 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 8924 0 -1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_1_94
timestamp 1676037725
transform 1 0 9752 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_106
timestamp 1676037725
transform 1 0 10856 0 -1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_1_113
timestamp 1676037725
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_125
timestamp 1676037725
transform 1 0 12604 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_137
timestamp 1676037725
transform 1 0 13708 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_141
timestamp 1676037725
transform 1 0 14076 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_166
timestamp 1676037725
transform 1 0 16376 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_169
timestamp 1676037725
transform 1 0 16652 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_174
timestamp 1676037725
transform 1 0 17112 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_181
timestamp 1676037725
transform 1 0 17756 0 -1 3264
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_1_210
timestamp 1676037725
transform 1 0 20424 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_222
timestamp 1676037725
transform 1 0 21528 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_225
timestamp 1676037725
transform 1 0 21804 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_229
timestamp 1676037725
transform 1 0 22172 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_233
timestamp 1676037725
transform 1 0 22540 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_245
timestamp 1676037725
transform 1 0 23644 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_257
timestamp 1676037725
transform 1 0 24748 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_269
timestamp 1676037725
transform 1 0 25852 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_277
timestamp 1676037725
transform 1 0 26588 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_1_281
timestamp 1676037725
transform 1 0 26956 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_293
timestamp 1676037725
transform 1 0 28060 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_305
timestamp 1676037725
transform 1 0 29164 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_317
timestamp 1676037725
transform 1 0 30268 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_329
timestamp 1676037725
transform 1 0 31372 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_335
timestamp 1676037725
transform 1 0 31924 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_337
timestamp 1676037725
transform 1 0 32108 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_349
timestamp 1676037725
transform 1 0 33212 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_355
timestamp 1676037725
transform 1 0 33764 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_358
timestamp 1676037725
transform 1 0 34040 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_363
timestamp 1676037725
transform 1 0 34500 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_375
timestamp 1676037725
transform 1 0 35604 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_387
timestamp 1676037725
transform 1 0 36708 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_391
timestamp 1676037725
transform 1 0 37076 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_393
timestamp 1676037725
transform 1 0 37260 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_405
timestamp 1676037725
transform 1 0 38364 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_417
timestamp 1676037725
transform 1 0 39468 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_429
timestamp 1676037725
transform 1 0 40572 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_441
timestamp 1676037725
transform 1 0 41676 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_447
timestamp 1676037725
transform 1 0 42228 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_449
timestamp 1676037725
transform 1 0 42412 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_461
timestamp 1676037725
transform 1 0 43516 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_467
timestamp 1676037725
transform 1 0 44068 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_471
timestamp 1676037725
transform 1 0 44436 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_3
timestamp 1676037725
transform 1 0 1380 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_8
timestamp 1676037725
transform 1 0 1840 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_20
timestamp 1676037725
transform 1 0 2944 0 1 3264
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_2_29
timestamp 1676037725
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_41
timestamp 1676037725
transform 1 0 4876 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_49
timestamp 1676037725
transform 1 0 5612 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_53
timestamp 1676037725
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_65
timestamp 1676037725
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_77
timestamp 1676037725
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 1676037725
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_85
timestamp 1676037725
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_97
timestamp 1676037725
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_109
timestamp 1676037725
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_121
timestamp 1676037725
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_133
timestamp 1676037725
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_139
timestamp 1676037725
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_141
timestamp 1676037725
transform 1 0 14076 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_145
timestamp 1676037725
transform 1 0 14444 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_149
timestamp 1676037725
transform 1 0 14812 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_155
timestamp 1676037725
transform 1 0 15364 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_159
timestamp 1676037725
transform 1 0 15732 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_167
timestamp 1676037725
transform 1 0 16468 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_2_190
timestamp 1676037725
transform 1 0 18584 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_2_197
timestamp 1676037725
transform 1 0 19228 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_202
timestamp 1676037725
transform 1 0 19688 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_214
timestamp 1676037725
transform 1 0 20792 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_226
timestamp 1676037725
transform 1 0 21896 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_233
timestamp 1676037725
transform 1 0 22540 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_245
timestamp 1676037725
transform 1 0 23644 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_251
timestamp 1676037725
transform 1 0 24196 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_253
timestamp 1676037725
transform 1 0 24380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_265
timestamp 1676037725
transform 1 0 25484 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_277
timestamp 1676037725
transform 1 0 26588 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_289
timestamp 1676037725
transform 1 0 27692 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_301
timestamp 1676037725
transform 1 0 28796 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_307
timestamp 1676037725
transform 1 0 29348 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_309
timestamp 1676037725
transform 1 0 29532 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_321
timestamp 1676037725
transform 1 0 30636 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_325
timestamp 1676037725
transform 1 0 31004 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_346
timestamp 1676037725
transform 1 0 32936 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_358
timestamp 1676037725
transform 1 0 34040 0 1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_2_365
timestamp 1676037725
transform 1 0 34684 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_377
timestamp 1676037725
transform 1 0 35788 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_389
timestamp 1676037725
transform 1 0 36892 0 1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_2_398
timestamp 1676037725
transform 1 0 37720 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_410
timestamp 1676037725
transform 1 0 38824 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_418
timestamp 1676037725
transform 1 0 39560 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_421
timestamp 1676037725
transform 1 0 39836 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_433
timestamp 1676037725
transform 1 0 40940 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_445
timestamp 1676037725
transform 1 0 42044 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_457
timestamp 1676037725
transform 1 0 43148 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_2_465
timestamp 1676037725
transform 1 0 43884 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_471
timestamp 1676037725
transform 1 0 44436 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3
timestamp 1676037725
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_15
timestamp 1676037725
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_27
timestamp 1676037725
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_39
timestamp 1676037725
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_51
timestamp 1676037725
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 1676037725
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_57
timestamp 1676037725
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_69
timestamp 1676037725
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_81
timestamp 1676037725
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_93
timestamp 1676037725
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_105
timestamp 1676037725
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 1676037725
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_113
timestamp 1676037725
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_125
timestamp 1676037725
transform 1 0 12604 0 -1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_3_132
timestamp 1676037725
transform 1 0 13248 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_3_144
timestamp 1676037725
transform 1 0 14352 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_166
timestamp 1676037725
transform 1 0 16376 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_169
timestamp 1676037725
transform 1 0 16652 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_174
timestamp 1676037725
transform 1 0 17112 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_181
timestamp 1676037725
transform 1 0 17756 0 -1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_3_205
timestamp 1676037725
transform 1 0 19964 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_217
timestamp 1676037725
transform 1 0 21068 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_223
timestamp 1676037725
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_225
timestamp 1676037725
transform 1 0 21804 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_230
timestamp 1676037725
transform 1 0 22264 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_234
timestamp 1676037725
transform 1 0 22632 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_238
timestamp 1676037725
transform 1 0 23000 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_250
timestamp 1676037725
transform 1 0 24104 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_262
timestamp 1676037725
transform 1 0 25208 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_274
timestamp 1676037725
transform 1 0 26312 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_3_281
timestamp 1676037725
transform 1 0 26956 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_285
timestamp 1676037725
transform 1 0 27324 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_295
timestamp 1676037725
transform 1 0 28244 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_307
timestamp 1676037725
transform 1 0 29348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_319
timestamp 1676037725
transform 1 0 30452 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_3_334
timestamp 1676037725
transform 1 0 31832 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_337
timestamp 1676037725
transform 1 0 32108 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_3_345
timestamp 1676037725
transform 1 0 32844 0 -1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_3_354
timestamp 1676037725
transform 1 0 33672 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_3_366
timestamp 1676037725
transform 1 0 34776 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_3_372
timestamp 1676037725
transform 1 0 35328 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_380
timestamp 1676037725
transform 1 0 36064 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_388
timestamp 1676037725
transform 1 0 36800 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_393
timestamp 1676037725
transform 1 0 37260 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_415
timestamp 1676037725
transform 1 0 39284 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_427
timestamp 1676037725
transform 1 0 40388 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_439
timestamp 1676037725
transform 1 0 41492 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_447
timestamp 1676037725
transform 1 0 42228 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_449
timestamp 1676037725
transform 1 0 42412 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_461
timestamp 1676037725
transform 1 0 43516 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3
timestamp 1676037725
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_15
timestamp 1676037725
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1676037725
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_29
timestamp 1676037725
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_46
timestamp 1676037725
transform 1 0 5336 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_58
timestamp 1676037725
transform 1 0 6440 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_70
timestamp 1676037725
transform 1 0 7544 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_4_82
timestamp 1676037725
transform 1 0 8648 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_85
timestamp 1676037725
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_97
timestamp 1676037725
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_109
timestamp 1676037725
transform 1 0 11132 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_115
timestamp 1676037725
transform 1 0 11684 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_132
timestamp 1676037725
transform 1 0 13248 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_4_141
timestamp 1676037725
transform 1 0 14076 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_149
timestamp 1676037725
transform 1 0 14812 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_154
timestamp 1676037725
transform 1 0 15272 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_178
timestamp 1676037725
transform 1 0 17480 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_186
timestamp 1676037725
transform 1 0 18216 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_4_190
timestamp 1676037725
transform 1 0 18584 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_4_197
timestamp 1676037725
transform 1 0 19228 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_4_202
timestamp 1676037725
transform 1 0 19688 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_210
timestamp 1676037725
transform 1 0 20424 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_231
timestamp 1676037725
transform 1 0 22356 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_241
timestamp 1676037725
transform 1 0 23276 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_4_249
timestamp 1676037725
transform 1 0 24012 0 1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_253
timestamp 1676037725
transform 1 0 24380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_265
timestamp 1676037725
transform 1 0 25484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_277
timestamp 1676037725
transform 1 0 26588 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_4_299
timestamp 1676037725
transform 1 0 28612 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_307
timestamp 1676037725
transform 1 0 29348 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_309
timestamp 1676037725
transform 1 0 29532 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_321
timestamp 1676037725
transform 1 0 30636 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_4_347
timestamp 1676037725
transform 1 0 33028 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_4_357
timestamp 1676037725
transform 1 0 33948 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_363
timestamp 1676037725
transform 1 0 34500 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_365
timestamp 1676037725
transform 1 0 34684 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_4_393
timestamp 1676037725
transform 1 0 37260 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_400
timestamp 1676037725
transform 1 0 37904 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_404
timestamp 1676037725
transform 1 0 38272 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_408
timestamp 1676037725
transform 1 0 38640 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_421
timestamp 1676037725
transform 1 0 39836 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_433
timestamp 1676037725
transform 1 0 40940 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_445
timestamp 1676037725
transform 1 0 42044 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_457
timestamp 1676037725
transform 1 0 43148 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_465
timestamp 1676037725
transform 1 0 43884 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_471
timestamp 1676037725
transform 1 0 44436 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_3
timestamp 1676037725
transform 1 0 1380 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_15
timestamp 1676037725
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_27
timestamp 1676037725
transform 1 0 3588 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_47
timestamp 1676037725
transform 1 0 5428 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1676037725
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_57
timestamp 1676037725
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_69
timestamp 1676037725
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_81
timestamp 1676037725
transform 1 0 8556 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_87
timestamp 1676037725
transform 1 0 9108 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_93
timestamp 1676037725
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_105
timestamp 1676037725
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1676037725
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_113
timestamp 1676037725
transform 1 0 11500 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_5_137
timestamp 1676037725
transform 1 0 13708 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_145
timestamp 1676037725
transform 1 0 14444 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_153
timestamp 1676037725
transform 1 0 15180 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_159
timestamp 1676037725
transform 1 0 15732 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 1676037725
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_169
timestamp 1676037725
transform 1 0 16652 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_191
timestamp 1676037725
transform 1 0 18676 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_5_198
timestamp 1676037725
transform 1 0 19320 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_210
timestamp 1676037725
transform 1 0 20424 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_5_219
timestamp 1676037725
transform 1 0 21252 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_223
timestamp 1676037725
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_225
timestamp 1676037725
transform 1 0 21804 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_5_237
timestamp 1676037725
transform 1 0 22908 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_255
timestamp 1676037725
transform 1 0 24564 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_267
timestamp 1676037725
transform 1 0 25668 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_5_279
timestamp 1676037725
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_281
timestamp 1676037725
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_293
timestamp 1676037725
transform 1 0 28060 0 -1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_5_319
timestamp 1676037725
transform 1 0 30452 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_331
timestamp 1676037725
transform 1 0 31556 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_335
timestamp 1676037725
transform 1 0 31924 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_5_337
timestamp 1676037725
transform 1 0 32108 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_5_347
timestamp 1676037725
transform 1 0 33028 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_5_375
timestamp 1676037725
transform 1 0 35604 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_384
timestamp 1676037725
transform 1 0 36432 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_5_393
timestamp 1676037725
transform 1 0 37260 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_5_402
timestamp 1676037725
transform 1 0 38088 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_411
timestamp 1676037725
transform 1 0 38916 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_419
timestamp 1676037725
transform 1 0 39652 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_425
timestamp 1676037725
transform 1 0 40204 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_430
timestamp 1676037725
transform 1 0 40664 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_437
timestamp 1676037725
transform 1 0 41308 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_5_445
timestamp 1676037725
transform 1 0 42044 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_449
timestamp 1676037725
transform 1 0 42412 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_5_456
timestamp 1676037725
transform 1 0 43056 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_468
timestamp 1676037725
transform 1 0 44160 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_472
timestamp 1676037725
transform 1 0 44528 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3
timestamp 1676037725
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_15
timestamp 1676037725
transform 1 0 2484 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_19
timestamp 1676037725
transform 1 0 2852 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_26
timestamp 1676037725
transform 1 0 3496 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_29
timestamp 1676037725
transform 1 0 3772 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_47
timestamp 1676037725
transform 1 0 5428 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_6_56
timestamp 1676037725
transform 1 0 6256 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_68
timestamp 1676037725
transform 1 0 7360 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_80
timestamp 1676037725
transform 1 0 8464 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_6_85
timestamp 1676037725
transform 1 0 8924 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_91
timestamp 1676037725
transform 1 0 9476 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_97
timestamp 1676037725
transform 1 0 10028 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_6_121
timestamp 1676037725
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_133
timestamp 1676037725
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1676037725
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_141
timestamp 1676037725
transform 1 0 14076 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_147
timestamp 1676037725
transform 1 0 14628 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_159
timestamp 1676037725
transform 1 0 15732 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_163
timestamp 1676037725
transform 1 0 16100 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_187
timestamp 1676037725
transform 1 0 18308 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_194
timestamp 1676037725
transform 1 0 18952 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_6_197
timestamp 1676037725
transform 1 0 19228 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_205
timestamp 1676037725
transform 1 0 19964 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_215
timestamp 1676037725
transform 1 0 20884 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_6_235
timestamp 1676037725
transform 1 0 22724 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_247
timestamp 1676037725
transform 1 0 23828 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_251
timestamp 1676037725
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_253
timestamp 1676037725
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_265
timestamp 1676037725
transform 1 0 25484 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_271
timestamp 1676037725
transform 1 0 26036 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_275
timestamp 1676037725
transform 1 0 26404 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_295
timestamp 1676037725
transform 1 0 28244 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_6_302
timestamp 1676037725
transform 1 0 28888 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_6_309
timestamp 1676037725
transform 1 0 29532 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_6_320
timestamp 1676037725
transform 1 0 30544 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_328
timestamp 1676037725
transform 1 0 31280 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_332
timestamp 1676037725
transform 1 0 31648 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_339
timestamp 1676037725
transform 1 0 32292 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_351
timestamp 1676037725
transform 1 0 33396 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_6_361
timestamp 1676037725
transform 1 0 34316 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_365
timestamp 1676037725
transform 1 0 34684 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_370
timestamp 1676037725
transform 1 0 35144 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_6_377
timestamp 1676037725
transform 1 0 35788 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_6_390
timestamp 1676037725
transform 1 0 36984 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_418
timestamp 1676037725
transform 1 0 39560 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_421
timestamp 1676037725
transform 1 0 39836 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_427
timestamp 1676037725
transform 1 0 40388 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_431
timestamp 1676037725
transform 1 0 40756 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_452
timestamp 1676037725
transform 1 0 42688 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_6_464
timestamp 1676037725
transform 1 0 43792 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_471
timestamp 1676037725
transform 1 0 44436 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_3
timestamp 1676037725
transform 1 0 1380 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_8
timestamp 1676037725
transform 1 0 1840 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_20
timestamp 1676037725
transform 1 0 2944 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_7_40
timestamp 1676037725
transform 1 0 4784 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_52
timestamp 1676037725
transform 1 0 5888 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_7_57
timestamp 1676037725
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_69
timestamp 1676037725
transform 1 0 7452 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_73
timestamp 1676037725
transform 1 0 7820 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_90
timestamp 1676037725
transform 1 0 9384 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_110
timestamp 1676037725
transform 1 0 11224 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_7_113
timestamp 1676037725
transform 1 0 11500 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_119
timestamp 1676037725
transform 1 0 12052 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_125
timestamp 1676037725
transform 1 0 12604 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_136
timestamp 1676037725
transform 1 0 13616 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_145
timestamp 1676037725
transform 1 0 14444 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_7_154
timestamp 1676037725
transform 1 0 15272 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_166
timestamp 1676037725
transform 1 0 16376 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_7_169
timestamp 1676037725
transform 1 0 16652 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_175
timestamp 1676037725
transform 1 0 17204 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_185
timestamp 1676037725
transform 1 0 18124 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_198
timestamp 1676037725
transform 1 0 19320 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_209
timestamp 1676037725
transform 1 0 20332 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_220
timestamp 1676037725
transform 1 0 21344 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_225
timestamp 1676037725
transform 1 0 21804 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_7_243
timestamp 1676037725
transform 1 0 23460 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_7_254
timestamp 1676037725
transform 1 0 24472 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_7_267
timestamp 1676037725
transform 1 0 25668 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_279
timestamp 1676037725
transform 1 0 26772 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_7_281
timestamp 1676037725
transform 1 0 26956 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_7_293
timestamp 1676037725
transform 1 0 28060 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_297
timestamp 1676037725
transform 1 0 28428 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_314
timestamp 1676037725
transform 1 0 29992 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_7_326
timestamp 1676037725
transform 1 0 31096 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_334
timestamp 1676037725
transform 1 0 31832 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_7_337
timestamp 1676037725
transform 1 0 32108 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_343
timestamp 1676037725
transform 1 0 32660 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_352
timestamp 1676037725
transform 1 0 33488 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_363
timestamp 1676037725
transform 1 0 34500 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_373
timestamp 1676037725
transform 1 0 35420 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_377
timestamp 1676037725
transform 1 0 35788 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_381
timestamp 1676037725
transform 1 0 36156 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_7_389
timestamp 1676037725
transform 1 0 36892 0 -1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_7_393
timestamp 1676037725
transform 1 0 37260 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_405
timestamp 1676037725
transform 1 0 38364 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_409
timestamp 1676037725
transform 1 0 38732 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_7_420
timestamp 1676037725
transform 1 0 39744 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_7_446
timestamp 1676037725
transform 1 0 42136 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_449
timestamp 1676037725
transform 1 0 42412 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_454
timestamp 1676037725
transform 1 0 42872 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_466
timestamp 1676037725
transform 1 0 43976 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_472
timestamp 1676037725
transform 1 0 44528 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_3
timestamp 1676037725
transform 1 0 1380 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_8_20
timestamp 1676037725
transform 1 0 2944 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_29
timestamp 1676037725
transform 1 0 3772 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_47
timestamp 1676037725
transform 1 0 5428 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_59
timestamp 1676037725
transform 1 0 6532 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_65
timestamp 1676037725
transform 1 0 7084 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_82
timestamp 1676037725
transform 1 0 8648 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_85
timestamp 1676037725
transform 1 0 8924 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_96
timestamp 1676037725
transform 1 0 9936 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_108
timestamp 1676037725
transform 1 0 11040 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_114
timestamp 1676037725
transform 1 0 11592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_118
timestamp 1676037725
transform 1 0 11960 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_138
timestamp 1676037725
transform 1 0 13800 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_141
timestamp 1676037725
transform 1 0 14076 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_150
timestamp 1676037725
transform 1 0 14904 0 1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_8_157
timestamp 1676037725
transform 1 0 15548 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_169
timestamp 1676037725
transform 1 0 16652 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_181
timestamp 1676037725
transform 1 0 17756 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_194
timestamp 1676037725
transform 1 0 18952 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_197
timestamp 1676037725
transform 1 0 19228 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_8_207
timestamp 1676037725
transform 1 0 20148 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_213
timestamp 1676037725
transform 1 0 20700 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_217
timestamp 1676037725
transform 1 0 21068 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_229
timestamp 1676037725
transform 1 0 22172 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_233
timestamp 1676037725
transform 1 0 22540 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_237
timestamp 1676037725
transform 1 0 22908 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_245
timestamp 1676037725
transform 1 0 23644 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_250
timestamp 1676037725
transform 1 0 24104 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_253
timestamp 1676037725
transform 1 0 24380 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_275
timestamp 1676037725
transform 1 0 26404 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_287
timestamp 1676037725
transform 1 0 27508 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_291
timestamp 1676037725
transform 1 0 27876 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_295
timestamp 1676037725
transform 1 0 28244 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_8_302
timestamp 1676037725
transform 1 0 28888 0 1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_8_309
timestamp 1676037725
transform 1 0 29532 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_321
timestamp 1676037725
transform 1 0 30636 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_8_330
timestamp 1676037725
transform 1 0 31464 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_338
timestamp 1676037725
transform 1 0 32200 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_349
timestamp 1676037725
transform 1 0 33212 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_360
timestamp 1676037725
transform 1 0 34224 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_8_365
timestamp 1676037725
transform 1 0 34684 0 1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_8_379
timestamp 1676037725
transform 1 0 35972 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_391
timestamp 1676037725
transform 1 0 37076 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_403
timestamp 1676037725
transform 1 0 38180 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_407
timestamp 1676037725
transform 1 0 38548 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_416
timestamp 1676037725
transform 1 0 39376 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_421
timestamp 1676037725
transform 1 0 39836 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_428
timestamp 1676037725
transform 1 0 40480 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_436
timestamp 1676037725
transform 1 0 41216 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_443
timestamp 1676037725
transform 1 0 41860 0 1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_8_450
timestamp 1676037725
transform 1 0 42504 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_462
timestamp 1676037725
transform 1 0 43608 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_8_470
timestamp 1676037725
transform 1 0 44344 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_3
timestamp 1676037725
transform 1 0 1380 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_9_8
timestamp 1676037725
transform 1 0 1840 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_9_36
timestamp 1676037725
transform 1 0 4416 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_53
timestamp 1676037725
transform 1 0 5980 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_57
timestamp 1676037725
transform 1 0 6348 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_9_64
timestamp 1676037725
transform 1 0 6992 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_72
timestamp 1676037725
transform 1 0 7728 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_93
timestamp 1676037725
transform 1 0 9660 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_106
timestamp 1676037725
transform 1 0 10856 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_9_113
timestamp 1676037725
transform 1 0 11500 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_121
timestamp 1676037725
transform 1 0 12236 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_126
timestamp 1676037725
transform 1 0 12696 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_146
timestamp 1676037725
transform 1 0 14536 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_9_153
timestamp 1676037725
transform 1 0 15180 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_165
timestamp 1676037725
transform 1 0 16284 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_169
timestamp 1676037725
transform 1 0 16652 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_180
timestamp 1676037725
transform 1 0 17664 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_184
timestamp 1676037725
transform 1 0 18032 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_9_194
timestamp 1676037725
transform 1 0 18952 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_200
timestamp 1676037725
transform 1 0 19504 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_209
timestamp 1676037725
transform 1 0 20332 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_220
timestamp 1676037725
transform 1 0 21344 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_225
timestamp 1676037725
transform 1 0 21804 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_232
timestamp 1676037725
transform 1 0 22448 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_239
timestamp 1676037725
transform 1 0 23092 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_245
timestamp 1676037725
transform 1 0 23644 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_252
timestamp 1676037725
transform 1 0 24288 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_262
timestamp 1676037725
transform 1 0 25208 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_269
timestamp 1676037725
transform 1 0 25852 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_277
timestamp 1676037725
transform 1 0 26588 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_281
timestamp 1676037725
transform 1 0 26956 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_293
timestamp 1676037725
transform 1 0 28060 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_297
timestamp 1676037725
transform 1 0 28428 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_314
timestamp 1676037725
transform 1 0 29992 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_327
timestamp 1676037725
transform 1 0 31188 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_335
timestamp 1676037725
transform 1 0 31924 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_337
timestamp 1676037725
transform 1 0 32108 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_355
timestamp 1676037725
transform 1 0 33764 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_366
timestamp 1676037725
transform 1 0 34776 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_9_383
timestamp 1676037725
transform 1 0 36340 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_391
timestamp 1676037725
transform 1 0 37076 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_393
timestamp 1676037725
transform 1 0 37260 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_9_398
timestamp 1676037725
transform 1 0 37720 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_406
timestamp 1676037725
transform 1 0 38456 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_413
timestamp 1676037725
transform 1 0 39100 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_423
timestamp 1676037725
transform 1 0 40020 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_432
timestamp 1676037725
transform 1 0 40848 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_439
timestamp 1676037725
transform 1 0 41492 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_447
timestamp 1676037725
transform 1 0 42228 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_449
timestamp 1676037725
transform 1 0 42412 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_454
timestamp 1676037725
transform 1 0 42872 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_466
timestamp 1676037725
transform 1 0 43976 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_471
timestamp 1676037725
transform 1 0 44436 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_10_3
timestamp 1676037725
transform 1 0 1380 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_9
timestamp 1676037725
transform 1 0 1932 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_26
timestamp 1676037725
transform 1 0 3496 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_29
timestamp 1676037725
transform 1 0 3772 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_47
timestamp 1676037725
transform 1 0 5428 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_59
timestamp 1676037725
transform 1 0 6532 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_71
timestamp 1676037725
transform 1 0 7636 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_80
timestamp 1676037725
transform 1 0 8464 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_85
timestamp 1676037725
transform 1 0 8924 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_103
timestamp 1676037725
transform 1 0 10580 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_115
timestamp 1676037725
transform 1 0 11684 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_10_124
timestamp 1676037725
transform 1 0 12512 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_130
timestamp 1676037725
transform 1 0 13064 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_136
timestamp 1676037725
transform 1 0 13616 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_141
timestamp 1676037725
transform 1 0 14076 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_145
timestamp 1676037725
transform 1 0 14444 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_149
timestamp 1676037725
transform 1 0 14812 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_156
timestamp 1676037725
transform 1 0 15456 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_163
timestamp 1676037725
transform 1 0 16100 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_170
timestamp 1676037725
transform 1 0 16744 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_194
timestamp 1676037725
transform 1 0 18952 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_197
timestamp 1676037725
transform 1 0 19228 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_201
timestamp 1676037725
transform 1 0 19596 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_211
timestamp 1676037725
transform 1 0 20516 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_218
timestamp 1676037725
transform 1 0 21160 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_238
timestamp 1676037725
transform 1 0 23000 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_10_245
timestamp 1676037725
transform 1 0 23644 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_251
timestamp 1676037725
transform 1 0 24196 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_253
timestamp 1676037725
transform 1 0 24380 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_262
timestamp 1676037725
transform 1 0 25208 0 1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_10_269
timestamp 1676037725
transform 1 0 25852 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_281
timestamp 1676037725
transform 1 0 26956 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_293
timestamp 1676037725
transform 1 0 28060 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_299
timestamp 1676037725
transform 1 0 28612 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_10_305
timestamp 1676037725
transform 1 0 29164 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_309
timestamp 1676037725
transform 1 0 29532 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_314
timestamp 1676037725
transform 1 0 29992 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_332
timestamp 1676037725
transform 1 0 31648 0 1 7616
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_10_343
timestamp 1676037725
transform 1 0 32660 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_355
timestamp 1676037725
transform 1 0 33764 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_363
timestamp 1676037725
transform 1 0 34500 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_365
timestamp 1676037725
transform 1 0 34684 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_376
timestamp 1676037725
transform 1 0 35696 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_388
timestamp 1676037725
transform 1 0 36800 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_10_400
timestamp 1676037725
transform 1 0 37904 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_409
timestamp 1676037725
transform 1 0 38732 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_413
timestamp 1676037725
transform 1 0 39100 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_418
timestamp 1676037725
transform 1 0 39560 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_421
timestamp 1676037725
transform 1 0 39836 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_443
timestamp 1676037725
transform 1 0 41860 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_10_467
timestamp 1676037725
transform 1 0 44068 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_11_3
timestamp 1676037725
transform 1 0 1380 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_11_27
timestamp 1676037725
transform 1 0 3588 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_47
timestamp 1676037725
transform 1 0 5428 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 1676037725
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_11_57
timestamp 1676037725
transform 1 0 6348 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_11_66
timestamp 1676037725
transform 1 0 7176 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_78
timestamp 1676037725
transform 1 0 8280 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_11_98
timestamp 1676037725
transform 1 0 10120 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_110
timestamp 1676037725
transform 1 0 11224 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_113
timestamp 1676037725
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_125
timestamp 1676037725
transform 1 0 12604 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_137
timestamp 1676037725
transform 1 0 13708 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_141
timestamp 1676037725
transform 1 0 14076 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_145
timestamp 1676037725
transform 1 0 14444 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_157
timestamp 1676037725
transform 1 0 15548 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_11_166
timestamp 1676037725
transform 1 0 16376 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_169
timestamp 1676037725
transform 1 0 16652 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_191
timestamp 1676037725
transform 1 0 18676 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_198
timestamp 1676037725
transform 1 0 19320 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_209
timestamp 1676037725
transform 1 0 20332 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_216
timestamp 1676037725
transform 1 0 20976 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_225
timestamp 1676037725
transform 1 0 21804 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_11_232
timestamp 1676037725
transform 1 0 22448 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_238
timestamp 1676037725
transform 1 0 23000 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_11_259
timestamp 1676037725
transform 1 0 24932 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_265
timestamp 1676037725
transform 1 0 25484 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_275
timestamp 1676037725
transform 1 0 26404 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_279
timestamp 1676037725
transform 1 0 26772 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_281
timestamp 1676037725
transform 1 0 26956 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_289
timestamp 1676037725
transform 1 0 27692 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_306
timestamp 1676037725
transform 1 0 29256 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_326
timestamp 1676037725
transform 1 0 31096 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_11_333
timestamp 1676037725
transform 1 0 31740 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_11_337
timestamp 1676037725
transform 1 0 32108 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_349
timestamp 1676037725
transform 1 0 33212 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_11_360
timestamp 1676037725
transform 1 0 34224 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_11_380
timestamp 1676037725
transform 1 0 36064 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_393
timestamp 1676037725
transform 1 0 37260 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_404
timestamp 1676037725
transform 1 0 38272 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_416
timestamp 1676037725
transform 1 0 39376 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_431
timestamp 1676037725
transform 1 0 40756 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_443
timestamp 1676037725
transform 1 0 41860 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_447
timestamp 1676037725
transform 1 0 42228 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_449
timestamp 1676037725
transform 1 0 42412 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_461
timestamp 1676037725
transform 1 0 43516 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_3
timestamp 1676037725
transform 1 0 1380 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_9
timestamp 1676037725
transform 1 0 1932 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_13
timestamp 1676037725
transform 1 0 2300 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_26
timestamp 1676037725
transform 1 0 3496 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_29
timestamp 1676037725
transform 1 0 3772 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_39
timestamp 1676037725
transform 1 0 4692 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_47
timestamp 1676037725
transform 1 0 5428 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_69
timestamp 1676037725
transform 1 0 7452 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_82
timestamp 1676037725
transform 1 0 8648 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_85
timestamp 1676037725
transform 1 0 8924 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_90
timestamp 1676037725
transform 1 0 9384 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_110
timestamp 1676037725
transform 1 0 11224 0 1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_12_117
timestamp 1676037725
transform 1 0 11868 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_129
timestamp 1676037725
transform 1 0 12972 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_12_137
timestamp 1676037725
transform 1 0 13708 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_141
timestamp 1676037725
transform 1 0 14076 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_152
timestamp 1676037725
transform 1 0 15088 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_167
timestamp 1676037725
transform 1 0 16468 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_12_194
timestamp 1676037725
transform 1 0 18952 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_197
timestamp 1676037725
transform 1 0 19228 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_208
timestamp 1676037725
transform 1 0 20240 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_220
timestamp 1676037725
transform 1 0 21344 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_230
timestamp 1676037725
transform 1 0 22264 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_250
timestamp 1676037725
transform 1 0 24104 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_253
timestamp 1676037725
transform 1 0 24380 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_277
timestamp 1676037725
transform 1 0 26588 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_283
timestamp 1676037725
transform 1 0 27140 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_293
timestamp 1676037725
transform 1 0 28060 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_301
timestamp 1676037725
transform 1 0 28796 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_306
timestamp 1676037725
transform 1 0 29256 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_309
timestamp 1676037725
transform 1 0 29532 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_12_321
timestamp 1676037725
transform 1 0 30636 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_342
timestamp 1676037725
transform 1 0 32568 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_12_349
timestamp 1676037725
transform 1 0 33212 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_357
timestamp 1676037725
transform 1 0 33948 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_362
timestamp 1676037725
transform 1 0 34408 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_365
timestamp 1676037725
transform 1 0 34684 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_12_384
timestamp 1676037725
transform 1 0 36432 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_12_392
timestamp 1676037725
transform 1 0 37168 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_12_411
timestamp 1676037725
transform 1 0 38916 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_419
timestamp 1676037725
transform 1 0 39652 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_421
timestamp 1676037725
transform 1 0 39836 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_433
timestamp 1676037725
transform 1 0 40940 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_445
timestamp 1676037725
transform 1 0 42044 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_457
timestamp 1676037725
transform 1 0 43148 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_12_465
timestamp 1676037725
transform 1 0 43884 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_471
timestamp 1676037725
transform 1 0 44436 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_13_3
timestamp 1676037725
transform 1 0 1380 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_9
timestamp 1676037725
transform 1 0 1932 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_13
timestamp 1676037725
transform 1 0 2300 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_20
timestamp 1676037725
transform 1 0 2944 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_40
timestamp 1676037725
transform 1 0 4784 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_13_53
timestamp 1676037725
transform 1 0 5980 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_13_57
timestamp 1676037725
transform 1 0 6348 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_65
timestamp 1676037725
transform 1 0 7084 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_82
timestamp 1676037725
transform 1 0 8648 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_13_90
timestamp 1676037725
transform 1 0 9384 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_13_109
timestamp 1676037725
transform 1 0 11132 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_113
timestamp 1676037725
transform 1 0 11500 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_13_118
timestamp 1676037725
transform 1 0 11960 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_126
timestamp 1676037725
transform 1 0 12696 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_13_144
timestamp 1676037725
transform 1 0 14352 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_13_166
timestamp 1676037725
transform 1 0 16376 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_169
timestamp 1676037725
transform 1 0 16652 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_175
timestamp 1676037725
transform 1 0 17204 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_182
timestamp 1676037725
transform 1 0 17848 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_13_207
timestamp 1676037725
transform 1 0 20148 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_219
timestamp 1676037725
transform 1 0 21252 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_223
timestamp 1676037725
transform 1 0 21620 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_225
timestamp 1676037725
transform 1 0 21804 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_13_256
timestamp 1676037725
transform 1 0 24656 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_13_265
timestamp 1676037725
transform 1 0 25484 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_276
timestamp 1676037725
transform 1 0 26496 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_13_281
timestamp 1676037725
transform 1 0 26956 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_293
timestamp 1676037725
transform 1 0 28060 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_317
timestamp 1676037725
transform 1 0 30268 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_327
timestamp 1676037725
transform 1 0 31188 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_334
timestamp 1676037725
transform 1 0 31832 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_337
timestamp 1676037725
transform 1 0 32108 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_342
timestamp 1676037725
transform 1 0 32568 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_369
timestamp 1676037725
transform 1 0 35052 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_382
timestamp 1676037725
transform 1 0 36248 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_386
timestamp 1676037725
transform 1 0 36616 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_390
timestamp 1676037725
transform 1 0 36984 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_393
timestamp 1676037725
transform 1 0 37260 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_399
timestamp 1676037725
transform 1 0 37812 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_411
timestamp 1676037725
transform 1 0 38916 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_423
timestamp 1676037725
transform 1 0 40020 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_435
timestamp 1676037725
transform 1 0 41124 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_13_447
timestamp 1676037725
transform 1 0 42228 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_449
timestamp 1676037725
transform 1 0 42412 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_461
timestamp 1676037725
transform 1 0 43516 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_3
timestamp 1676037725
transform 1 0 1380 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_14_9
timestamp 1676037725
transform 1 0 1932 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_26
timestamp 1676037725
transform 1 0 3496 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_14_29
timestamp 1676037725
transform 1 0 3772 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_14_53
timestamp 1676037725
transform 1 0 5980 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_14_75
timestamp 1676037725
transform 1 0 8004 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_82
timestamp 1676037725
transform 1 0 8648 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_85
timestamp 1676037725
transform 1 0 8924 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_96
timestamp 1676037725
transform 1 0 9936 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_100
timestamp 1676037725
transform 1 0 10304 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_121
timestamp 1676037725
transform 1 0 12236 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_138
timestamp 1676037725
transform 1 0 13800 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_141
timestamp 1676037725
transform 1 0 14076 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_145
timestamp 1676037725
transform 1 0 14444 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_14_151
timestamp 1676037725
transform 1 0 14996 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_157
timestamp 1676037725
transform 1 0 15548 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_14_178
timestamp 1676037725
transform 1 0 17480 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_14_193
timestamp 1676037725
transform 1 0 18860 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_197
timestamp 1676037725
transform 1 0 19228 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_202
timestamp 1676037725
transform 1 0 19688 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_214
timestamp 1676037725
transform 1 0 20792 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_238
timestamp 1676037725
transform 1 0 23000 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_14_247
timestamp 1676037725
transform 1 0 23828 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_251
timestamp 1676037725
transform 1 0 24196 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_253
timestamp 1676037725
transform 1 0 24380 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_14_258
timestamp 1676037725
transform 1 0 24840 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_266
timestamp 1676037725
transform 1 0 25576 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_283
timestamp 1676037725
transform 1 0 27140 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_295
timestamp 1676037725
transform 1 0 28244 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_307
timestamp 1676037725
transform 1 0 29348 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_309
timestamp 1676037725
transform 1 0 29532 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_327
timestamp 1676037725
transform 1 0 31188 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_338
timestamp 1676037725
transform 1 0 32200 0 1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_14_347
timestamp 1676037725
transform 1 0 33028 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_359
timestamp 1676037725
transform 1 0 34132 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_363
timestamp 1676037725
transform 1 0 34500 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_365
timestamp 1676037725
transform 1 0 34684 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_377
timestamp 1676037725
transform 1 0 35788 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_14_385
timestamp 1676037725
transform 1 0 36524 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_14_404
timestamp 1676037725
transform 1 0 38272 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_411
timestamp 1676037725
transform 1 0 38916 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_419
timestamp 1676037725
transform 1 0 39652 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_421
timestamp 1676037725
transform 1 0 39836 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_433
timestamp 1676037725
transform 1 0 40940 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_445
timestamp 1676037725
transform 1 0 42044 0 1 9792
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_14_456
timestamp 1676037725
transform 1 0 43056 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_468
timestamp 1676037725
transform 1 0 44160 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_472
timestamp 1676037725
transform 1 0 44528 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_3
timestamp 1676037725
transform 1 0 1380 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_15_15
timestamp 1676037725
transform 1 0 2484 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_27
timestamp 1676037725
transform 1 0 3588 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_15_47
timestamp 1676037725
transform 1 0 5428 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_55
timestamp 1676037725
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_15_57
timestamp 1676037725
transform 1 0 6348 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_15_79
timestamp 1676037725
transform 1 0 8372 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_15_96
timestamp 1676037725
transform 1 0 9936 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_15_109
timestamp 1676037725
transform 1 0 11132 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_113
timestamp 1676037725
transform 1 0 11500 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_131
timestamp 1676037725
transform 1 0 13156 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_144
timestamp 1676037725
transform 1 0 14352 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_148
timestamp 1676037725
transform 1 0 14720 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_152
timestamp 1676037725
transform 1 0 15088 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_159
timestamp 1676037725
transform 1 0 15732 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_166
timestamp 1676037725
transform 1 0 16376 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_169
timestamp 1676037725
transform 1 0 16652 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_15_181
timestamp 1676037725
transform 1 0 17756 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_189
timestamp 1676037725
transform 1 0 18492 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_15_194
timestamp 1676037725
transform 1 0 18952 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_15_202
timestamp 1676037725
transform 1 0 19688 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_209
timestamp 1676037725
transform 1 0 20332 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_15_216
timestamp 1676037725
transform 1 0 20976 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_15_225
timestamp 1676037725
transform 1 0 21804 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_231
timestamp 1676037725
transform 1 0 22356 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_235
timestamp 1676037725
transform 1 0 22724 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_259
timestamp 1676037725
transform 1 0 24932 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_263
timestamp 1676037725
transform 1 0 25300 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_267
timestamp 1676037725
transform 1 0 25668 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_15_274
timestamp 1676037725
transform 1 0 26312 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_15_281
timestamp 1676037725
transform 1 0 26956 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_15_289
timestamp 1676037725
transform 1 0 27692 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_297
timestamp 1676037725
transform 1 0 28428 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_319
timestamp 1676037725
transform 1 0 30452 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_15_329
timestamp 1676037725
transform 1 0 31372 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_335
timestamp 1676037725
transform 1 0 31924 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_337
timestamp 1676037725
transform 1 0 32108 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_15_342
timestamp 1676037725
transform 1 0 32568 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_15_354
timestamp 1676037725
transform 1 0 33672 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_375
timestamp 1676037725
transform 1 0 35604 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_15_386
timestamp 1676037725
transform 1 0 36616 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_15_393
timestamp 1676037725
transform 1 0 37260 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_411
timestamp 1676037725
transform 1 0 38916 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_421
timestamp 1676037725
transform 1 0 39836 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_433
timestamp 1676037725
transform 1 0 40940 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_15_445
timestamp 1676037725
transform 1 0 42044 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_449
timestamp 1676037725
transform 1 0 42412 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_15_458
timestamp 1676037725
transform 1 0 43240 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_15_470
timestamp 1676037725
transform 1 0 44344 0 -1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_16_3
timestamp 1676037725
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_15
timestamp 1676037725
transform 1 0 2484 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_16_26
timestamp 1676037725
transform 1 0 3496 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_29
timestamp 1676037725
transform 1 0 3772 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_49
timestamp 1676037725
transform 1 0 5612 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_56
timestamp 1676037725
transform 1 0 6256 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_60
timestamp 1676037725
transform 1 0 6624 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_70
timestamp 1676037725
transform 1 0 7544 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_82
timestamp 1676037725
transform 1 0 8648 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_16_85
timestamp 1676037725
transform 1 0 8924 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_16_93
timestamp 1676037725
transform 1 0 9660 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_16_112
timestamp 1676037725
transform 1 0 11408 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_120
timestamp 1676037725
transform 1 0 12144 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_138
timestamp 1676037725
transform 1 0 13800 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_141
timestamp 1676037725
transform 1 0 14076 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_16_148
timestamp 1676037725
transform 1 0 14720 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_16_156
timestamp 1676037725
transform 1 0 15456 0 1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_16_175
timestamp 1676037725
transform 1 0 17204 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_187
timestamp 1676037725
transform 1 0 18308 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_195
timestamp 1676037725
transform 1 0 19044 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_197
timestamp 1676037725
transform 1 0 19228 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_219
timestamp 1676037725
transform 1 0 21252 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_231
timestamp 1676037725
transform 1 0 22356 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_235
timestamp 1676037725
transform 1 0 22724 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_247
timestamp 1676037725
transform 1 0 23828 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_251
timestamp 1676037725
transform 1 0 24196 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_253
timestamp 1676037725
transform 1 0 24380 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_260
timestamp 1676037725
transform 1 0 25024 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_267
timestamp 1676037725
transform 1 0 25668 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_16_274
timestamp 1676037725
transform 1 0 26312 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_286
timestamp 1676037725
transform 1 0 27416 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_298
timestamp 1676037725
transform 1 0 28520 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_306
timestamp 1676037725
transform 1 0 29256 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_16_309
timestamp 1676037725
transform 1 0 29532 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_16_338
timestamp 1676037725
transform 1 0 32200 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_16_346
timestamp 1676037725
transform 1 0 32936 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_358
timestamp 1676037725
transform 1 0 34040 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_16_365
timestamp 1676037725
transform 1 0 34684 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_16_373
timestamp 1676037725
transform 1 0 35420 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_381
timestamp 1676037725
transform 1 0 36156 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_389
timestamp 1676037725
transform 1 0 36892 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_397
timestamp 1676037725
transform 1 0 37628 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_410
timestamp 1676037725
transform 1 0 38824 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_418
timestamp 1676037725
transform 1 0 39560 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_421
timestamp 1676037725
transform 1 0 39836 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_433
timestamp 1676037725
transform 1 0 40940 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_437
timestamp 1676037725
transform 1 0 41308 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_454
timestamp 1676037725
transform 1 0 42872 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_16_466
timestamp 1676037725
transform 1 0 43976 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_471
timestamp 1676037725
transform 1 0 44436 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_3
timestamp 1676037725
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_15
timestamp 1676037725
transform 1 0 2484 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_17_26
timestamp 1676037725
transform 1 0 3496 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_30
timestamp 1676037725
transform 1 0 3864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_34
timestamp 1676037725
transform 1 0 4232 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_54
timestamp 1676037725
transform 1 0 6072 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_17_57
timestamp 1676037725
transform 1 0 6348 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_63
timestamp 1676037725
transform 1 0 6900 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_73
timestamp 1676037725
transform 1 0 7820 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_17_86
timestamp 1676037725
transform 1 0 9016 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_101
timestamp 1676037725
transform 1 0 10396 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_17_109
timestamp 1676037725
transform 1 0 11132 0 -1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_17_113
timestamp 1676037725
transform 1 0 11500 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_125
timestamp 1676037725
transform 1 0 12604 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_17_147
timestamp 1676037725
transform 1 0 14628 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_17_154
timestamp 1676037725
transform 1 0 15272 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_166
timestamp 1676037725
transform 1 0 16376 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_169
timestamp 1676037725
transform 1 0 16652 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_180
timestamp 1676037725
transform 1 0 17664 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_17_192
timestamp 1676037725
transform 1 0 18768 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_198
timestamp 1676037725
transform 1 0 19320 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_211
timestamp 1676037725
transform 1 0 20516 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_222
timestamp 1676037725
transform 1 0 21528 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_225
timestamp 1676037725
transform 1 0 21804 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_232
timestamp 1676037725
transform 1 0 22448 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_17_239
timestamp 1676037725
transform 1 0 23092 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_251
timestamp 1676037725
transform 1 0 24196 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_257
timestamp 1676037725
transform 1 0 24748 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_278
timestamp 1676037725
transform 1 0 26680 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_281
timestamp 1676037725
transform 1 0 26956 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_293
timestamp 1676037725
transform 1 0 28060 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_17_303
timestamp 1676037725
transform 1 0 28980 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_313
timestamp 1676037725
transform 1 0 29900 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_17_333
timestamp 1676037725
transform 1 0 31740 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_337
timestamp 1676037725
transform 1 0 32108 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_344
timestamp 1676037725
transform 1 0 32752 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_353
timestamp 1676037725
transform 1 0 33580 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_373
timestamp 1676037725
transform 1 0 35420 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_380
timestamp 1676037725
transform 1 0 36064 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_390
timestamp 1676037725
transform 1 0 36984 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_393
timestamp 1676037725
transform 1 0 37260 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_403
timestamp 1676037725
transform 1 0 38180 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_17_416
timestamp 1676037725
transform 1 0 39376 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_17_428
timestamp 1676037725
transform 1 0 40480 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_434
timestamp 1676037725
transform 1 0 41032 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_444
timestamp 1676037725
transform 1 0 41952 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_17_449
timestamp 1676037725
transform 1 0 42412 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_461
timestamp 1676037725
transform 1 0 43516 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_3
timestamp 1676037725
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_15
timestamp 1676037725
transform 1 0 2484 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_19
timestamp 1676037725
transform 1 0 2852 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_23
timestamp 1676037725
transform 1 0 3220 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1676037725
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_29
timestamp 1676037725
transform 1 0 3772 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_33
timestamp 1676037725
transform 1 0 4140 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_43
timestamp 1676037725
transform 1 0 5060 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_63
timestamp 1676037725
transform 1 0 6900 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_67
timestamp 1676037725
transform 1 0 7268 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_18_77
timestamp 1676037725
transform 1 0 8188 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp 1676037725
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_85
timestamp 1676037725
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_97
timestamp 1676037725
transform 1 0 10028 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_101
timestamp 1676037725
transform 1 0 10396 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_121
timestamp 1676037725
transform 1 0 12236 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_138
timestamp 1676037725
transform 1 0 13800 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_18_141
timestamp 1676037725
transform 1 0 14076 0 1 11968
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_18_156
timestamp 1676037725
transform 1 0 15456 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_168
timestamp 1676037725
transform 1 0 16560 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_180
timestamp 1676037725
transform 1 0 17664 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_18_188
timestamp 1676037725
transform 1 0 18400 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_194
timestamp 1676037725
transform 1 0 18952 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_197
timestamp 1676037725
transform 1 0 19228 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_219
timestamp 1676037725
transform 1 0 21252 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_231
timestamp 1676037725
transform 1 0 22356 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_242
timestamp 1676037725
transform 1 0 23368 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_250
timestamp 1676037725
transform 1 0 24104 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_253
timestamp 1676037725
transform 1 0 24380 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_275
timestamp 1676037725
transform 1 0 26404 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_18_282
timestamp 1676037725
transform 1 0 27048 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_294
timestamp 1676037725
transform 1 0 28152 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_18_306
timestamp 1676037725
transform 1 0 29256 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_309
timestamp 1676037725
transform 1 0 29532 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_321
timestamp 1676037725
transform 1 0 30636 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_329
timestamp 1676037725
transform 1 0 31372 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_340
timestamp 1676037725
transform 1 0 32384 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_349
timestamp 1676037725
transform 1 0 33212 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_357
timestamp 1676037725
transform 1 0 33948 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_362
timestamp 1676037725
transform 1 0 34408 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_18_365
timestamp 1676037725
transform 1 0 34684 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_18_376
timestamp 1676037725
transform 1 0 35696 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_385
timestamp 1676037725
transform 1 0 36524 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_397
timestamp 1676037725
transform 1 0 37628 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_406
timestamp 1676037725
transform 1 0 38456 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_18_417
timestamp 1676037725
transform 1 0 39468 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_421
timestamp 1676037725
transform 1 0 39836 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_433
timestamp 1676037725
transform 1 0 40940 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_439
timestamp 1676037725
transform 1 0 41492 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_448
timestamp 1676037725
transform 1 0 42320 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_460
timestamp 1676037725
transform 1 0 43424 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_472
timestamp 1676037725
transform 1 0 44528 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_3
timestamp 1676037725
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_15
timestamp 1676037725
transform 1 0 2484 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_19
timestamp 1676037725
transform 1 0 2852 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_23
timestamp 1676037725
transform 1 0 3220 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_31
timestamp 1676037725
transform 1 0 3956 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_48
timestamp 1676037725
transform 1 0 5520 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_57
timestamp 1676037725
transform 1 0 6348 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_75
timestamp 1676037725
transform 1 0 8004 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_19_82
timestamp 1676037725
transform 1 0 8648 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_19_110
timestamp 1676037725
transform 1 0 11224 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_113
timestamp 1676037725
transform 1 0 11500 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_19_124
timestamp 1676037725
transform 1 0 12512 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_130
timestamp 1676037725
transform 1 0 13064 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_147
timestamp 1676037725
transform 1 0 14628 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_19_154
timestamp 1676037725
transform 1 0 15272 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_19_166
timestamp 1676037725
transform 1 0 16376 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_169
timestamp 1676037725
transform 1 0 16652 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_19_181
timestamp 1676037725
transform 1 0 17756 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_185
timestamp 1676037725
transform 1 0 18124 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_209
timestamp 1676037725
transform 1 0 20332 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_19_221
timestamp 1676037725
transform 1 0 21436 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_225
timestamp 1676037725
transform 1 0 21804 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_232
timestamp 1676037725
transform 1 0 22448 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_244
timestamp 1676037725
transform 1 0 23552 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_19_256
timestamp 1676037725
transform 1 0 24656 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_261
timestamp 1676037725
transform 1 0 25116 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_19_274
timestamp 1676037725
transform 1 0 26312 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_19_281
timestamp 1676037725
transform 1 0 26956 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_287
timestamp 1676037725
transform 1 0 27508 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_299
timestamp 1676037725
transform 1 0 28612 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_19_321
timestamp 1676037725
transform 1 0 30636 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_19_334
timestamp 1676037725
transform 1 0 31832 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_337
timestamp 1676037725
transform 1 0 32108 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_347
timestamp 1676037725
transform 1 0 33028 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_356
timestamp 1676037725
transform 1 0 33856 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_360
timestamp 1676037725
transform 1 0 34224 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_365
timestamp 1676037725
transform 1 0 34684 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_19_376
timestamp 1676037725
transform 1 0 35696 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_19_389
timestamp 1676037725
transform 1 0 36892 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_393
timestamp 1676037725
transform 1 0 37260 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_401
timestamp 1676037725
transform 1 0 37996 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_411
timestamp 1676037725
transform 1 0 38916 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_418
timestamp 1676037725
transform 1 0 39560 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_422
timestamp 1676037725
transform 1 0 39928 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_428
timestamp 1676037725
transform 1 0 40480 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_19_444
timestamp 1676037725
transform 1 0 41952 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_19_449
timestamp 1676037725
transform 1 0 42412 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_461
timestamp 1676037725
transform 1 0 43516 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_467
timestamp 1676037725
transform 1 0 44068 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_471
timestamp 1676037725
transform 1 0 44436 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_3
timestamp 1676037725
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_15
timestamp 1676037725
transform 1 0 2484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1676037725
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_20_29
timestamp 1676037725
transform 1 0 3772 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_35
timestamp 1676037725
transform 1 0 4324 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_39
timestamp 1676037725
transform 1 0 4692 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_59
timestamp 1676037725
transform 1 0 6532 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_20_72
timestamp 1676037725
transform 1 0 7728 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_85
timestamp 1676037725
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_20_97
timestamp 1676037725
transform 1 0 10028 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_108
timestamp 1676037725
transform 1 0 11040 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_20_128
timestamp 1676037725
transform 1 0 12880 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_20_141
timestamp 1676037725
transform 1 0 14076 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_148
timestamp 1676037725
transform 1 0 14720 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_160
timestamp 1676037725
transform 1 0 15824 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_20_172
timestamp 1676037725
transform 1 0 16928 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_194
timestamp 1676037725
transform 1 0 18952 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_197
timestamp 1676037725
transform 1 0 19228 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_207
timestamp 1676037725
transform 1 0 20148 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_217
timestamp 1676037725
transform 1 0 21068 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_224
timestamp 1676037725
transform 1 0 21712 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_228
timestamp 1676037725
transform 1 0 22080 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_234
timestamp 1676037725
transform 1 0 22632 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_242
timestamp 1676037725
transform 1 0 23368 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_247
timestamp 1676037725
transform 1 0 23828 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_251
timestamp 1676037725
transform 1 0 24196 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_253
timestamp 1676037725
transform 1 0 24380 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_275
timestamp 1676037725
transform 1 0 26404 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_20_282
timestamp 1676037725
transform 1 0 27048 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_294
timestamp 1676037725
transform 1 0 28152 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_20_303
timestamp 1676037725
transform 1 0 28980 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_307
timestamp 1676037725
transform 1 0 29348 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_309
timestamp 1676037725
transform 1 0 29532 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_20_315
timestamp 1676037725
transform 1 0 30084 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_20_330
timestamp 1676037725
transform 1 0 31464 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_335
timestamp 1676037725
transform 1 0 31924 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_345
timestamp 1676037725
transform 1 0 32844 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_20_352
timestamp 1676037725
transform 1 0 33488 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_365
timestamp 1676037725
transform 1 0 34684 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_20_376
timestamp 1676037725
transform 1 0 35696 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_385
timestamp 1676037725
transform 1 0 36524 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_20_405
timestamp 1676037725
transform 1 0 38364 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_20_417
timestamp 1676037725
transform 1 0 39468 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_421
timestamp 1676037725
transform 1 0 39836 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_429
timestamp 1676037725
transform 1 0 40572 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_449
timestamp 1676037725
transform 1 0 42412 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_20_459
timestamp 1676037725
transform 1 0 43332 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_20_471
timestamp 1676037725
transform 1 0 44436 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_3
timestamp 1676037725
transform 1 0 1380 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_8
timestamp 1676037725
transform 1 0 1840 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_20
timestamp 1676037725
transform 1 0 2944 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_32
timestamp 1676037725
transform 1 0 4048 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_49
timestamp 1676037725
transform 1 0 5612 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_55
timestamp 1676037725
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_57
timestamp 1676037725
transform 1 0 6348 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_68
timestamp 1676037725
transform 1 0 7360 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_80
timestamp 1676037725
transform 1 0 8464 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_92
timestamp 1676037725
transform 1 0 9568 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_104
timestamp 1676037725
transform 1 0 10672 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_21_113
timestamp 1676037725
transform 1 0 11500 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_121
timestamp 1676037725
transform 1 0 12236 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_126
timestamp 1676037725
transform 1 0 12696 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_21_146
timestamp 1676037725
transform 1 0 14536 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_158
timestamp 1676037725
transform 1 0 15640 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_166
timestamp 1676037725
transform 1 0 16376 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_21_169
timestamp 1676037725
transform 1 0 16652 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_21_178
timestamp 1676037725
transform 1 0 17480 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_202
timestamp 1676037725
transform 1 0 19688 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_212
timestamp 1676037725
transform 1 0 20608 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_21_221
timestamp 1676037725
transform 1 0 21436 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_225
timestamp 1676037725
transform 1 0 21804 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_229
timestamp 1676037725
transform 1 0 22172 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_233
timestamp 1676037725
transform 1 0 22540 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_253
timestamp 1676037725
transform 1 0 24380 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_266
timestamp 1676037725
transform 1 0 25576 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_270
timestamp 1676037725
transform 1 0 25944 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_276
timestamp 1676037725
transform 1 0 26496 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_281
timestamp 1676037725
transform 1 0 26956 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_292
timestamp 1676037725
transform 1 0 27968 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_312
timestamp 1676037725
transform 1 0 29808 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_21_324
timestamp 1676037725
transform 1 0 30912 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_21_334
timestamp 1676037725
transform 1 0 31832 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_337
timestamp 1676037725
transform 1 0 32108 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_21_361
timestamp 1676037725
transform 1 0 34316 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_365
timestamp 1676037725
transform 1 0 34684 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_369
timestamp 1676037725
transform 1 0 35052 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_21_376
timestamp 1676037725
transform 1 0 35696 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_21_390
timestamp 1676037725
transform 1 0 36984 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_393
timestamp 1676037725
transform 1 0 37260 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_399
timestamp 1676037725
transform 1 0 37812 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_21_406
timestamp 1676037725
transform 1 0 38456 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_418
timestamp 1676037725
transform 1 0 39560 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_446
timestamp 1676037725
transform 1 0 42136 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_449
timestamp 1676037725
transform 1 0 42412 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_461
timestamp 1676037725
transform 1 0 43516 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_3
timestamp 1676037725
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_15
timestamp 1676037725
transform 1 0 2484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 1676037725
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_29
timestamp 1676037725
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_41
timestamp 1676037725
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_53
timestamp 1676037725
transform 1 0 5980 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_65
timestamp 1676037725
transform 1 0 7084 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_77
timestamp 1676037725
transform 1 0 8188 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_83
timestamp 1676037725
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_85
timestamp 1676037725
transform 1 0 8924 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_93
timestamp 1676037725
transform 1 0 9660 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_111
timestamp 1676037725
transform 1 0 11316 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_123
timestamp 1676037725
transform 1 0 12420 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_135
timestamp 1676037725
transform 1 0 13524 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_139
timestamp 1676037725
transform 1 0 13892 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_141
timestamp 1676037725
transform 1 0 14076 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_153
timestamp 1676037725
transform 1 0 15180 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_165
timestamp 1676037725
transform 1 0 16284 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_177
timestamp 1676037725
transform 1 0 17388 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_183
timestamp 1676037725
transform 1 0 17940 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_187
timestamp 1676037725
transform 1 0 18308 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_194
timestamp 1676037725
transform 1 0 18952 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_197
timestamp 1676037725
transform 1 0 19228 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_22_202
timestamp 1676037725
transform 1 0 19688 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_208
timestamp 1676037725
transform 1 0 20240 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_225
timestamp 1676037725
transform 1 0 21804 0 1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_22_238
timestamp 1676037725
transform 1 0 23000 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_22_250
timestamp 1676037725
transform 1 0 24104 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_253
timestamp 1676037725
transform 1 0 24380 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_265
timestamp 1676037725
transform 1 0 25484 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_271
timestamp 1676037725
transform 1 0 26036 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_288
timestamp 1676037725
transform 1 0 27600 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_300
timestamp 1676037725
transform 1 0 28704 0 1 14144
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_22_309
timestamp 1676037725
transform 1 0 29532 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_321
timestamp 1676037725
transform 1 0 30636 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_327
timestamp 1676037725
transform 1 0 31188 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_344
timestamp 1676037725
transform 1 0 32752 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_356
timestamp 1676037725
transform 1 0 33856 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_365
timestamp 1676037725
transform 1 0 34684 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_22_370
timestamp 1676037725
transform 1 0 35144 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_378
timestamp 1676037725
transform 1 0 35880 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_384
timestamp 1676037725
transform 1 0 36432 0 1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_22_404
timestamp 1676037725
transform 1 0 38272 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_416
timestamp 1676037725
transform 1 0 39376 0 1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_22_421
timestamp 1676037725
transform 1 0 39836 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_440
timestamp 1676037725
transform 1 0 41584 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_22_447
timestamp 1676037725
transform 1 0 42228 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_22_456
timestamp 1676037725
transform 1 0 43056 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_22_464
timestamp 1676037725
transform 1 0 43792 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_471
timestamp 1676037725
transform 1 0 44436 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_23_3
timestamp 1676037725
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_15
timestamp 1676037725
transform 1 0 2484 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_27
timestamp 1676037725
transform 1 0 3588 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_39
timestamp 1676037725
transform 1 0 4692 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_51
timestamp 1676037725
transform 1 0 5796 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_55
timestamp 1676037725
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_57
timestamp 1676037725
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_69
timestamp 1676037725
transform 1 0 7452 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_81
timestamp 1676037725
transform 1 0 8556 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_93
timestamp 1676037725
transform 1 0 9660 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_105
timestamp 1676037725
transform 1 0 10764 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_111
timestamp 1676037725
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_113
timestamp 1676037725
transform 1 0 11500 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_125
timestamp 1676037725
transform 1 0 12604 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_137
timestamp 1676037725
transform 1 0 13708 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_149
timestamp 1676037725
transform 1 0 14812 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_161
timestamp 1676037725
transform 1 0 15916 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_167
timestamp 1676037725
transform 1 0 16468 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_169
timestamp 1676037725
transform 1 0 16652 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_181
timestamp 1676037725
transform 1 0 17756 0 -1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_23_205
timestamp 1676037725
transform 1 0 19964 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_217
timestamp 1676037725
transform 1 0 21068 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_223
timestamp 1676037725
transform 1 0 21620 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_225
timestamp 1676037725
transform 1 0 21804 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_23_233
timestamp 1676037725
transform 1 0 22540 0 -1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_23_245
timestamp 1676037725
transform 1 0 23644 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_257
timestamp 1676037725
transform 1 0 24748 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_278
timestamp 1676037725
transform 1 0 26680 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_23_281
timestamp 1676037725
transform 1 0 26956 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_293
timestamp 1676037725
transform 1 0 28060 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_305
timestamp 1676037725
transform 1 0 29164 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_317
timestamp 1676037725
transform 1 0 30268 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_23_329
timestamp 1676037725
transform 1 0 31372 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_334
timestamp 1676037725
transform 1 0 31832 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_337
timestamp 1676037725
transform 1 0 32108 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_347
timestamp 1676037725
transform 1 0 33028 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_357
timestamp 1676037725
transform 1 0 33948 0 -1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_23_366
timestamp 1676037725
transform 1 0 34776 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_378
timestamp 1676037725
transform 1 0 35880 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_382
timestamp 1676037725
transform 1 0 36248 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_23_386
timestamp 1676037725
transform 1 0 36616 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_23_393
timestamp 1676037725
transform 1 0 37260 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_23_398
timestamp 1676037725
transform 1 0 37720 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_410
timestamp 1676037725
transform 1 0 38824 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_422
timestamp 1676037725
transform 1 0 39928 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_434
timestamp 1676037725
transform 1 0 41032 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_446
timestamp 1676037725
transform 1 0 42136 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_23_449
timestamp 1676037725
transform 1 0 42412 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_461
timestamp 1676037725
transform 1 0 43516 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_24_3
timestamp 1676037725
transform 1 0 1380 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_9
timestamp 1676037725
transform 1 0 1932 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_21
timestamp 1676037725
transform 1 0 3036 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1676037725
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_29
timestamp 1676037725
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_41
timestamp 1676037725
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_53
timestamp 1676037725
transform 1 0 5980 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_65
timestamp 1676037725
transform 1 0 7084 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_77
timestamp 1676037725
transform 1 0 8188 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_83
timestamp 1676037725
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_85
timestamp 1676037725
transform 1 0 8924 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_97
timestamp 1676037725
transform 1 0 10028 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_109
timestamp 1676037725
transform 1 0 11132 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_121
timestamp 1676037725
transform 1 0 12236 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_133
timestamp 1676037725
transform 1 0 13340 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_139
timestamp 1676037725
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_141
timestamp 1676037725
transform 1 0 14076 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_153
timestamp 1676037725
transform 1 0 15180 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_165
timestamp 1676037725
transform 1 0 16284 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_177
timestamp 1676037725
transform 1 0 17388 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_189
timestamp 1676037725
transform 1 0 18492 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_195
timestamp 1676037725
transform 1 0 19044 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_197
timestamp 1676037725
transform 1 0 19228 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_209
timestamp 1676037725
transform 1 0 20332 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_221
timestamp 1676037725
transform 1 0 21436 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_233
timestamp 1676037725
transform 1 0 22540 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_245
timestamp 1676037725
transform 1 0 23644 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_251
timestamp 1676037725
transform 1 0 24196 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_253
timestamp 1676037725
transform 1 0 24380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_265
timestamp 1676037725
transform 1 0 25484 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_277
timestamp 1676037725
transform 1 0 26588 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_289
timestamp 1676037725
transform 1 0 27692 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_301
timestamp 1676037725
transform 1 0 28796 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_307
timestamp 1676037725
transform 1 0 29348 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_309
timestamp 1676037725
transform 1 0 29532 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_321
timestamp 1676037725
transform 1 0 30636 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_333
timestamp 1676037725
transform 1 0 31740 0 1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_24_342
timestamp 1676037725
transform 1 0 32568 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_354
timestamp 1676037725
transform 1 0 33672 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_362
timestamp 1676037725
transform 1 0 34408 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_365
timestamp 1676037725
transform 1 0 34684 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_377
timestamp 1676037725
transform 1 0 35788 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_389
timestamp 1676037725
transform 1 0 36892 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_401
timestamp 1676037725
transform 1 0 37996 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_413
timestamp 1676037725
transform 1 0 39100 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_419
timestamp 1676037725
transform 1 0 39652 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_421
timestamp 1676037725
transform 1 0 39836 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_433
timestamp 1676037725
transform 1 0 40940 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_445
timestamp 1676037725
transform 1 0 42044 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_457
timestamp 1676037725
transform 1 0 43148 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_469
timestamp 1676037725
transform 1 0 44252 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_3
timestamp 1676037725
transform 1 0 1380 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_8
timestamp 1676037725
transform 1 0 1840 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_20
timestamp 1676037725
transform 1 0 2944 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_32
timestamp 1676037725
transform 1 0 4048 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_44
timestamp 1676037725
transform 1 0 5152 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_57
timestamp 1676037725
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_69
timestamp 1676037725
transform 1 0 7452 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_81
timestamp 1676037725
transform 1 0 8556 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_93
timestamp 1676037725
transform 1 0 9660 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_105
timestamp 1676037725
transform 1 0 10764 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_111
timestamp 1676037725
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_113
timestamp 1676037725
transform 1 0 11500 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_125
timestamp 1676037725
transform 1 0 12604 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_137
timestamp 1676037725
transform 1 0 13708 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_149
timestamp 1676037725
transform 1 0 14812 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_161
timestamp 1676037725
transform 1 0 15916 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_167
timestamp 1676037725
transform 1 0 16468 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_169
timestamp 1676037725
transform 1 0 16652 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_181
timestamp 1676037725
transform 1 0 17756 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_193
timestamp 1676037725
transform 1 0 18860 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_205
timestamp 1676037725
transform 1 0 19964 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_217
timestamp 1676037725
transform 1 0 21068 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_223
timestamp 1676037725
transform 1 0 21620 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_225
timestamp 1676037725
transform 1 0 21804 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_237
timestamp 1676037725
transform 1 0 22908 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_249
timestamp 1676037725
transform 1 0 24012 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_261
timestamp 1676037725
transform 1 0 25116 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_273
timestamp 1676037725
transform 1 0 26220 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_279
timestamp 1676037725
transform 1 0 26772 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_281
timestamp 1676037725
transform 1 0 26956 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_293
timestamp 1676037725
transform 1 0 28060 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_305
timestamp 1676037725
transform 1 0 29164 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_317
timestamp 1676037725
transform 1 0 30268 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_329
timestamp 1676037725
transform 1 0 31372 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_335
timestamp 1676037725
transform 1 0 31924 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_337
timestamp 1676037725
transform 1 0 32108 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_349
timestamp 1676037725
transform 1 0 33212 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_361
timestamp 1676037725
transform 1 0 34316 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_373
timestamp 1676037725
transform 1 0 35420 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_385
timestamp 1676037725
transform 1 0 36524 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_391
timestamp 1676037725
transform 1 0 37076 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_393
timestamp 1676037725
transform 1 0 37260 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_405
timestamp 1676037725
transform 1 0 38364 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_417
timestamp 1676037725
transform 1 0 39468 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_429
timestamp 1676037725
transform 1 0 40572 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_441
timestamp 1676037725
transform 1 0 41676 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_447
timestamp 1676037725
transform 1 0 42228 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_449
timestamp 1676037725
transform 1 0 42412 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_456
timestamp 1676037725
transform 1 0 43056 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_25_460
timestamp 1676037725
transform 1 0 43424 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_471
timestamp 1676037725
transform 1 0 44436 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_3
timestamp 1676037725
transform 1 0 1380 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_9
timestamp 1676037725
transform 1 0 1932 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_21
timestamp 1676037725
transform 1 0 3036 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 1676037725
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_29
timestamp 1676037725
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_41
timestamp 1676037725
transform 1 0 4876 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_53
timestamp 1676037725
transform 1 0 5980 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_65
timestamp 1676037725
transform 1 0 7084 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_77
timestamp 1676037725
transform 1 0 8188 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_83
timestamp 1676037725
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_85
timestamp 1676037725
transform 1 0 8924 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_97
timestamp 1676037725
transform 1 0 10028 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_109
timestamp 1676037725
transform 1 0 11132 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_121
timestamp 1676037725
transform 1 0 12236 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_133
timestamp 1676037725
transform 1 0 13340 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_139
timestamp 1676037725
transform 1 0 13892 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_26_141
timestamp 1676037725
transform 1 0 14076 0 1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_26_147
timestamp 1676037725
transform 1 0 14628 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_159
timestamp 1676037725
transform 1 0 15732 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_171
timestamp 1676037725
transform 1 0 16836 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_183
timestamp 1676037725
transform 1 0 17940 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_195
timestamp 1676037725
transform 1 0 19044 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_197
timestamp 1676037725
transform 1 0 19228 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_209
timestamp 1676037725
transform 1 0 20332 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_221
timestamp 1676037725
transform 1 0 21436 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_233
timestamp 1676037725
transform 1 0 22540 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_245
timestamp 1676037725
transform 1 0 23644 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_251
timestamp 1676037725
transform 1 0 24196 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_253
timestamp 1676037725
transform 1 0 24380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_265
timestamp 1676037725
transform 1 0 25484 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_277
timestamp 1676037725
transform 1 0 26588 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_289
timestamp 1676037725
transform 1 0 27692 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_295
timestamp 1676037725
transform 1 0 28244 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_299
timestamp 1676037725
transform 1 0 28612 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_307
timestamp 1676037725
transform 1 0 29348 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_309
timestamp 1676037725
transform 1 0 29532 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_321
timestamp 1676037725
transform 1 0 30636 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_333
timestamp 1676037725
transform 1 0 31740 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_345
timestamp 1676037725
transform 1 0 32844 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_357
timestamp 1676037725
transform 1 0 33948 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_363
timestamp 1676037725
transform 1 0 34500 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_365
timestamp 1676037725
transform 1 0 34684 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_377
timestamp 1676037725
transform 1 0 35788 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_389
timestamp 1676037725
transform 1 0 36892 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_401
timestamp 1676037725
transform 1 0 37996 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_413
timestamp 1676037725
transform 1 0 39100 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_419
timestamp 1676037725
transform 1 0 39652 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_421
timestamp 1676037725
transform 1 0 39836 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_433
timestamp 1676037725
transform 1 0 40940 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_445
timestamp 1676037725
transform 1 0 42044 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_457
timestamp 1676037725
transform 1 0 43148 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_464
timestamp 1676037725
transform 1 0 43792 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_471
timestamp 1676037725
transform 1 0 44436 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_3
timestamp 1676037725
transform 1 0 1380 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_9
timestamp 1676037725
transform 1 0 1932 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_17
timestamp 1676037725
transform 1 0 2668 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_21
timestamp 1676037725
transform 1 0 3036 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_26
timestamp 1676037725
transform 1 0 3496 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_27_29
timestamp 1676037725
transform 1 0 3772 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_37
timestamp 1676037725
transform 1 0 4508 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_42
timestamp 1676037725
transform 1 0 4968 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_54
timestamp 1676037725
transform 1 0 6072 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_57
timestamp 1676037725
transform 1 0 6348 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_27_62
timestamp 1676037725
transform 1 0 6808 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_70
timestamp 1676037725
transform 1 0 7544 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_27_76
timestamp 1676037725
transform 1 0 8096 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_27_85
timestamp 1676037725
transform 1 0 8924 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_93
timestamp 1676037725
transform 1 0 9660 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_97
timestamp 1676037725
transform 1 0 10028 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_27_109
timestamp 1676037725
transform 1 0 11132 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_113
timestamp 1676037725
transform 1 0 11500 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_27_119
timestamp 1676037725
transform 1 0 12052 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_127
timestamp 1676037725
transform 1 0 12788 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_27_132
timestamp 1676037725
transform 1 0 13248 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_141
timestamp 1676037725
transform 1 0 14076 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_27_146
timestamp 1676037725
transform 1 0 14536 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_158
timestamp 1676037725
transform 1 0 15640 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_166
timestamp 1676037725
transform 1 0 16376 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_27_169
timestamp 1676037725
transform 1 0 16652 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_177
timestamp 1676037725
transform 1 0 17388 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_182
timestamp 1676037725
transform 1 0 17848 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_194
timestamp 1676037725
transform 1 0 18952 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_197
timestamp 1676037725
transform 1 0 19228 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_27_202
timestamp 1676037725
transform 1 0 19688 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_210
timestamp 1676037725
transform 1 0 20424 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_27_217
timestamp 1676037725
transform 1 0 21068 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_223
timestamp 1676037725
transform 1 0 21620 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_225
timestamp 1676037725
transform 1 0 21804 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_233
timestamp 1676037725
transform 1 0 22540 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_237
timestamp 1676037725
transform 1 0 22908 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_27_249
timestamp 1676037725
transform 1 0 24012 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_253
timestamp 1676037725
transform 1 0 24380 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_27_258
timestamp 1676037725
transform 1 0 24840 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_266
timestamp 1676037725
transform 1 0 25576 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_27_272
timestamp 1676037725
transform 1 0 26128 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_27_281
timestamp 1676037725
transform 1 0 26956 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_289
timestamp 1676037725
transform 1 0 27692 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_293
timestamp 1676037725
transform 1 0 28060 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_27_305
timestamp 1676037725
transform 1 0 29164 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_309
timestamp 1676037725
transform 1 0 29532 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_27_314
timestamp 1676037725
transform 1 0 29992 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_322
timestamp 1676037725
transform 1 0 30728 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_27_328
timestamp 1676037725
transform 1 0 31280 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_337
timestamp 1676037725
transform 1 0 32108 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_27_343
timestamp 1676037725
transform 1 0 32660 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_355
timestamp 1676037725
transform 1 0 33764 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_363
timestamp 1676037725
transform 1 0 34500 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_365
timestamp 1676037725
transform 1 0 34684 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_370
timestamp 1676037725
transform 1 0 35144 0 -1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_27_377
timestamp 1676037725
transform 1 0 35788 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_27_389
timestamp 1676037725
transform 1 0 36892 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_393
timestamp 1676037725
transform 1 0 37260 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_27_398
timestamp 1676037725
transform 1 0 37720 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_406
timestamp 1676037725
transform 1 0 38456 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_27_413
timestamp 1676037725
transform 1 0 39100 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_419
timestamp 1676037725
transform 1 0 39652 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_421
timestamp 1676037725
transform 1 0 39836 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_429
timestamp 1676037725
transform 1 0 40572 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_434
timestamp 1676037725
transform 1 0 41032 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_446
timestamp 1676037725
transform 1 0 42136 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_449
timestamp 1676037725
transform 1 0 42412 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_27_454
timestamp 1676037725
transform 1 0 42872 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_27_463
timestamp 1676037725
transform 1 0 43700 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_471
timestamp 1676037725
transform 1 0 44436 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1676037725
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1676037725
transform -1 0 44896 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1676037725
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1676037725
transform -1 0 44896 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1676037725
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1676037725
transform -1 0 44896 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1676037725
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1676037725
transform -1 0 44896 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1676037725
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1676037725
transform -1 0 44896 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1676037725
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1676037725
transform -1 0 44896 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1676037725
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1676037725
transform -1 0 44896 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1676037725
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1676037725
transform -1 0 44896 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1676037725
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1676037725
transform -1 0 44896 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1676037725
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1676037725
transform -1 0 44896 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1676037725
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1676037725
transform -1 0 44896 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1676037725
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1676037725
transform -1 0 44896 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1676037725
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1676037725
transform -1 0 44896 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1676037725
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1676037725
transform -1 0 44896 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1676037725
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1676037725
transform -1 0 44896 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1676037725
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1676037725
transform -1 0 44896 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1676037725
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1676037725
transform -1 0 44896 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1676037725
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1676037725
transform -1 0 44896 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1676037725
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1676037725
transform -1 0 44896 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1676037725
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1676037725
transform -1 0 44896 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1676037725
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1676037725
transform -1 0 44896 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1676037725
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1676037725
transform -1 0 44896 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1676037725
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1676037725
transform -1 0 44896 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1676037725
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1676037725
transform -1 0 44896 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1676037725
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1676037725
transform -1 0 44896 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1676037725
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1676037725
transform -1 0 44896 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1676037725
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1676037725
transform -1 0 44896 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1676037725
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1676037725
transform -1 0 44896 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_56 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_57
timestamp 1676037725
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_58
timestamp 1676037725
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_59
timestamp 1676037725
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_60
timestamp 1676037725
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_61
timestamp 1676037725
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_62
timestamp 1676037725
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_63
timestamp 1676037725
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_64
timestamp 1676037725
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_65
timestamp 1676037725
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_66
timestamp 1676037725
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_67
timestamp 1676037725
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_68
timestamp 1676037725
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_69
timestamp 1676037725
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_70
timestamp 1676037725
transform 1 0 39744 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_71
timestamp 1676037725
transform 1 0 42320 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_72
timestamp 1676037725
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_73
timestamp 1676037725
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_74
timestamp 1676037725
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_75
timestamp 1676037725
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_76
timestamp 1676037725
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_77
timestamp 1676037725
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_78
timestamp 1676037725
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_79
timestamp 1676037725
transform 1 0 42320 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_80
timestamp 1676037725
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_81
timestamp 1676037725
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_82
timestamp 1676037725
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_83
timestamp 1676037725
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_84
timestamp 1676037725
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_85
timestamp 1676037725
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_86
timestamp 1676037725
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_87
timestamp 1676037725
transform 1 0 39744 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_88
timestamp 1676037725
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_89
timestamp 1676037725
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_90
timestamp 1676037725
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_91
timestamp 1676037725
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_92
timestamp 1676037725
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_93
timestamp 1676037725
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94
timestamp 1676037725
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1676037725
transform 1 0 42320 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 1676037725
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 1676037725
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 1676037725
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 1676037725
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 1676037725
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_101
timestamp 1676037725
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102
timestamp 1676037725
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 1676037725
transform 1 0 39744 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 1676037725
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 1676037725
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 1676037725
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 1676037725
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 1676037725
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1676037725
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1676037725
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1676037725
transform 1 0 42320 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1676037725
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1676037725
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1676037725
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1676037725
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 1676037725
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1676037725
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1676037725
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1676037725
transform 1 0 39744 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1676037725
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_121
timestamp 1676037725
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_122
timestamp 1676037725
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_123
timestamp 1676037725
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_124
timestamp 1676037725
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_125
timestamp 1676037725
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_126
timestamp 1676037725
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_127
timestamp 1676037725
transform 1 0 42320 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_128
timestamp 1676037725
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_129
timestamp 1676037725
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130
timestamp 1676037725
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1676037725
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1676037725
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1676037725
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1676037725
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1676037725
transform 1 0 39744 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1676037725
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1676037725
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1676037725
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1676037725
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1676037725
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1676037725
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1676037725
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1676037725
transform 1 0 42320 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1676037725
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1676037725
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1676037725
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1676037725
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1676037725
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1676037725
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1676037725
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1676037725
transform 1 0 39744 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1676037725
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1676037725
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1676037725
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1676037725
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1676037725
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1676037725
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1676037725
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1676037725
transform 1 0 42320 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1676037725
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1676037725
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1676037725
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1676037725
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1676037725
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1676037725
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1676037725
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1676037725
transform 1 0 39744 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1676037725
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1676037725
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1676037725
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1676037725
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1676037725
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1676037725
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1676037725
transform 1 0 37168 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1676037725
transform 1 0 42320 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1676037725
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1676037725
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1676037725
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1676037725
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1676037725
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1676037725
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1676037725
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1676037725
transform 1 0 39744 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1676037725
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1676037725
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1676037725
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1676037725
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1676037725
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1676037725
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1676037725
transform 1 0 37168 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1676037725
transform 1 0 42320 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1676037725
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1676037725
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1676037725
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1676037725
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1676037725
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1676037725
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1676037725
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1676037725
transform 1 0 39744 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1676037725
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1676037725
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1676037725
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1676037725
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1676037725
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1676037725
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1676037725
transform 1 0 37168 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1676037725
transform 1 0 42320 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1676037725
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1676037725
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1676037725
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1676037725
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1676037725
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1676037725
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1676037725
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1676037725
transform 1 0 39744 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1676037725
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1676037725
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1676037725
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1676037725
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1676037725
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1676037725
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1676037725
transform 1 0 37168 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1676037725
transform 1 0 42320 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1676037725
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1676037725
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1676037725
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1676037725
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1676037725
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1676037725
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1676037725
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1676037725
transform 1 0 39744 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1676037725
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1676037725
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1676037725
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1676037725
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1676037725
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1676037725
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1676037725
transform 1 0 37168 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1676037725
transform 1 0 42320 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1676037725
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1676037725
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1676037725
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1676037725
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1676037725
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1676037725
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1676037725
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1676037725
transform 1 0 39744 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1676037725
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1676037725
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1676037725
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1676037725
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1676037725
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1676037725
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1676037725
transform 1 0 37168 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1676037725
transform 1 0 42320 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1676037725
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1676037725
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1676037725
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1676037725
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1676037725
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1676037725
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1676037725
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1676037725
transform 1 0 39744 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1676037725
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1676037725
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1676037725
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1676037725
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1676037725
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1676037725
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1676037725
transform 1 0 37168 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1676037725
transform 1 0 42320 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1676037725
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1676037725
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1676037725
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1676037725
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1676037725
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1676037725
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1676037725
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1676037725
transform 1 0 39744 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1676037725
transform 1 0 3680 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1676037725
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1676037725
transform 1 0 8832 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1676037725
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1676037725
transform 1 0 13984 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1676037725
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1676037725
transform 1 0 19136 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1676037725
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1676037725
transform 1 0 24288 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1676037725
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1676037725
transform 1 0 29440 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1676037725
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1676037725
transform 1 0 34592 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1676037725
transform 1 0 37168 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1676037725
transform 1 0 39744 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1676037725
transform 1 0 42320 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _345_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 31372 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _346_
timestamp 1676037725
transform 1 0 35512 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _347_
timestamp 1676037725
transform 1 0 34868 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _348_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 33580 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _349_
timestamp 1676037725
transform 1 0 37444 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _350_
timestamp 1676037725
transform 1 0 38456 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _351_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 34132 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _352_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 35236 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _353_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 38088 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _354_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 35512 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _355_
timestamp 1676037725
transform 1 0 31188 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _356_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 33856 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__o2bb2a_1  _357_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 32660 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _358_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 32752 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__nand3b_1  _359_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 34868 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__a211oi_1  _360_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 33764 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_2  _361_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 31372 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _362_
timestamp 1676037725
transform 1 0 36156 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _363_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 40020 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _364_
timestamp 1676037725
transform 1 0 41584 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _365_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 38272 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _366_
timestamp 1676037725
transform 1 0 38916 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _367_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 35880 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _368_
timestamp 1676037725
transform 1 0 32016 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__a21boi_1  _369_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 33396 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _370_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 32292 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__a221oi_1  _371_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 32384 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _372_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 36524 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _373_
timestamp 1676037725
transform 1 0 35972 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _374_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 35052 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _375_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 39284 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _376_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 39100 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _377_
timestamp 1676037725
transform 1 0 38456 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _378_
timestamp 1676037725
transform 1 0 38364 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _379_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 40848 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _380_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 40296 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _381_
timestamp 1676037725
transform 1 0 40020 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _382_
timestamp 1676037725
transform 1 0 41032 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _383_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 39468 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _384_
timestamp 1676037725
transform 1 0 40388 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _385_
timestamp 1676037725
transform 1 0 41216 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _386_
timestamp 1676037725
transform 1 0 39192 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _387_
timestamp 1676037725
transform 1 0 38732 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _388_
timestamp 1676037725
transform 1 0 17480 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _389_
timestamp 1676037725
transform 1 0 16836 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _390_
timestamp 1676037725
transform 1 0 16836 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _391_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 17296 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _392_
timestamp 1676037725
transform 1 0 15824 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _393_
timestamp 1676037725
transform 1 0 18492 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _394_
timestamp 1676037725
transform 1 0 19044 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _395_
timestamp 1676037725
transform 1 0 24840 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _396_
timestamp 1676037725
transform 1 0 23828 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _397_
timestamp 1676037725
transform 1 0 18124 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _398_
timestamp 1676037725
transform 1 0 15824 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _399_
timestamp 1676037725
transform 1 0 18032 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _400_
timestamp 1676037725
transform 1 0 16928 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _401_
timestamp 1676037725
transform 1 0 16836 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _402_
timestamp 1676037725
transform 1 0 16192 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _403_
timestamp 1676037725
transform 1 0 19412 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _404_
timestamp 1676037725
transform 1 0 18676 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _405_
timestamp 1676037725
transform 1 0 25576 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _406_
timestamp 1676037725
transform 1 0 25208 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _407_
timestamp 1676037725
transform 1 0 20700 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _408_
timestamp 1676037725
transform 1 0 19044 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _409_
timestamp 1676037725
transform 1 0 19688 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _410_
timestamp 1676037725
transform 1 0 20700 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _411_
timestamp 1676037725
transform 1 0 24196 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _412_
timestamp 1676037725
transform 1 0 22632 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_1  _413_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 19412 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _414_
timestamp 1676037725
transform 1 0 15272 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _415_
timestamp 1676037725
transform 1 0 19688 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _416_
timestamp 1676037725
transform 1 0 24564 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _417_
timestamp 1676037725
transform 1 0 19688 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__or3b_1  _418_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 20700 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _419_
timestamp 1676037725
transform 1 0 14536 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__o2bb2a_1  _420_
timestamp 1676037725
transform 1 0 17020 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _421_
timestamp 1676037725
transform 1 0 18124 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__or4b_1  _422_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 19596 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _423_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 19964 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _424_
timestamp 1676037725
transform 1 0 19688 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _425_
timestamp 1676037725
transform 1 0 19044 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _426_
timestamp 1676037725
transform 1 0 19596 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _427_
timestamp 1676037725
transform 1 0 21436 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _428_
timestamp 1676037725
transform 1 0 35420 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__and4b_1  _429_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 40204 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__and4b_1  _430_
timestamp 1676037725
transform 1 0 37444 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _431_
timestamp 1676037725
transform 1 0 32752 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _432_
timestamp 1676037725
transform 1 0 40756 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _433_
timestamp 1676037725
transform 1 0 42596 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _434_
timestamp 1676037725
transform 1 0 35420 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _435_
timestamp 1676037725
transform 1 0 38180 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _436_
timestamp 1676037725
transform 1 0 42780 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _437_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 39284 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__a221oi_1  _438_
timestamp 1676037725
transform 1 0 38824 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__o2111a_1  _439_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 38548 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _440_
timestamp 1676037725
transform 1 0 34776 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _441_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 36064 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _442_
timestamp 1676037725
transform 1 0 36064 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _443_
timestamp 1676037725
transform 1 0 35420 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _444_
timestamp 1676037725
transform 1 0 30820 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _445_
timestamp 1676037725
transform 1 0 36064 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _446_
timestamp 1676037725
transform 1 0 38640 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _447_
timestamp 1676037725
transform 1 0 31556 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _448_
timestamp 1676037725
transform 1 0 37996 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__o211a_1  _449_
timestamp 1676037725
transform 1 0 36892 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _450_
timestamp 1676037725
transform 1 0 39284 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__and4b_1  _451_
timestamp 1676037725
transform 1 0 32292 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _452_
timestamp 1676037725
transform -1 0 32844 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _453_
timestamp 1676037725
transform 1 0 33212 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _454_
timestamp 1676037725
transform 1 0 37444 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__or4b_1  _455_
timestamp 1676037725
transform 1 0 33120 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__a21bo_1  _456_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 32292 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _457_
timestamp 1676037725
transform 1 0 32292 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _458_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 29716 0 1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__nand2_1  _459_
timestamp 1676037725
transform 1 0 22816 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _460_
timestamp 1676037725
transform 1 0 22724 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _461_
timestamp 1676037725
transform 1 0 20056 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _462_
timestamp 1676037725
transform 1 0 25392 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _463_
timestamp 1676037725
transform 1 0 24840 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _464_
timestamp 1676037725
transform 1 0 26036 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__a31oi_1  _465_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 24564 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _466_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 20700 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _467_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 34040 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _468_
timestamp 1676037725
transform 1 0 31556 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _469_
timestamp 1676037725
transform 1 0 30820 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__a32o_1  _470_
timestamp 1676037725
transform 1 0 21620 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _471_
timestamp 1676037725
transform 1 0 2116 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _472_
timestamp 1676037725
transform 1 0 15272 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _473_
timestamp 1676037725
transform 1 0 14996 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _474_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 27140 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_2  _475_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 9108 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _476_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 9476 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _477_
timestamp 1676037725
transform 1 0 6532 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _478_
timestamp 1676037725
transform -1 0 43056 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _479_
timestamp 1676037725
transform 1 0 9568 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _480_
timestamp 1676037725
transform -1 0 34500 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _481_
timestamp 1676037725
transform 1 0 14536 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _482_
timestamp 1676037725
transform 1 0 16100 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _483_
timestamp 1676037725
transform 1 0 9200 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _484_
timestamp 1676037725
transform 1 0 42780 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _485_
timestamp 1676037725
transform 1 0 4876 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _486_
timestamp 1676037725
transform 1 0 5704 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _487_
timestamp 1676037725
transform 1 0 5796 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _488_
timestamp 1676037725
transform 1 0 7544 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _489_
timestamp 1676037725
transform 1 0 3036 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _490_
timestamp 1676037725
transform 1 0 2944 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _491_
timestamp 1676037725
transform 1 0 27232 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _492_
timestamp 1676037725
transform 1 0 27140 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _493_
timestamp 1676037725
transform 1 0 28336 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _494_
timestamp 1676037725
transform 1 0 14260 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _495_
timestamp 1676037725
transform 1 0 13524 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _496_
timestamp 1676037725
transform 1 0 14352 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _497_
timestamp 1676037725
transform 1 0 25852 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _498_
timestamp 1676037725
transform 1 0 24748 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _499_
timestamp 1676037725
transform 1 0 2944 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _500_
timestamp 1676037725
transform 1 0 22816 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _501_
timestamp 1676037725
transform 1 0 22172 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _502_
timestamp 1676037725
transform 1 0 22264 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _503_
timestamp 1676037725
transform 1 0 32568 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _504_
timestamp 1676037725
transform 1 0 32292 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _505_
timestamp 1676037725
transform 1 0 22172 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _506_
timestamp 1676037725
transform 1 0 23552 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _507_
timestamp 1676037725
transform 1 0 21988 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _508_
timestamp 1676037725
transform 1 0 22448 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _509_
timestamp 1676037725
transform 1 0 20976 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _510_
timestamp 1676037725
transform 1 0 18032 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _511_
timestamp 1676037725
transform 1 0 25852 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _512_
timestamp 1676037725
transform 1 0 27140 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _513_
timestamp 1676037725
transform 1 0 26036 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _514_
timestamp 1676037725
transform 1 0 26772 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _515_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 21988 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _516_
timestamp 1676037725
transform 1 0 22264 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _517_
timestamp 1676037725
transform 1 0 22724 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _518_
timestamp 1676037725
transform 1 0 22724 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _519_
timestamp 1676037725
transform 1 0 30636 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _520_
timestamp 1676037725
transform 1 0 31464 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _521_
timestamp 1676037725
transform 1 0 21988 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  _522_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 31096 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _523_
timestamp 1676037725
transform 1 0 20700 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _524_
timestamp 1676037725
transform 1 0 32292 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _525_
timestamp 1676037725
transform 1 0 19412 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _526_
timestamp 1676037725
transform 1 0 17848 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _527_
timestamp 1676037725
transform 1 0 18676 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _528_
timestamp 1676037725
transform 1 0 22080 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _529_
timestamp 1676037725
transform 1 0 25392 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _530_
timestamp 1676037725
transform 1 0 18676 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _531_
timestamp 1676037725
transform 1 0 32936 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _532_
timestamp 1676037725
transform 1 0 17204 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _533_
timestamp 1676037725
transform 1 0 24656 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _534_
timestamp 1676037725
transform 1 0 24564 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _535_
timestamp 1676037725
transform 1 0 23552 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _536_
timestamp 1676037725
transform 1 0 26036 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _537_
timestamp 1676037725
transform 1 0 26772 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _538_
timestamp 1676037725
transform 1 0 29808 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _539_
timestamp 1676037725
transform 1 0 25852 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _540_
timestamp 1676037725
transform 1 0 16928 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _541_
timestamp 1676037725
transform 1 0 16836 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _542_
timestamp 1676037725
transform 1 0 15456 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _543_
timestamp 1676037725
transform 1 0 14628 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _544_
timestamp 1676037725
transform 1 0 12972 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _545_
timestamp 1676037725
transform 1 0 14996 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _546_
timestamp 1676037725
transform 1 0 11684 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _547_
timestamp 1676037725
transform 1 0 10212 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _548_
timestamp 1676037725
transform 1 0 10120 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _549_
timestamp 1676037725
transform 1 0 7360 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _550_
timestamp 1676037725
transform 1 0 6900 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _551_
timestamp 1676037725
transform 1 0 8372 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _552_
timestamp 1676037725
transform 1 0 6992 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _553_
timestamp 1676037725
transform 1 0 6716 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _554_
timestamp 1676037725
transform 1 0 5980 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _555_
timestamp 1676037725
transform 1 0 8188 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _556_
timestamp 1676037725
transform 1 0 4232 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _557_
timestamp 1676037725
transform 1 0 3956 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _558_
timestamp 1676037725
transform 1 0 10304 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _559_
timestamp 1676037725
transform 1 0 9108 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _560_
timestamp 1676037725
transform 1 0 10120 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _561_
timestamp 1676037725
transform 1 0 25576 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _562_
timestamp 1676037725
transform 1 0 19412 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _563_
timestamp 1676037725
transform 1 0 16100 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _564_
timestamp 1676037725
transform 1 0 17572 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _565_
timestamp 1676037725
transform 1 0 16468 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _566_
timestamp 1676037725
transform 1 0 25576 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _567_
timestamp 1676037725
transform 1 0 23736 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _568_
timestamp 1676037725
transform 1 0 18308 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _569_
timestamp 1676037725
transform 1 0 18676 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _570__1
timestamp 1676037725
transform 1 0 14536 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _571__2
timestamp 1676037725
transform 1 0 16836 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _572__3
timestamp 1676037725
transform 1 0 19412 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _573_
timestamp 1676037725
transform 1 0 32384 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _574_
timestamp 1676037725
transform 1 0 32384 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _575_
timestamp 1676037725
transform 1 0 35420 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _576_
timestamp 1676037725
transform 1 0 34132 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _577_
timestamp 1676037725
transform 1 0 34868 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _578_
timestamp 1676037725
transform 1 0 33948 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _579_
timestamp 1676037725
transform 1 0 37444 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _580_
timestamp 1676037725
transform 1 0 37536 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _581_
timestamp 1676037725
transform 1 0 30360 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _582_
timestamp 1676037725
transform 1 0 28612 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _583_
timestamp 1676037725
transform 1 0 27232 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _584_
timestamp 1676037725
transform 1 0 26128 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _585_
timestamp 1676037725
transform 1 0 27416 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _586_
timestamp 1676037725
transform 1 0 28612 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _587_
timestamp 1676037725
transform 1 0 29716 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _588_
timestamp 1676037725
transform 1 0 27968 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _589_
timestamp 1676037725
transform 1 0 28980 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _590_
timestamp 1676037725
transform 1 0 28704 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _591_
timestamp 1676037725
transform 1 0 29716 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _592_
timestamp 1676037725
transform 1 0 30176 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _593_
timestamp 1676037725
transform 1 0 31464 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _594_
timestamp 1676037725
transform 1 0 32108 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__nor3_1  _595_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 31464 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _596_
timestamp 1676037725
transform 1 0 34316 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _597_
timestamp 1676037725
transform 1 0 34868 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _598_
timestamp 1676037725
transform 1 0 33396 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _599_
timestamp 1676037725
transform 1 0 36340 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _600_
timestamp 1676037725
transform 1 0 35972 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__and4b_1  _601_
timestamp 1676037725
transform 1 0 36248 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _602_
timestamp 1676037725
transform 1 0 37444 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _603_
timestamp 1676037725
transform 1 0 33396 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _604_
timestamp 1676037725
transform 1 0 34316 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _605_
timestamp 1676037725
transform 1 0 38364 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _606_
timestamp 1676037725
transform 1 0 37444 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _607_
timestamp 1676037725
transform 1 0 37996 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _608_
timestamp 1676037725
transform 1 0 39192 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__a211oi_1  _609_
timestamp 1676037725
transform 1 0 36432 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _610_
timestamp 1676037725
transform 1 0 36340 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _611_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 37260 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__and3b_1  _612_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 35972 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _613_
timestamp 1676037725
transform 1 0 36708 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _614_
timestamp 1676037725
transform 1 0 35788 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _615_
timestamp 1676037725
transform 1 0 35236 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _616_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 31740 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a211oi_1  _617_
timestamp 1676037725
transform 1 0 34868 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _618_
timestamp 1676037725
transform 1 0 31004 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _619_
timestamp 1676037725
transform 1 0 29348 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _620_
timestamp 1676037725
transform 1 0 28612 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _621_
timestamp 1676037725
transform 1 0 33120 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _622_
timestamp 1676037725
transform 1 0 31188 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__nor3_1  _623_
timestamp 1676037725
transform 1 0 32568 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _624_
timestamp 1676037725
transform 1 0 41400 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _625_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 41584 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _626_
timestamp 1676037725
transform 1 0 42780 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__nand4_1  _627_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 40020 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _628_
timestamp 1676037725
transform 1 0 40940 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _629_
timestamp 1676037725
transform 1 0 41952 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__a41o_1  _630_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 41216 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _631_
timestamp 1676037725
transform 1 0 40204 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _632_
timestamp 1676037725
transform 1 0 28704 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _633_
timestamp 1676037725
transform 1 0 29716 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _634_
timestamp 1676037725
transform 1 0 13340 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _635_
timestamp 1676037725
transform 1 0 14812 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _636_
timestamp 1676037725
transform 1 0 14260 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _637_
timestamp 1676037725
transform 1 0 14996 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _638_
timestamp 1676037725
transform 1 0 14260 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _639_
timestamp 1676037725
transform 1 0 12420 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _640_
timestamp 1676037725
transform 1 0 5152 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _641_
timestamp 1676037725
transform 1 0 4416 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _642_
timestamp 1676037725
transform 1 0 8004 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _643_
timestamp 1676037725
transform 1 0 8372 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _644_
timestamp 1676037725
transform 1 0 6532 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _645_
timestamp 1676037725
transform 1 0 2668 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _646_
timestamp 1676037725
transform 1 0 12052 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _647_
timestamp 1676037725
transform 1 0 11592 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _648_
timestamp 1676037725
transform 1 0 2668 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _649_
timestamp 1676037725
transform 1 0 2024 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _650_
timestamp 1676037725
transform 1 0 5152 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _651_
timestamp 1676037725
transform 1 0 3220 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _652_
timestamp 1676037725
transform 1 0 9108 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _653_
timestamp 1676037725
transform 1 0 9108 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _654_
timestamp 1676037725
transform 1 0 7820 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _655_
timestamp 1676037725
transform 1 0 11684 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _656_
timestamp 1676037725
transform 1 0 10028 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _657_
timestamp 1676037725
transform 1 0 6900 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _658_
timestamp 1676037725
transform 1 0 2116 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _659_
timestamp 1676037725
transform 1 0 2576 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _660_
timestamp 1676037725
transform 1 0 5152 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _661_
timestamp 1676037725
transform 1 0 3220 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _662_
timestamp 1676037725
transform 1 0 2668 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _663_
timestamp 1676037725
transform 1 0 2024 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _664_
timestamp 1676037725
transform 1 0 17480 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _665_
timestamp 1676037725
transform 1 0 19412 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _666_
timestamp 1676037725
transform 1 0 21988 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _667_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 20516 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_2  _668_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 20884 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _669_
timestamp 1676037725
transform 1 0 21712 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _670_
timestamp 1676037725
transform 1 0 22816 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _671_
timestamp 1676037725
transform 1 0 21988 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _672_
timestamp 1676037725
transform 1 0 20884 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _673_
timestamp 1676037725
transform 1 0 21988 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _674_
timestamp 1676037725
transform 1 0 23368 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _675_
timestamp 1676037725
transform 1 0 14904 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _676_
timestamp 1676037725
transform 1 0 14168 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _677_
timestamp 1676037725
transform 1 0 14260 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _678_
timestamp 1676037725
transform 1 0 15180 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _679_
timestamp 1676037725
transform 1 0 13156 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _680_
timestamp 1676037725
transform 1 0 13984 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _681_
timestamp 1676037725
transform 1 0 12972 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _682_
timestamp 1676037725
transform 1 0 12420 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _683_
timestamp 1676037725
transform 1 0 12144 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _684_
timestamp 1676037725
transform 1 0 14260 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _685_
timestamp 1676037725
transform 1 0 11684 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _686_
timestamp 1676037725
transform 1 0 14812 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _687_
timestamp 1676037725
transform 1 0 14076 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _688_
timestamp 1676037725
transform 1 0 12972 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _689_
timestamp 1676037725
transform 1 0 20976 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _690_
timestamp 1676037725
transform 1 0 20148 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _691_
timestamp 1676037725
transform 1 0 20792 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _692_
timestamp 1676037725
transform 1 0 21436 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _693_
timestamp 1676037725
transform 1 0 40480 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _694_
timestamp 1676037725
transform 1 0 42596 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _695_
timestamp 1676037725
transform 1 0 42596 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _696_
timestamp 1676037725
transform 1 0 42228 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _697_
timestamp 1676037725
transform 1 0 37812 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _698_
timestamp 1676037725
transform 1 0 37628 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _699_
timestamp 1676037725
transform 1 0 33396 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _700_
timestamp 1676037725
transform 1 0 31556 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _701_
timestamp 1676037725
transform 1 0 37444 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _702_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 19412 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  _703_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 30268 0 1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _704_
timestamp 1676037725
transform 1 0 17848 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _705_
timestamp 1676037725
transform 1 0 18492 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _706_
timestamp 1676037725
transform 1 0 19412 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _707_
timestamp 1676037725
transform 1 0 21160 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _708_
timestamp 1676037725
transform 1 0 24564 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _709_
timestamp 1676037725
transform 1 0 18124 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _710_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 32936 0 -1 9792
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _711_
timestamp 1676037725
transform 1 0 17112 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _712_
timestamp 1676037725
transform 1 0 22816 0 -1 10880
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _713_
timestamp 1676037725
transform 1 0 22540 0 -1 9792
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _714_
timestamp 1676037725
transform 1 0 24840 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _715_
timestamp 1676037725
transform 1 0 24564 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfxtp_1  _716_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 25668 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _717_
timestamp 1676037725
transform 1 0 15732 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _718_
timestamp 1676037725
transform 1 0 13156 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _719_
timestamp 1676037725
transform 1 0 9752 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _720_
timestamp 1676037725
transform 1 0 6532 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _721_
timestamp 1676037725
transform 1 0 5428 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _722_
timestamp 1676037725
transform 1 0 4600 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _723_
timestamp 1676037725
transform 1 0 9936 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfrtp_1  _724_
timestamp 1676037725
transform 1 0 24748 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  _725_
timestamp 1676037725
transform 1 0 18216 0 -1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _726_
timestamp 1676037725
transform 1 0 16836 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  _727_
timestamp 1676037725
transform 1 0 17020 0 1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _728_
timestamp 1676037725
transform 1 0 17112 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _729_
timestamp 1676037725
transform 1 0 24564 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _730_
timestamp 1676037725
transform 1 0 16836 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _731_
timestamp 1676037725
transform 1 0 16468 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__conb_1  _732__42 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 15456 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__dfstp_1  _732_
timestamp 1676037725
transform 1 0 14444 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_1  _733_
timestamp 1676037725
transform 1 0 16652 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_1  _734_
timestamp 1676037725
transform 1 0 18492 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__dfxtp_1  _735_
timestamp 1676037725
transform 1 0 27784 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _736_
timestamp 1676037725
transform 1 0 12880 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _737_
timestamp 1676037725
transform 1 0 12328 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _738_
timestamp 1676037725
transform 1 0 13064 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _739_
timestamp 1676037725
transform 1 0 4048 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _740_
timestamp 1676037725
transform 1 0 7176 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _741_
timestamp 1676037725
transform 1 0 3956 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _742_
timestamp 1676037725
transform 1 0 9752 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _743_
timestamp 1676037725
transform 1 0 32292 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _744_
timestamp 1676037725
transform 1 0 34960 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _745_
timestamp 1676037725
transform 1 0 34592 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _746_
timestamp 1676037725
transform 1 0 37444 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _747_
timestamp 1676037725
transform 1 0 28520 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _748_
timestamp 1676037725
transform 1 0 26772 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _749_
timestamp 1676037725
transform 1 0 27140 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _750_
timestamp 1676037725
transform 1 0 28520 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfrtp_1  _751_
timestamp 1676037725
transform 1 0 28428 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfxtp_1  _752_
timestamp 1676037725
transform 1 0 28336 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _753_
timestamp 1676037725
transform 1 0 31280 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _754_
timestamp 1676037725
transform 1 0 32844 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _755_
timestamp 1676037725
transform 1 0 36800 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _756_
timestamp 1676037725
transform 1 0 36892 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _757_
timestamp 1676037725
transform 1 0 37444 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _758_
timestamp 1676037725
transform 1 0 36800 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _759_
timestamp 1676037725
transform 1 0 33948 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _760_
timestamp 1676037725
transform 1 0 29164 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _761_
timestamp 1676037725
transform 1 0 30268 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _762_
timestamp 1676037725
transform 1 0 41400 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _763_
timestamp 1676037725
transform 1 0 40664 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _764_
timestamp 1676037725
transform 1 0 40940 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _765_
timestamp 1676037725
transform 1 0 26128 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _766_
timestamp 1676037725
transform 1 0 11684 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _767_
timestamp 1676037725
transform 1 0 22908 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _768_
timestamp 1676037725
transform 1 0 20332 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _769_
timestamp 1676037725
transform 1 0 29624 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _770_
timestamp 1676037725
transform 1 0 14904 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _771_
timestamp 1676037725
transform 1 0 13156 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _772_
timestamp 1676037725
transform 1 0 10764 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _773_
timestamp 1676037725
transform 1 0 5060 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _774_
timestamp 1676037725
transform 1 0 6900 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _775_
timestamp 1676037725
transform 1 0 3956 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _776_
timestamp 1676037725
transform 1 0 9660 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _777_
timestamp 1676037725
transform 1 0 3312 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _778_
timestamp 1676037725
transform 1 0 4508 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _779_
timestamp 1676037725
transform 1 0 6532 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _780_
timestamp 1676037725
transform 1 0 7176 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _781_
timestamp 1676037725
transform 1 0 9108 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _782_
timestamp 1676037725
transform 1 0 3312 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _783_
timestamp 1676037725
transform 1 0 2024 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _784_
timestamp 1676037725
transform 1 0 3956 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _785_
timestamp 1676037725
transform 1 0 3956 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _786_
timestamp 1676037725
transform 1 0 4140 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _787_
timestamp 1676037725
transform 1 0 8648 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _788_
timestamp 1676037725
transform 1 0 9752 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _789_
timestamp 1676037725
transform 1 0 7912 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _790_
timestamp 1676037725
transform 1 0 3956 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _791_
timestamp 1676037725
transform 1 0 3956 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _792_
timestamp 1676037725
transform 1 0 2116 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfrtp_1  _793_
timestamp 1676037725
transform 1 0 14536 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _794_
timestamp 1676037725
transform 1 0 18124 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _795_
timestamp 1676037725
transform 1 0 20516 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfxtp_2  _796_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 23000 0 -1 5440
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _797_
timestamp 1676037725
transform 1 0 22632 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _798_
timestamp 1676037725
transform 1 0 21528 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _799_
timestamp 1676037725
transform 1 0 13064 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _800_
timestamp 1676037725
transform 1 0 12328 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _801_
timestamp 1676037725
transform 1 0 11776 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _802_
timestamp 1676037725
transform 1 0 12236 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _803_
timestamp 1676037725
transform 1 0 21252 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _804_
timestamp 1676037725
transform 1 0 21988 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _805_
timestamp 1676037725
transform 1 0 31004 0 1 8704
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _806_
timestamp 1676037725
transform 1 0 9844 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _807_
timestamp 1676037725
transform 1 0 11408 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _808_
timestamp 1676037725
transform 1 0 29716 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfrtp_1  _809_
timestamp 1676037725
transform 1 0 40020 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _810_
timestamp 1676037725
transform 1 0 42228 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _811_
timestamp 1676037725
transform 1 0 40296 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _812_
timestamp 1676037725
transform 1 0 40848 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _813_
timestamp 1676037725
transform 1 0 37720 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _814_
timestamp 1676037725
transform 1 0 35420 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _815_
timestamp 1676037725
transform 1 0 31188 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _816_
timestamp 1676037725
transform 1 0 31096 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _817_
timestamp 1676037725
transform 1 0 37444 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_1  _857_
timestamp 1676037725
transform 1 0 42780 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 23092 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_scan_clk_in
timestamp 1676037725
transform 1 0 5612 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_scan_clk_in
timestamp 1676037725
transform 1 0 2576 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_scan_clk_in
timestamp 1676037725
transform 1 0 7820 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_0__f_clk
timestamp 1676037725
transform 1 0 10396 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_1__f_clk
timestamp 1676037725
transform 1 0 15640 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_2__f_clk
timestamp 1676037725
transform 1 0 10396 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_3__f_clk
timestamp 1676037725
transform 1 0 15640 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_4__f_clk
timestamp 1676037725
transform 1 0 28612 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_5__f_clk
timestamp 1676037725
transform 1 0 33764 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_6__f_clk
timestamp 1676037725
transform 1 0 28612 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_7__f_clk
timestamp 1676037725
transform 1 0 33764 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3956 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold2
timestamp 1676037725
transform 1 0 5796 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold3
timestamp 1676037725
transform 1 0 2208 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold4
timestamp 1676037725
transform 1 0 7544 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold5
timestamp 1676037725
transform 1 0 7912 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold6
timestamp 1676037725
transform 1 0 2852 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold7
timestamp 1676037725
transform 1 0 6900 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold8
timestamp 1676037725
transform 1 0 10948 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  input1
timestamp 1676037725
transform 1 0 1564 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1676037725
transform 1 0 43424 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1676037725
transform 1 0 44160 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1676037725
transform 1 0 37444 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1676037725
transform 1 0 31004 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1676037725
transform 1 0 25852 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1676037725
transform 1 0 44160 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input8
timestamp 1676037725
transform 1 0 2300 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input9
timestamp 1676037725
transform 1 0 3128 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input10
timestamp 1676037725
transform 1 0 27140 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input11
timestamp 1676037725
transform 1 0 1564 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input12
timestamp 1676037725
transform 1 0 32292 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input13
timestamp 1676037725
transform 1 0 11684 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input14
timestamp 1676037725
transform 1 0 32292 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input15
timestamp 1676037725
transform 1 0 38732 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input16
timestamp 1676037725
transform 1 0 4600 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input17
timestamp 1676037725
transform 1 0 12880 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input18
timestamp 1676037725
transform 1 0 1564 0 -1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input19
timestamp 1676037725
transform 1 0 42596 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input20
timestamp 1676037725
transform 1 0 44160 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input21
timestamp 1676037725
transform 1 0 1564 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input22
timestamp 1676037725
transform 1 0 24564 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input23
timestamp 1676037725
transform 1 0 34868 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input24
timestamp 1676037725
transform 1 0 17480 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input25
timestamp 1676037725
transform 1 0 16008 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input26
timestamp 1676037725
transform 1 0 9752 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output27
timestamp 1676037725
transform 1 0 44068 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  output28
timestamp 1676037725
transform 1 0 13800 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output29
timestamp 1676037725
transform 1 0 44068 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output30
timestamp 1676037725
transform 1 0 35512 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output31
timestamp 1676037725
transform 1 0 17480 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output32
timestamp 1676037725
transform 1 0 44068 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output33
timestamp 1676037725
transform 1 0 6532 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output34
timestamp 1676037725
transform 1 0 9752 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output35
timestamp 1676037725
transform 1 0 1564 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output36
timestamp 1676037725
transform 1 0 44068 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output37
timestamp 1676037725
transform 1 0 40664 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output38
timestamp 1676037725
transform 1 0 20700 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output39
timestamp 1676037725
transform 1 0 22632 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output40
timestamp 1676037725
transform 1 0 1564 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output41
timestamp 1676037725
transform 1 0 44068 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  scan_controller_43
timestamp 1676037725
transform 1 0 12972 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  scan_controller_44
timestamp 1676037725
transform 1 0 15456 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  scan_controller_45
timestamp 1676037725
transform 1 0 44160 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  scan_controller_46
timestamp 1676037725
transform 1 0 35512 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  scan_controller_47
timestamp 1676037725
transform 1 0 44160 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  scan_controller_48
timestamp 1676037725
transform 1 0 19412 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  scan_controller_49
timestamp 1676037725
transform 1 0 4600 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  scan_controller_50
timestamp 1676037725
transform 1 0 1564 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  scan_controller_51
timestamp 1676037725
transform 1 0 43516 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  scan_controller_52
timestamp 1676037725
transform 1 0 1564 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  scan_controller_53
timestamp 1676037725
transform 1 0 20700 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  scan_controller_54
timestamp 1676037725
transform 1 0 44160 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  scan_controller_55
timestamp 1676037725
transform 1 0 44160 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  scan_controller_56
timestamp 1676037725
transform 1 0 29716 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  scan_controller_57
timestamp 1676037725
transform 1 0 37444 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  scan_controller_58
timestamp 1676037725
transform 1 0 3956 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  scan_controller_59
timestamp 1676037725
transform 1 0 7820 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  scan_controller_60
timestamp 1676037725
transform 1 0 11684 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  scan_controller_61
timestamp 1676037725
transform 1 0 43424 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  scan_controller_62
timestamp 1676037725
transform 1 0 44160 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  scan_controller_63
timestamp 1676037725
transform 1 0 42596 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  scan_controller_64
timestamp 1676037725
transform 1 0 7820 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  scan_controller_65
timestamp 1676037725
transform 1 0 24564 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  scan_controller_66
timestamp 1676037725
transform 1 0 40020 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  scan_controller_67
timestamp 1676037725
transform 1 0 6532 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  scan_controller_68
timestamp 1676037725
transform 1 0 19412 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  scan_controller_69
timestamp 1676037725
transform 1 0 14260 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  scan_controller_70
timestamp 1676037725
transform 1 0 30360 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  scan_controller_71
timestamp 1676037725
transform 1 0 25852 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  scan_controller_72
timestamp 1676037725
transform 1 0 38732 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  scan_controller_73
timestamp 1676037725
transform 1 0 1564 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  scan_controller_74
timestamp 1676037725
transform 1 0 1564 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  scan_controller_75
timestamp 1676037725
transform 1 0 22632 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  scan_controller_76
timestamp 1676037725
transform 1 0 29716 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  scan_controller_77
timestamp 1676037725
transform 1 0 1564 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  scan_controller_78
timestamp 1676037725
transform 1 0 2208 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  scan_controller_79
timestamp 1676037725
transform 1 0 1564 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  scan_controller_80
timestamp 1676037725
transform 1 0 27784 0 -1 17408
box -38 -48 314 592
<< labels >>
flabel metal2 s 1278 19200 1390 20000 0 FreeSans 448 90 0 0 active_select[0]
port 0 nsew signal input
flabel metal2 s 43782 0 43894 800 0 FreeSans 448 90 0 0 active_select[1]
port 1 nsew signal input
flabel metal2 s 45070 0 45182 800 0 FreeSans 448 90 0 0 active_select[2]
port 2 nsew signal input
flabel metal2 s 36698 0 36810 800 0 FreeSans 448 90 0 0 active_select[3]
port 3 nsew signal input
flabel metal2 s 30902 19200 31014 20000 0 FreeSans 448 90 0 0 active_select[4]
port 4 nsew signal input
flabel metal2 s 25750 0 25862 800 0 FreeSans 448 90 0 0 active_select[5]
port 5 nsew signal input
flabel metal3 s 45200 7428 46000 7668 0 FreeSans 960 0 0 0 active_select[6]
port 6 nsew signal input
flabel metal3 s 0 16948 800 17188 0 FreeSans 960 0 0 0 active_select[7]
port 7 nsew signal input
flabel metal2 s 3210 19200 3322 20000 0 FreeSans 448 90 0 0 active_select[8]
port 8 nsew signal input
flabel metal2 s 33478 0 33590 800 0 FreeSans 448 90 0 0 clk
port 9 nsew signal input
flabel metal2 s 27038 0 27150 800 0 FreeSans 448 90 0 0 driver_sel[0]
port 10 nsew signal input
flabel metal2 s -10 19200 102 20000 0 FreeSans 448 90 0 0 driver_sel[1]
port 11 nsew signal input
flabel metal2 s 32190 0 32302 800 0 FreeSans 448 90 0 0 inputs[0]
port 12 nsew signal input
flabel metal2 s 10938 19200 11050 20000 0 FreeSans 448 90 0 0 inputs[1]
port 13 nsew signal input
flabel metal2 s 32190 19200 32302 20000 0 FreeSans 448 90 0 0 inputs[2]
port 14 nsew signal input
flabel metal2 s 38630 19200 38742 20000 0 FreeSans 448 90 0 0 inputs[3]
port 15 nsew signal input
flabel metal2 s 4498 19200 4610 20000 0 FreeSans 448 90 0 0 inputs[4]
port 16 nsew signal input
flabel metal2 s 12870 0 12982 800 0 FreeSans 448 90 0 0 inputs[5]
port 17 nsew signal input
flabel metal3 s 0 4708 800 4948 0 FreeSans 960 0 0 0 inputs[6]
port 18 nsew signal input
flabel metal2 s 41850 0 41962 800 0 FreeSans 448 90 0 0 inputs[7]
port 19 nsew signal input
flabel metal3 s 45200 8788 46000 9028 0 FreeSans 960 0 0 0 la_scan_clk_in
port 20 nsew signal input
flabel metal3 s 0 8108 800 8348 0 FreeSans 960 0 0 0 la_scan_data_in
port 21 nsew signal input
flabel metal3 s 45200 14228 46000 14468 0 FreeSans 960 0 0 0 la_scan_data_out
port 22 nsew signal tristate
flabel metal2 s 23818 19200 23930 20000 0 FreeSans 448 90 0 0 la_scan_latch_en
port 23 nsew signal input
flabel metal2 s 34122 19200 34234 20000 0 FreeSans 448 90 0 0 la_scan_select
port 24 nsew signal input
flabel metal2 s 12870 19200 12982 20000 0 FreeSans 448 90 0 0 oeb[0]
port 25 nsew signal tristate
flabel metal2 s 20598 0 20710 800 0 FreeSans 448 90 0 0 oeb[10]
port 26 nsew signal tristate
flabel metal3 s 45200 12188 46000 12428 0 FreeSans 960 0 0 0 oeb[11]
port 27 nsew signal tristate
flabel metal3 s 45200 15588 46000 15828 0 FreeSans 960 0 0 0 oeb[12]
port 28 nsew signal tristate
flabel metal2 s 28970 0 29082 800 0 FreeSans 448 90 0 0 oeb[13]
port 29 nsew signal tristate
flabel metal2 s 37342 19200 37454 20000 0 FreeSans 448 90 0 0 oeb[14]
port 30 nsew signal tristate
flabel metal2 s 3210 0 3322 800 0 FreeSans 448 90 0 0 oeb[15]
port 31 nsew signal tristate
flabel metal2 s 7718 19200 7830 20000 0 FreeSans 448 90 0 0 oeb[16]
port 32 nsew signal tristate
flabel metal2 s 10938 0 11050 800 0 FreeSans 448 90 0 0 oeb[17]
port 33 nsew signal tristate
flabel metal2 s 43782 19200 43894 20000 0 FreeSans 448 90 0 0 oeb[18]
port 34 nsew signal tristate
flabel metal3 s 45200 10828 46000 11068 0 FreeSans 960 0 0 0 oeb[19]
port 35 nsew signal tristate
flabel metal2 s 16090 0 16202 800 0 FreeSans 448 90 0 0 oeb[1]
port 36 nsew signal tristate
flabel metal2 s 41850 19200 41962 20000 0 FreeSans 448 90 0 0 oeb[20]
port 37 nsew signal tristate
flabel metal2 s 7718 0 7830 800 0 FreeSans 448 90 0 0 oeb[21]
port 38 nsew signal tristate
flabel metal2 s 23818 0 23930 800 0 FreeSans 448 90 0 0 oeb[22]
port 39 nsew signal tristate
flabel metal2 s 39918 0 40030 800 0 FreeSans 448 90 0 0 oeb[23]
port 40 nsew signal tristate
flabel metal2 s 6430 19200 6542 20000 0 FreeSans 448 90 0 0 oeb[24]
port 41 nsew signal tristate
flabel metal2 s 19310 0 19422 800 0 FreeSans 448 90 0 0 oeb[25]
port 42 nsew signal tristate
flabel metal2 s 14158 19200 14270 20000 0 FreeSans 448 90 0 0 oeb[26]
port 43 nsew signal tristate
flabel metal2 s 30258 0 30370 800 0 FreeSans 448 90 0 0 oeb[27]
port 44 nsew signal tristate
flabel metal2 s 25750 19200 25862 20000 0 FreeSans 448 90 0 0 oeb[28]
port 45 nsew signal tristate
flabel metal2 s 38630 0 38742 800 0 FreeSans 448 90 0 0 oeb[29]
port 46 nsew signal tristate
flabel metal3 s 45200 628 46000 868 0 FreeSans 960 0 0 0 oeb[2]
port 47 nsew signal tristate
flabel metal3 s 0 6748 800 6988 0 FreeSans 960 0 0 0 oeb[30]
port 48 nsew signal tristate
flabel metal3 s 0 1308 800 1548 0 FreeSans 960 0 0 0 oeb[31]
port 49 nsew signal tristate
flabel metal2 s 22530 19200 22642 20000 0 FreeSans 448 90 0 0 oeb[32]
port 50 nsew signal tristate
flabel metal2 s 28970 19200 29082 20000 0 FreeSans 448 90 0 0 oeb[33]
port 51 nsew signal tristate
flabel metal3 s 0 3348 800 3588 0 FreeSans 960 0 0 0 oeb[34]
port 52 nsew signal tristate
flabel metal2 s -10 0 102 800 0 FreeSans 448 90 0 0 oeb[35]
port 53 nsew signal tristate
flabel metal3 s 0 18308 800 18548 0 FreeSans 960 0 0 0 oeb[36]
port 54 nsew signal tristate
flabel metal2 s 27682 19200 27794 20000 0 FreeSans 448 90 0 0 oeb[37]
port 55 nsew signal tristate
flabel metal2 s 35410 19200 35522 20000 0 FreeSans 448 90 0 0 oeb[3]
port 56 nsew signal tristate
flabel metal2 s 45070 19200 45182 20000 0 FreeSans 448 90 0 0 oeb[4]
port 57 nsew signal tristate
flabel metal2 s 19310 19200 19422 20000 0 FreeSans 448 90 0 0 oeb[5]
port 58 nsew signal tristate
flabel metal2 s 4498 0 4610 800 0 FreeSans 448 90 0 0 oeb[6]
port 59 nsew signal tristate
flabel metal2 s 1278 0 1390 800 0 FreeSans 448 90 0 0 oeb[7]
port 60 nsew signal tristate
flabel metal3 s 45200 18988 46000 19228 0 FreeSans 960 0 0 0 oeb[8]
port 61 nsew signal tristate
flabel metal3 s 0 13548 800 13788 0 FreeSans 960 0 0 0 oeb[9]
port 62 nsew signal tristate
flabel metal2 s 14158 0 14270 800 0 FreeSans 448 90 0 0 outputs[0]
port 63 nsew signal tristate
flabel metal3 s 45200 17628 46000 17868 0 FreeSans 960 0 0 0 outputs[1]
port 64 nsew signal tristate
flabel metal2 s 35410 0 35522 800 0 FreeSans 448 90 0 0 outputs[2]
port 65 nsew signal tristate
flabel metal2 s 17378 19200 17490 20000 0 FreeSans 448 90 0 0 outputs[3]
port 66 nsew signal tristate
flabel metal3 s 45200 4028 46000 4268 0 FreeSans 960 0 0 0 outputs[4]
port 67 nsew signal tristate
flabel metal2 s 6430 0 6542 800 0 FreeSans 448 90 0 0 outputs[5]
port 68 nsew signal tristate
flabel metal2 s 9650 0 9762 800 0 FreeSans 448 90 0 0 outputs[6]
port 69 nsew signal tristate
flabel metal3 s 0 14908 800 15148 0 FreeSans 960 0 0 0 outputs[7]
port 70 nsew signal tristate
flabel metal3 s 45200 5388 46000 5628 0 FreeSans 960 0 0 0 ready
port 71 nsew signal tristate
flabel metal2 s 17378 0 17490 800 0 FreeSans 448 90 0 0 reset
port 72 nsew signal input
flabel metal3 s 0 11508 800 11748 0 FreeSans 960 0 0 0 scan_clk_in
port 73 nsew signal input
flabel metal2 s 40562 19200 40674 20000 0 FreeSans 448 90 0 0 scan_clk_out
port 74 nsew signal tristate
flabel metal2 s 16090 19200 16202 20000 0 FreeSans 448 90 0 0 scan_data_in
port 75 nsew signal input
flabel metal2 s 20598 19200 20710 20000 0 FreeSans 448 90 0 0 scan_data_out
port 76 nsew signal tristate
flabel metal2 s 22530 0 22642 800 0 FreeSans 448 90 0 0 scan_latch_en
port 77 nsew signal tristate
flabel metal3 s 0 10148 800 10388 0 FreeSans 960 0 0 0 scan_select
port 78 nsew signal tristate
flabel metal2 s 9650 19200 9762 20000 0 FreeSans 448 90 0 0 set_clk_div
port 79 nsew signal input
flabel metal3 s 45200 1988 46000 2228 0 FreeSans 960 0 0 0 slow_clk
port 80 nsew signal tristate
flabel metal4 s 6417 2128 6737 17456 0 FreeSans 1920 90 0 0 vccd1
port 81 nsew power bidirectional
flabel metal4 s 17364 2128 17684 17456 0 FreeSans 1920 90 0 0 vccd1
port 81 nsew power bidirectional
flabel metal4 s 28311 2128 28631 17456 0 FreeSans 1920 90 0 0 vccd1
port 81 nsew power bidirectional
flabel metal4 s 39258 2128 39578 17456 0 FreeSans 1920 90 0 0 vccd1
port 81 nsew power bidirectional
flabel metal4 s 11890 2128 12210 17456 0 FreeSans 1920 90 0 0 vssd1
port 82 nsew ground bidirectional
flabel metal4 s 22837 2128 23157 17456 0 FreeSans 1920 90 0 0 vssd1
port 82 nsew ground bidirectional
flabel metal4 s 33784 2128 34104 17456 0 FreeSans 1920 90 0 0 vssd1
port 82 nsew ground bidirectional
flabel metal4 s 44731 2128 45051 17456 0 FreeSans 1920 90 0 0 vssd1
port 82 nsew ground bidirectional
rlabel metal1 23000 16864 23000 16864 0 vccd1
rlabel via1 23077 17408 23077 17408 0 vssd1
rlabel metal1 26634 13498 26634 13498 0 _000_
rlabel metal1 22754 13974 22754 13974 0 _001_
rlabel metal1 23046 3978 23046 3978 0 _002_
rlabel metal2 14858 4318 14858 4318 0 _003_
rlabel metal1 17434 13192 17434 13192 0 _004_
rlabel metal1 23184 10710 23184 10710 0 _005_
rlabel metal1 24886 13192 24886 13192 0 _006_
rlabel metal1 30774 10778 30774 10778 0 _007_
rlabel metal1 19090 13498 19090 13498 0 _008_
rlabel metal1 19780 12750 19780 12750 0 _009_
rlabel metal1 20700 12274 20700 12274 0 _010_
rlabel metal1 23506 10132 23506 10132 0 _011_
rlabel metal1 24104 12138 24104 12138 0 _012_
rlabel metal2 20102 14484 20102 14484 0 _013_
rlabel metal2 31510 8738 31510 8738 0 _014_
rlabel metal2 20838 10948 20838 10948 0 _015_
rlabel metal2 32430 10914 32430 10914 0 _016_
rlabel metal2 19550 14110 19550 14110 0 _017_
rlabel metal1 18623 12886 18623 12886 0 _018_
rlabel metal1 19320 12070 19320 12070 0 _019_
rlabel metal2 22218 10200 22218 10200 0 _020_
rlabel metal2 25530 11730 25530 11730 0 _021_
rlabel metal1 18860 14518 18860 14518 0 _022_
rlabel metal1 33396 9146 33396 9146 0 _023_
rlabel metal1 17664 14042 17664 14042 0 _024_
rlabel metal2 24702 10472 24702 10472 0 _025_
rlabel metal2 23598 9758 23598 9758 0 _026_
rlabel metal2 26174 11526 26174 11526 0 _027_
rlabel metal1 26503 13226 26503 13226 0 _028_
rlabel metal2 25714 8466 25714 8466 0 _029_
rlabel metal2 19550 9758 19550 9758 0 _030_
rlabel metal1 16238 8296 16238 8296 0 _031_
rlabel metal1 17756 9350 17756 9350 0 _032_
rlabel metal1 17066 7718 17066 7718 0 _033_
rlabel metal1 25668 7174 25668 7174 0 _034_
rlabel metal2 18446 5032 18446 5032 0 _035_
rlabel metal1 18407 5610 18407 5610 0 _036_
rlabel metal2 15870 3502 15870 3502 0 _037_
rlabel metal1 17066 2618 17066 2618 0 _039_
rlabel metal1 18400 3162 18400 3162 0 _041_
rlabel metal1 29164 9078 29164 9078 0 _043_
rlabel metal2 17618 4046 17618 4046 0 _044_
rlabel metal1 19504 4454 19504 4454 0 _045_
rlabel metal2 22126 4318 22126 4318 0 _046_
rlabel metal2 41446 8092 41446 8092 0 _047_
rlabel metal1 42872 7514 42872 7514 0 _048_
rlabel metal1 42281 6358 42281 6358 0 _049_
rlabel metal2 42274 6154 42274 6154 0 _050_
rlabel metal1 38318 5202 38318 5202 0 _051_
rlabel metal1 37359 4522 37359 4522 0 _052_
rlabel metal2 33534 4318 33534 4318 0 _053_
rlabel metal2 31694 3672 31694 3672 0 _054_
rlabel metal1 37904 3706 37904 3706 0 _055_
rlabel metal2 19734 11356 19734 11356 0 _056_
rlabel metal2 26450 9826 26450 9826 0 _057_
rlabel metal1 15686 10778 15686 10778 0 _058_
rlabel metal1 14255 12886 14255 12886 0 _059_
rlabel via1 10069 12818 10069 12818 0 _060_
rlabel metal1 8418 12750 8418 12750 0 _061_
rlabel metal2 6026 11730 6026 11730 0 _062_
rlabel metal1 5055 11730 5055 11730 0 _063_
rlabel via1 10253 11118 10253 11118 0 _064_
rlabel metal2 25070 9180 25070 9180 0 _065_
rlabel metal1 18676 9554 18676 9554 0 _066_
rlabel metal1 16698 8398 16698 8398 0 _067_
rlabel metal1 17204 9010 17204 9010 0 _068_
rlabel metal1 16652 7786 16652 7786 0 _069_
rlabel metal1 24886 6664 24886 6664 0 _070_
rlabel metal1 18124 5134 18124 5134 0 _071_
rlabel metal2 16790 5559 16790 5559 0 _072_
rlabel metal1 32506 7446 32506 7446 0 _073_
rlabel metal1 34714 8874 34714 8874 0 _074_
rlabel metal1 34438 8534 34438 8534 0 _075_
rlabel metal1 37664 8942 37664 8942 0 _076_
rlabel metal1 28750 6970 28750 6970 0 _077_
rlabel metal1 26618 5610 26618 5610 0 _078_
rlabel metal1 27825 4590 27825 4590 0 _079_
rlabel metal1 28412 6358 28412 6358 0 _080_
rlabel metal1 29435 13906 29435 13906 0 _081_
rlabel metal1 31500 14382 31500 14382 0 _082_
rlabel metal1 33299 13906 33299 13906 0 _083_
rlabel metal1 37301 14382 37301 14382 0 _084_
rlabel metal1 37347 13294 37347 13294 0 _085_
rlabel metal1 37664 10642 37664 10642 0 _086_
rlabel metal2 36754 9826 36754 9826 0 _087_
rlabel metal2 35282 11526 35282 11526 0 _088_
rlabel via1 29481 12818 29481 12818 0 _089_
rlabel metal1 32246 11322 32246 11322 0 _090_
rlabel via1 41717 11118 41717 11118 0 _091_
rlabel metal2 41998 14110 41998 14110 0 _092_
rlabel metal1 41160 13294 41160 13294 0 _093_
rlabel metal2 29762 8262 29762 8262 0 _094_
rlabel via1 15221 9622 15221 9622 0 _095_
rlabel metal1 14255 11798 14255 11798 0 _096_
rlabel metal2 12466 12920 12466 12920 0 _097_
rlabel metal1 4906 13226 4906 13226 0 _098_
rlabel metal2 8418 10438 8418 10438 0 _099_
rlabel metal2 4278 9996 4278 9996 0 _100_
rlabel metal2 11638 9350 11638 9350 0 _101_
rlabel metal2 2070 8976 2070 8976 0 _102_
rlabel metal1 4360 11118 4360 11118 0 _103_
rlabel via1 8965 8534 8965 8534 0 _104_
rlabel metal1 10207 8942 10207 8942 0 _105_
rlabel metal1 7574 6358 7574 6358 0 _106_
rlabel metal1 2622 5576 2622 5576 0 _107_
rlabel metal2 3266 6290 3266 6290 0 _108_
rlabel metal1 2336 8466 2336 8466 0 _109_
rlabel metal1 22816 7514 22816 7514 0 _110_
rlabel metal1 23414 7752 23414 7752 0 _111_
rlabel metal1 14301 7446 14301 7446 0 _112_
rlabel metal1 12548 6766 12548 6766 0 _113_
rlabel metal1 11852 4522 11852 4522 0 _114_
rlabel metal2 13110 4726 13110 4726 0 _115_
rlabel metal1 20868 5610 20868 5610 0 _116_
rlabel metal2 21482 6494 21482 6494 0 _117_
rlabel metal1 39560 7242 39560 7242 0 _118_
rlabel metal2 42550 7650 42550 7650 0 _119_
rlabel metal1 40894 5338 40894 5338 0 _120_
rlabel metal1 40756 5066 40756 5066 0 _121_
rlabel metal1 38226 4794 38226 4794 0 _122_
rlabel metal2 35098 4250 35098 4250 0 _123_
rlabel metal2 31510 4828 31510 4828 0 _124_
rlabel metal2 32062 3808 32062 3808 0 _125_
rlabel metal1 36754 4012 36754 4012 0 _126_
rlabel metal1 33488 5542 33488 5542 0 _127_
rlabel metal1 33442 5678 33442 5678 0 _128_
rlabel metal1 33626 6800 33626 6800 0 _129_
rlabel metal1 34132 5882 34132 5882 0 _130_
rlabel metal1 36110 7412 36110 7412 0 _131_
rlabel metal2 38502 6596 38502 6596 0 _132_
rlabel metal2 35282 6970 35282 6970 0 _133_
rlabel metal2 35006 6460 35006 6460 0 _134_
rlabel metal2 35558 7548 35558 7548 0 _135_
rlabel metal1 35190 6324 35190 6324 0 _136_
rlabel metal1 32844 5542 32844 5542 0 _137_
rlabel metal1 33258 6256 33258 6256 0 _138_
rlabel metal1 33074 5882 33074 5882 0 _139_
rlabel metal1 35098 6324 35098 6324 0 _140_
rlabel metal1 34776 5746 34776 5746 0 _141_
rlabel metal2 32890 5678 32890 5678 0 _142_
rlabel metal1 40342 5712 40342 5712 0 _143_
rlabel metal1 40434 6664 40434 6664 0 _144_
rlabel metal1 40296 7174 40296 7174 0 _145_
rlabel metal1 38786 6630 38786 6630 0 _146_
rlabel metal1 39606 5202 39606 5202 0 _147_
rlabel metal1 36110 4998 36110 4998 0 _148_
rlabel metal1 32292 5202 32292 5202 0 _149_
rlabel metal1 32844 4114 32844 4114 0 _150_
rlabel metal1 36583 5338 36583 5338 0 _151_
rlabel metal1 35604 4114 35604 4114 0 _152_
rlabel metal1 38686 5032 38686 5032 0 _153_
rlabel metal1 38929 5338 38929 5338 0 _154_
rlabel metal1 38732 4590 38732 4590 0 _155_
rlabel metal1 40526 5270 40526 5270 0 _156_
rlabel metal2 41078 5372 41078 5372 0 _157_
rlabel metal1 40074 7514 40074 7514 0 _158_
rlabel metal1 41446 7310 41446 7310 0 _159_
rlabel metal2 38778 7582 38778 7582 0 _160_
rlabel metal2 16054 5882 16054 5882 0 _161_
rlabel metal2 19274 5644 19274 5644 0 _162_
rlabel metal1 24472 6426 24472 6426 0 _163_
rlabel metal2 18170 7718 18170 7718 0 _164_
rlabel metal1 17158 9588 17158 9588 0 _165_
rlabel metal2 16882 8228 16882 8228 0 _166_
rlabel metal2 19458 9894 19458 9894 0 _167_
rlabel metal2 25622 9078 25622 9078 0 _168_
rlabel metal1 20424 8534 20424 8534 0 _169_
rlabel metal1 19458 8466 19458 8466 0 _170_
rlabel metal2 20102 7820 20102 7820 0 _171_
rlabel metal1 21114 6154 21114 6154 0 _172_
rlabel metal2 19734 6188 19734 6188 0 _173_
rlabel metal1 20102 6732 20102 6732 0 _174_
rlabel metal1 20240 6630 20240 6630 0 _175_
rlabel metal1 17572 6834 17572 6834 0 _176_
rlabel metal1 20562 6426 20562 6426 0 _177_
rlabel metal1 19734 7956 19734 7956 0 _178_
rlabel metal2 20746 7548 20746 7548 0 _179_
rlabel metal1 20010 7276 20010 7276 0 _180_
rlabel metal1 17894 6630 17894 6630 0 _181_
rlabel metal1 17756 6766 17756 6766 0 _182_
rlabel metal2 18906 7106 18906 7106 0 _183_
rlabel metal1 20240 7514 20240 7514 0 _184_
rlabel metal1 21390 12682 21390 12682 0 _185_
rlabel metal1 19504 11730 19504 11730 0 _186_
rlabel metal1 22402 13362 22402 13362 0 _187_
rlabel metal1 37398 13974 37398 13974 0 _188_
rlabel metal1 39434 11798 39434 11798 0 _189_
rlabel metal2 38134 11968 38134 11968 0 _190_
rlabel metal1 33212 13294 33212 13294 0 _191_
rlabel metal1 39330 11628 39330 11628 0 _192_
rlabel metal1 40250 11696 40250 11696 0 _193_
rlabel metal1 37766 14042 37766 14042 0 _194_
rlabel metal1 38640 13838 38640 13838 0 _195_
rlabel metal1 38456 11118 38456 11118 0 _196_
rlabel metal1 39422 10778 39422 10778 0 _197_
rlabel metal2 38870 11900 38870 11900 0 _198_
rlabel metal1 39514 12750 39514 12750 0 _199_
rlabel metal2 36662 13260 36662 13260 0 _200_
rlabel metal2 36478 12988 36478 12988 0 _201_
rlabel metal1 36386 12410 36386 12410 0 _202_
rlabel metal1 35972 12750 35972 12750 0 _203_
rlabel metal1 32062 13192 32062 13192 0 _204_
rlabel metal1 37122 12614 37122 12614 0 _205_
rlabel metal2 38778 10710 38778 10710 0 _206_
rlabel metal1 35052 10234 35052 10234 0 _207_
rlabel metal1 38364 11050 38364 11050 0 _208_
rlabel metal1 38180 12818 38180 12818 0 _209_
rlabel metal1 24886 12852 24886 12852 0 _210_
rlabel metal2 32798 14042 32798 14042 0 _211_
rlabel metal1 32798 13498 32798 13498 0 _212_
rlabel metal2 32706 12988 32706 12988 0 _213_
rlabel metal1 33948 12818 33948 12818 0 _214_
rlabel metal1 32798 12886 32798 12886 0 _215_
rlabel metal1 33304 12614 33304 12614 0 _216_
rlabel metal2 29762 12036 29762 12036 0 _217_
rlabel metal2 28934 12784 28934 12784 0 _218_
rlabel metal1 22862 11866 22862 11866 0 _219_
rlabel metal1 10994 13362 10994 13362 0 _220_
rlabel metal1 23598 12750 23598 12750 0 _221_
rlabel metal1 25760 10778 25760 10778 0 _222_
rlabel metal1 30360 13226 30360 13226 0 _223_
rlabel metal1 31510 9690 31510 9690 0 _224_
rlabel metal1 15042 5202 15042 5202 0 _225_
rlabel metal2 15226 4794 15226 4794 0 _226_
rlabel metal2 11362 14042 11362 14042 0 _227_
rlabel metal1 9476 3026 9476 3026 0 _228_
rlabel metal2 6854 14960 6854 14960 0 _229_
rlabel metal1 34086 3026 34086 3026 0 _230_
rlabel metal1 15640 10166 15640 10166 0 _231_
rlabel metal2 13570 4624 13570 4624 0 _232_
rlabel metal2 5934 3978 5934 3978 0 _233_
rlabel metal2 7774 4284 7774 4284 0 _234_
rlabel metal2 3450 11764 3450 11764 0 _235_
rlabel metal1 27416 9078 27416 9078 0 _236_
rlabel metal1 27186 13804 27186 13804 0 _237_
rlabel metal1 14122 9146 14122 9146 0 _238_
rlabel metal1 14398 16558 14398 16558 0 _239_
rlabel metal2 25162 14416 25162 14416 0 _240_
rlabel via2 3174 12835 3174 12835 0 _241_
rlabel metal1 22724 14246 22724 14246 0 _242_
rlabel metal1 22310 14246 22310 14246 0 _243_
rlabel metal2 32522 9724 32522 9724 0 _244_
rlabel metal1 23184 13294 23184 13294 0 _245_
rlabel metal2 22678 11322 22678 11322 0 _246_
rlabel metal1 20792 14042 20792 14042 0 _247_
rlabel metal1 26772 12818 26772 12818 0 _248_
rlabel metal1 27278 12954 27278 12954 0 _249_
rlabel metal2 27002 13498 27002 13498 0 _250_
rlabel metal1 22448 12954 22448 12954 0 _251_
rlabel metal1 23092 4114 23092 4114 0 _252_
rlabel metal2 31694 8908 31694 8908 0 _253_
rlabel metal1 33350 4114 33350 4114 0 _254_
rlabel metal1 19090 14382 19090 14382 0 _255_
rlabel metal1 19550 10030 19550 10030 0 _256_
rlabel metal2 29854 9214 29854 9214 0 _257_
rlabel metal1 17020 10778 17020 10778 0 _258_
rlabel metal1 15686 10676 15686 10676 0 _259_
rlabel metal1 14076 12070 14076 12070 0 _260_
rlabel metal1 14536 12818 14536 12818 0 _261_
rlabel metal2 11730 13056 11730 13056 0 _262_
rlabel metal1 10304 13158 10304 13158 0 _263_
rlabel metal2 7406 12784 7406 12784 0 _264_
rlabel metal2 8602 13124 8602 13124 0 _265_
rlabel metal2 7222 11356 7222 11356 0 _266_
rlabel metal1 6486 11118 6486 11118 0 _267_
rlabel metal2 8234 12002 8234 12002 0 _268_
rlabel metal1 4232 11730 4232 11730 0 _269_
rlabel metal1 9982 10778 9982 10778 0 _270_
rlabel metal1 9752 10506 9752 10506 0 _271_
rlabel metal1 22034 4148 22034 4148 0 _272_
rlabel metal1 32522 6970 32522 6970 0 _273_
rlabel metal2 34362 9146 34362 9146 0 _274_
rlabel metal1 34730 8058 34730 8058 0 _275_
rlabel metal1 37628 8602 37628 8602 0 _276_
rlabel metal1 29440 6766 29440 6766 0 _277_
rlabel metal2 26358 5882 26358 5882 0 _278_
rlabel metal2 27462 4828 27462 4828 0 _279_
rlabel metal2 29762 6290 29762 6290 0 _280_
rlabel metal1 30682 13940 30682 13940 0 _281_
rlabel metal2 30866 13702 30866 13702 0 _282_
rlabel via1 31605 14042 31605 14042 0 _283_
rlabel metal2 32522 15164 32522 15164 0 _284_
rlabel metal2 34914 14586 34914 14586 0 _285_
rlabel metal1 34270 14586 34270 14586 0 _286_
rlabel metal2 36662 14416 36662 14416 0 _287_
rlabel metal1 36582 13974 36582 13974 0 _288_
rlabel metal2 36938 14518 36938 14518 0 _289_
rlabel metal1 34132 12886 34132 12886 0 _290_
rlabel metal1 39514 12886 39514 12886 0 _291_
rlabel metal1 37996 12954 37996 12954 0 _292_
rlabel metal1 37398 11118 37398 11118 0 _293_
rlabel metal2 36754 11424 36754 11424 0 _294_
rlabel metal2 36386 10710 36386 10710 0 _295_
rlabel metal1 36432 10778 36432 10778 0 _296_
rlabel metal2 36938 9996 36938 9996 0 _297_
rlabel metal1 35098 11152 35098 11152 0 _298_
rlabel metal1 34516 11798 34516 11798 0 _299_
rlabel metal1 32798 12206 32798 12206 0 _300_
rlabel metal2 29578 12036 29578 12036 0 _301_
rlabel metal1 32223 11254 32223 11254 0 _302_
rlabel via2 31602 12835 31602 12835 0 _303_
rlabel via2 41906 12733 41906 12733 0 _304_
rlabel metal2 41446 12036 41446 12036 0 _305_
rlabel metal1 42780 13498 42780 13498 0 _306_
rlabel metal2 40526 13770 40526 13770 0 _307_
rlabel metal1 41860 14382 41860 14382 0 _308_
rlabel metal1 41170 12954 41170 12954 0 _309_
rlabel metal1 29946 7820 29946 7820 0 _310_
rlabel metal1 13892 10166 13892 10166 0 _311_
rlabel metal2 14674 11526 14674 11526 0 _312_
rlabel metal2 14674 13736 14674 13736 0 _313_
rlabel metal1 4646 13328 4646 13328 0 _314_
rlabel metal1 8510 8058 8510 8058 0 _315_
rlabel metal1 6348 7514 6348 7514 0 _316_
rlabel metal1 12144 8058 12144 8058 0 _317_
rlabel metal2 2254 9724 2254 9724 0 _318_
rlabel metal1 4876 9418 4876 9418 0 _319_
rlabel metal2 9338 9418 9338 9418 0 _320_
rlabel metal1 9292 9146 9292 9146 0 _321_
rlabel metal1 9798 7514 9798 7514 0 _322_
rlabel metal2 2162 6154 2162 6154 0 _323_
rlabel metal1 4324 5678 4324 5678 0 _324_
rlabel metal1 2484 8942 2484 8942 0 _325_
rlabel metal1 21206 11730 21206 11730 0 _326_
rlabel metal1 21528 9078 21528 9078 0 _327_
rlabel metal1 22862 7378 22862 7378 0 _328_
rlabel metal2 22218 7718 22218 7718 0 _329_
rlabel metal2 14950 7888 14950 7888 0 _330_
rlabel metal2 22402 7684 22402 7684 0 _331_
rlabel metal1 13754 6358 13754 6358 0 _332_
rlabel metal2 14674 7616 14674 7616 0 _333_
rlabel metal1 15088 6630 15088 6630 0 _334_
rlabel metal2 13018 6936 13018 6936 0 _335_
rlabel metal1 13386 6120 13386 6120 0 _336_
rlabel metal1 13110 6426 13110 6426 0 _337_
rlabel metal2 12558 5984 12558 5984 0 _338_
rlabel metal2 14490 6290 14490 6290 0 _339_
rlabel metal1 15272 6086 15272 6086 0 _340_
rlabel metal1 13018 4080 13018 4080 0 _341_
rlabel metal1 21482 5338 21482 5338 0 _342_
rlabel metal1 21942 6800 21942 6800 0 _343_
rlabel metal2 32798 9826 32798 9826 0 active
rlabel metal1 1518 17238 1518 17238 0 active_select[0]
rlabel metal2 43838 1588 43838 1588 0 active_select[1]
rlabel metal1 44758 3026 44758 3026 0 active_select[2]
rlabel metal2 36754 840 36754 840 0 active_select[3]
rlabel metal1 31096 17170 31096 17170 0 active_select[4]
rlabel metal2 25806 1588 25806 1588 0 active_select[5]
rlabel via2 44390 7395 44390 7395 0 active_select[6]
rlabel metal3 820 17068 820 17068 0 active_select[7]
rlabel metal2 3266 18234 3266 18234 0 active_select[8]
rlabel metal1 30636 8602 30636 8602 0 aio_input_reg\[0\]
rlabel metal1 16376 9418 16376 9418 0 aio_input_reg\[1\]
rlabel metal1 13984 11866 13984 11866 0 aio_input_reg\[2\]
rlabel metal1 11224 13226 11224 13226 0 aio_input_reg\[3\]
rlabel metal1 6693 13158 6693 13158 0 aio_input_reg\[4\]
rlabel metal2 8326 10914 8326 10914 0 aio_input_reg\[5\]
rlabel metal1 5014 10778 5014 10778 0 aio_input_reg\[6\]
rlabel metal1 11040 9418 11040 9418 0 aio_input_reg\[7\]
rlabel metal1 25576 12818 25576 12818 0 aio_input_sh
rlabel metal1 17434 10540 17434 10540 0 aio_input_shift\[0\]
rlabel metal2 17158 11696 17158 11696 0 aio_input_shift\[1\]
rlabel metal1 13386 12954 13386 12954 0 aio_input_shift\[2\]
rlabel metal1 11638 12818 11638 12818 0 aio_input_shift\[3\]
rlabel metal1 7866 12614 7866 12614 0 aio_input_shift\[4\]
rlabel metal2 7406 11968 7406 11968 0 aio_input_shift\[5\]
rlabel metal1 7314 11730 7314 11730 0 aio_input_shift\[6\]
rlabel metal2 11362 10846 11362 10846 0 aio_input_shift\[7\]
rlabel metal1 29072 7854 29072 7854 0 aio_input_sync\[0\]
rlabel metal2 14306 9860 14306 9860 0 aio_input_sync\[1\]
rlabel metal1 14490 11152 14490 11152 0 aio_input_sync\[2\]
rlabel metal2 14490 13498 14490 13498 0 aio_input_sync\[3\]
rlabel metal1 5428 12954 5428 12954 0 aio_input_sync\[4\]
rlabel metal2 8602 7412 8602 7412 0 aio_input_sync\[5\]
rlabel metal2 5382 6324 5382 6324 0 aio_input_sync\[6\]
rlabel metal2 11178 7106 11178 7106 0 aio_input_sync\[7\]
rlabel metal1 9798 10132 9798 10132 0 aio_output_cap
rlabel metal1 5382 8568 5382 8568 0 aio_output_reg\[0\]
rlabel metal1 6348 13974 6348 13974 0 aio_output_reg\[1\]
rlabel metal2 10074 9248 10074 9248 0 aio_output_reg\[2\]
rlabel metal2 13662 9588 13662 9588 0 aio_output_reg\[3\]
rlabel metal2 9338 6902 9338 6902 0 aio_output_reg\[4\]
rlabel metal1 5336 5882 5336 5882 0 aio_output_reg\[5\]
rlabel metal1 5704 6630 5704 6630 0 aio_output_reg\[6\]
rlabel metal1 3174 8874 3174 8874 0 aio_output_reg\[7\]
rlabel metal1 4728 10030 4728 10030 0 aio_output_shift\[0\]
rlabel metal2 5934 8908 5934 8908 0 aio_output_shift\[1\]
rlabel metal2 7958 10676 7958 10676 0 aio_output_shift\[2\]
rlabel metal1 8004 8398 8004 8398 0 aio_output_shift\[3\]
rlabel metal2 10534 7038 10534 7038 0 aio_output_shift\[4\]
rlabel via1 2341 7786 2341 7786 0 aio_output_shift\[5\]
rlabel metal1 5607 7854 5607 7854 0 aio_output_shift\[6\]
rlabel metal2 5382 8500 5382 8500 0 aio_output_shift\[7\]
rlabel metal1 29854 13702 29854 13702 0 bit_cnt\[0\]
rlabel metal2 32706 14110 32706 14110 0 bit_cnt\[1\]
rlabel metal1 33902 15028 33902 15028 0 bit_cnt\[2\]
rlabel metal1 32752 14314 32752 14314 0 bit_cnt\[3\]
rlabel metal2 33534 2166 33534 2166 0 clk
rlabel metal2 30682 9758 30682 9758 0 clk_divider_I.active
rlabel metal2 31970 7514 31970 7514 0 clk_divider_I.ce
rlabel metal1 33626 7174 33626 7174 0 clk_divider_I.compare\[0\]
rlabel metal2 36386 9350 36386 9350 0 clk_divider_I.compare\[1\]
rlabel metal1 35466 7854 35466 7854 0 clk_divider_I.compare\[2\]
rlabel metal1 37904 8466 37904 8466 0 clk_divider_I.compare\[3\]
rlabel metal1 30360 7514 30360 7514 0 clk_divider_I.compare\[4\]
rlabel metal1 33350 5780 33350 5780 0 clk_divider_I.compare\[5\]
rlabel metal2 33166 5508 33166 5508 0 clk_divider_I.compare\[6\]
rlabel metal1 33488 5610 33488 5610 0 clk_divider_I.compare\[7\]
rlabel metal1 39054 7446 39054 7446 0 clk_divider_I.counter\[0\]
rlabel metal1 39698 7344 39698 7344 0 clk_divider_I.counter\[1\]
rlabel metal1 40066 5712 40066 5712 0 clk_divider_I.counter\[2\]
rlabel metal2 39146 7412 39146 7412 0 clk_divider_I.counter\[3\]
rlabel metal1 34362 6290 34362 6290 0 clk_divider_I.counter\[4\]
rlabel metal1 36984 5610 36984 5610 0 clk_divider_I.counter\[5\]
rlabel metal1 33350 4794 33350 4794 0 clk_divider_I.counter\[6\]
rlabel metal1 32798 4012 32798 4012 0 clk_divider_I.counter\[7\]
rlabel metal2 22126 3298 22126 3298 0 clk_divider_I.reset
rlabel metal1 35650 7922 35650 7922 0 clk_divider_I.set_now
rlabel metal1 11490 13294 11490 13294 0 clk_divider_I.set_sync\[0\]
rlabel metal2 12834 11577 12834 11577 0 clk_divider_I.set_sync\[1\]
rlabel metal2 15686 9282 15686 9282 0 clknet_0_clk
rlabel metal1 6900 8806 6900 8806 0 clknet_0_scan_clk_in
rlabel metal2 3358 9792 3358 9792 0 clknet_1_0__leaf_scan_clk_in
rlabel metal2 7222 9792 7222 9792 0 clknet_1_1__leaf_scan_clk_in
rlabel metal1 2162 8500 2162 8500 0 clknet_3_0__leaf_clk
rlabel metal2 21574 8432 21574 8432 0 clknet_3_1__leaf_clk
rlabel metal1 4048 12818 4048 12818 0 clknet_3_2__leaf_clk
rlabel metal2 18170 14688 18170 14688 0 clknet_3_3__leaf_clk
rlabel metal2 24610 6018 24610 6018 0 clknet_3_4__leaf_clk
rlabel metal2 34638 8704 34638 8704 0 clknet_3_5__leaf_clk
rlabel metal1 26542 14348 26542 14348 0 clknet_3_6__leaf_clk
rlabel metal1 36892 13362 36892 13362 0 clknet_3_7__leaf_clk
rlabel metal2 27094 1588 27094 1588 0 driver_sel[0]
rlabel metal1 874 16558 874 16558 0 driver_sel[1]
rlabel metal2 32246 1588 32246 1588 0 inputs[0]
rlabel metal1 11454 17238 11454 17238 0 inputs[1]
rlabel metal1 32338 17238 32338 17238 0 inputs[2]
rlabel metal1 38778 17238 38778 17238 0 inputs[3]
rlabel metal1 4646 17238 4646 17238 0 inputs[4]
rlabel metal2 12926 1588 12926 1588 0 inputs[5]
rlabel metal3 820 4828 820 4828 0 inputs[6]
rlabel metal2 41906 1554 41906 1554 0 inputs[7]
rlabel metal1 27600 14042 27600 14042 0 int_scan_clk_out
rlabel metal1 13570 10778 13570 10778 0 int_scan_data_out
rlabel metal1 22379 14314 22379 14314 0 int_scan_latch_en
rlabel metal1 24794 13974 24794 13974 0 int_scan_select
rlabel via2 44390 8925 44390 8925 0 la_scan_clk_in
rlabel metal3 820 8228 820 8228 0 la_scan_data_in
rlabel metal2 44298 14297 44298 14297 0 la_scan_data_out
rlabel metal1 24334 17170 24334 17170 0 la_scan_latch_en
rlabel metal2 35098 18122 35098 18122 0 la_scan_select
rlabel metal2 1886 15402 1886 15402 0 net1
rlabel metal1 26588 14926 26588 14926 0 net10
rlabel metal1 1932 16626 1932 16626 0 net11
rlabel metal1 32752 6698 32752 6698 0 net12
rlabel metal1 12558 17034 12558 17034 0 net13
rlabel metal2 32246 14926 32246 14926 0 net14
rlabel metal1 23230 14926 23230 14926 0 net15
rlabel via1 4365 12818 4365 12818 0 net16
rlabel metal1 13018 2482 13018 2482 0 net17
rlabel metal2 18998 5474 18998 5474 0 net18
rlabel metal1 36570 2550 36570 2550 0 net19
rlabel metal1 43148 10030 43148 10030 0 net2
rlabel via2 27738 8891 27738 8891 0 net20
rlabel metal1 13110 7208 13110 7208 0 net21
rlabel metal1 23966 16966 23966 16966 0 net22
rlabel metal2 34914 16048 34914 16048 0 net23
rlabel metal1 16836 2414 16836 2414 0 net24
rlabel metal2 43010 14433 43010 14433 0 net25
rlabel metal1 9890 16966 9890 16966 0 net26
rlabel metal1 44114 14416 44114 14416 0 net27
rlabel metal1 13225 3026 13225 3026 0 net28
rlabel metal1 43562 16218 43562 16218 0 net29
rlabel metal2 38686 10370 38686 10370 0 net3
rlabel metal1 35006 2822 35006 2822 0 net30
rlabel metal1 17066 17170 17066 17170 0 net31
rlabel metal2 44114 4794 44114 4794 0 net32
rlabel metal1 6164 2414 6164 2414 0 net33
rlabel metal1 9706 2414 9706 2414 0 net34
rlabel metal1 2300 15470 2300 15470 0 net35
rlabel metal1 34086 9486 34086 9486 0 net36
rlabel metal2 40710 16796 40710 16796 0 net37
rlabel metal1 17572 16422 17572 16422 0 net38
rlabel metal1 22494 2822 22494 2822 0 net39
rlabel metal1 37812 2618 37812 2618 0 net4
rlabel metal1 2898 12614 2898 12614 0 net40
rlabel metal2 36386 3774 36386 3774 0 net41
rlabel metal2 14858 3264 14858 3264 0 net42
rlabel metal1 13064 17170 13064 17170 0 net43
rlabel metal2 16146 1588 16146 1588 0 net44
rlabel metal3 44996 748 44996 748 0 net45
rlabel metal1 35604 17170 35604 17170 0 net46
rlabel metal1 44758 16762 44758 16762 0 net47
rlabel metal1 19504 17170 19504 17170 0 net48
rlabel metal2 4554 1588 4554 1588 0 net49
rlabel metal1 31004 16966 31004 16966 0 net5
rlabel metal2 1334 1588 1334 1588 0 net50
rlabel metal2 43746 17374 43746 17374 0 net51
rlabel metal3 820 13668 820 13668 0 net52
rlabel metal2 20654 823 20654 823 0 net53
rlabel metal1 44712 12614 44712 12614 0 net54
rlabel metal2 44390 15793 44390 15793 0 net55
rlabel metal2 29026 1588 29026 1588 0 net56
rlabel metal1 37536 17170 37536 17170 0 net57
rlabel metal2 3266 840 3266 840 0 net58
rlabel metal1 7912 17170 7912 17170 0 net59
rlabel metal1 28888 2278 28888 2278 0 net6
rlabel metal2 10994 823 10994 823 0 net60
rlabel metal1 43746 17170 43746 17170 0 net61
rlabel metal1 44712 11118 44712 11118 0 net62
rlabel metal2 42826 18122 42826 18122 0 net63
rlabel metal2 7774 1588 7774 1588 0 net64
rlabel metal2 23874 1588 23874 1588 0 net65
rlabel metal2 39974 823 39974 823 0 net66
rlabel metal1 6624 17170 6624 17170 0 net67
rlabel metal2 19366 1588 19366 1588 0 net68
rlabel metal1 14352 17170 14352 17170 0 net69
rlabel metal1 43608 10574 43608 10574 0 net7
rlabel metal2 30314 823 30314 823 0 net70
rlabel metal1 25944 17170 25944 17170 0 net71
rlabel metal2 38686 1588 38686 1588 0 net72
rlabel metal1 1380 6290 1380 6290 0 net73
rlabel metal3 820 1428 820 1428 0 net74
rlabel metal1 22724 17170 22724 17170 0 net75
rlabel metal1 29486 17170 29486 17170 0 net76
rlabel metal3 820 3468 820 3468 0 net77
rlabel metal2 46 1622 46 1622 0 net78
rlabel metal3 866 18428 866 18428 0 net79
rlabel metal2 2530 16864 2530 16864 0 net8
rlabel metal1 27876 17170 27876 17170 0 net80
rlabel metal2 14490 3196 14490 3196 0 net81
rlabel metal2 16974 3332 16974 3332 0 net82
rlabel metal1 18584 3026 18584 3026 0 net83
rlabel metal1 3910 8806 3910 8806 0 net84
rlabel metal1 6394 8058 6394 8058 0 net85
rlabel metal2 2898 6528 2898 6528 0 net86
rlabel metal2 8234 8772 8234 8772 0 net87
rlabel metal2 9614 10540 9614 10540 0 net88
rlabel metal2 3174 10268 3174 10268 0 net89
rlabel metal1 3772 17034 3772 17034 0 net9
rlabel metal2 5658 7616 5658 7616 0 net90
rlabel metal1 11086 7514 11086 7514 0 net91
rlabel metal1 14030 2822 14030 2822 0 outputs[0]
rlabel metal2 44298 17527 44298 17527 0 outputs[1]
rlabel metal2 35466 1520 35466 1520 0 outputs[2]
rlabel metal1 17572 17306 17572 17306 0 outputs[3]
rlabel metal2 44298 4301 44298 4301 0 outputs[4]
rlabel metal2 6486 1520 6486 1520 0 outputs[5]
rlabel metal2 9706 1520 9706 1520 0 outputs[6]
rlabel metal3 820 15028 820 15028 0 outputs[7]
rlabel metal1 38732 12818 38732 12818 0 proj_cnt\[0\]
rlabel metal2 37766 11968 37766 11968 0 proj_cnt\[1\]
rlabel metal2 36570 11492 36570 11492 0 proj_cnt\[2\]
rlabel metal2 35650 12619 35650 12619 0 proj_cnt\[3\]
rlabel metal1 30820 13294 30820 13294 0 proj_cnt\[4\]
rlabel metal2 31786 10778 31786 10778 0 proj_cnt\[5\]
rlabel metal1 41768 12750 41768 12750 0 proj_cnt\[6\]
rlabel metal2 42090 13328 42090 13328 0 proj_cnt\[7\]
rlabel metal1 41952 12818 41952 12818 0 proj_cnt\[8\]
rlabel metal1 44666 5542 44666 5542 0 ready
rlabel metal2 17434 1588 17434 1588 0 reset
rlabel metal1 16583 3162 16583 3162 0 rst_shift\[0\]
rlabel metal2 18906 3230 18906 3230 0 rst_shift\[1\]
rlabel metal2 4094 11577 4094 11577 0 scan_clk_in
rlabel metal1 40756 17306 40756 17306 0 scan_clk_out
rlabel metal2 16146 18234 16146 18234 0 scan_data_in
rlabel metal1 20838 17306 20838 17306 0 scan_data_out
rlabel metal2 22586 1520 22586 1520 0 scan_latch_en
rlabel metal1 1380 10234 1380 10234 0 scan_select
rlabel metal1 9844 17170 9844 17170 0 set_clk_div
rlabel metal2 44298 2125 44298 2125 0 slow_clk
rlabel metal1 41446 12682 41446 12682 0 state\[0\]
rlabel metal1 26036 12818 26036 12818 0 state\[12\]
rlabel metal1 22448 12614 22448 12614 0 state\[13\]
rlabel metal1 22126 12716 22126 12716 0 state\[1\]
rlabel metal2 20792 13362 20792 13362 0 state\[2\]
rlabel metal1 20976 12410 20976 12410 0 state\[3\]
rlabel metal1 22816 9622 22816 9622 0 state\[4\]
rlabel metal2 25162 11934 25162 11934 0 state\[5\]
rlabel metal2 20470 14382 20470 14382 0 state\[6\]
rlabel metal2 21482 11900 21482 11900 0 state\[8\]
rlabel metal2 20286 13668 20286 13668 0 state\[9\]
rlabel metal2 25990 8704 25990 8704 0 ws_cfg\[0\]
rlabel metal1 20286 8874 20286 8874 0 ws_cfg\[1\]
rlabel metal1 18676 6766 18676 6766 0 ws_cfg\[2\]
rlabel metal1 18653 9146 18653 9146 0 ws_cfg\[3\]
rlabel metal1 19458 7718 19458 7718 0 ws_cfg\[4\]
rlabel metal2 25254 6528 25254 6528 0 ws_cfg\[5\]
rlabel metal1 19918 6358 19918 6358 0 ws_cfg\[6\]
rlabel metal2 18446 6834 18446 6834 0 ws_cfg\[7\]
rlabel metal1 21436 8874 21436 8874 0 ws_cnt\[0\]
rlabel metal2 22034 8092 22034 8092 0 ws_cnt\[1\]
rlabel metal2 14490 7684 14490 7684 0 ws_cnt\[2\]
rlabel metal2 19918 8160 19918 8160 0 ws_cnt\[3\]
rlabel metal1 13754 5678 13754 5678 0 ws_cnt\[4\]
rlabel metal2 19918 6528 19918 6528 0 ws_cnt\[5\]
rlabel metal2 21206 5372 21206 5372 0 ws_cnt\[6\]
rlabel metal1 23046 6426 23046 6426 0 ws_cnt\[7\]
rlabel metal2 19182 6018 19182 6018 0 ws_set_now
rlabel metal1 18354 4046 18354 4046 0 ws_set_sync\[0\]
rlabel metal1 20378 4046 20378 4046 0 ws_set_sync\[1\]
rlabel metal1 22540 4658 22540 4658 0 ws_set_sync\[2\]
<< properties >>
string FIXED_BBOX 0 0 46000 20000
<< end >>
