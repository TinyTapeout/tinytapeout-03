/* Automatically generated from https://wokwi.com/projects/358370685977079809 */

`default_nettype none

module user_module_358370685977079809(
  input [7:0] io_in,
  output [7:0] io_out
);
  wire net1 = io_in[0];
  wire net2 = io_in[1];
  wire net3 = io_in[2];
  wire net4 = io_in[3];
  wire net5 = io_in[4];
  wire net6 = io_in[5];
  wire net7 = io_in[6];
  wire net8 = io_in[7];
  wire net9;
  wire net10;
  wire net11;
  wire net12;
  wire net13;
  wire net14;
  wire net15;
  wire net16;
  wire net17 = 1'b0;
  wire net18 = 1'b1;
  wire net19 = 1'b1;
  wire net20;
  wire net21;
  wire net22;
  wire net23;
  wire net24;
  wire net25;
  wire net26;
  wire net27;
  wire net28;
  wire net29;
  wire net30;
  wire net31;
  wire net32;
  wire net33;
  wire net34;
  wire net35;
  wire net36;
  wire net37;
  wire net38;
  wire net39;
  wire net40;
  wire net41;
  wire net42;
  wire net43;
  wire net44;
  wire net45;
  wire net46;
  wire net47;
  wire net48;
  wire net49;
  wire net50;
  wire net51;
  wire net52;
  wire net53;
  wire net54;
  wire net55;
  wire net56;
  wire net57;
  wire net58;
  wire net59;
  wire net60;
  wire net61;
  wire net62;
  wire net63;
  wire net64;
  wire net65;
  wire net66;
  wire net67;
  wire net68;
  wire net69;
  wire net70;
  wire net71;
  wire net72;
  wire net73;
  wire net74;
  wire net75;
  wire net76;
  wire net77;
  wire net78;
  wire net79;
  wire net80;
  wire net81;
  wire net82;
  wire net83;
  wire net84;
  wire net85;
  wire net86;
  wire net87;
  wire net88;
  wire net89;
  wire net90;
  wire net91;
  wire net92;
  wire net93;
  wire net94;
  wire net95;
  wire net96;
  wire net97;
  wire net98;
  wire net99;
  wire net100;
  wire net101;
  wire net102;
  wire net103;
  wire net104;
  wire net105;
  wire net106;
  wire net107;
  wire net108;
  wire net109;
  wire net110;
  wire net111;
  wire net112;
  wire net113;
  wire net114;
  wire net115;
  wire net116;
  wire net117;
  wire net118;
  wire net119;
  wire net120;
  wire net121;
  wire net122;
  wire net123;
  wire net124;
  wire net125;
  wire net126;
  wire net127;
  wire net128;
  wire net129;
  wire net130;
  wire net131;
  wire net132;
  wire net133;
  wire net134;
  wire net135;
  wire net136;
  wire net137;
  wire net138;
  wire net139;
  wire net140;
  wire net141;
  wire net142;
  wire net143;
  wire net144;
  wire net145;
  wire net146;
  wire net147;
  wire net148;
  wire net149;
  wire net150;
  wire net151;
  wire net152;
  wire net153;
  wire net154;
  wire net155;
  wire net156;
  wire net157;
  wire net158;
  wire net159;
  wire net160;
  wire net161;
  wire net162;
  wire net163;
  wire net164;
  wire net165;
  wire net166;
  wire net167;
  wire net168;
  wire net169;
  wire net170;
  wire net171;
  wire net172;
  wire net173;
  wire net174;
  wire net175;
  wire net176;
  wire net177;
  wire net178;
  wire net179;
  wire net180;
  wire net181;
  wire net182;
  wire net183;
  wire net184;
  wire net185;
  wire net186;
  wire net187;
  wire net188;
  wire net189;
  wire net190;
  wire net191;
  wire net192;
  wire net193;
  wire net194;
  wire net195;
  wire net196;
  wire net197;
  wire net198;
  wire net199;
  wire net200;
  wire net201;
  wire net202;
  wire net203;
  wire net204;
  wire net205 = 1'b0;
  wire net206;
  wire net207;
  wire net208;
  wire net209;
  wire net210;
  wire net211;
  wire net212;
  wire net213;
  wire net214;
  wire net215;
  wire net216;
  wire net217;
  wire net218;
  wire net219;
  wire net220;
  wire net221;
  wire net222;
  wire net223;
  wire net224;
  wire net225;
  wire net226;
  wire net227;
  wire net228;
  wire net229;
  wire net230;
  wire net231;
  wire net232;
  wire net233;
  wire net234;
  wire net235;
  wire net236;
  wire net237;
  wire net238;
  wire net239;
  wire net240;
  wire net241;
  wire net242;
  wire net243;
  wire net244;
  wire net245;
  wire net246;
  wire net247;
  wire net248;
  wire net249;
  wire net250;
  wire net251;
  wire net252;
  wire net253;
  wire net254;
  wire net255;
  wire net256;
  wire net257;
  wire net258;
  wire net259;
  wire net260;
  wire net261;
  wire net262;
  wire net263 = 1'b0;

  assign io_out[0] = net9;
  assign io_out[1] = net10;
  assign io_out[2] = net11;
  assign io_out[3] = net12;
  assign io_out[4] = net13;
  assign io_out[5] = net14;
  assign io_out[6] = net15;
  assign io_out[7] = net16;

  mux_cell mux1 (
    .a (net20),
    .b (net21),
    .sel (net22),
    .out (net9)
  );
  mux_cell mux5 (
    .a (net23),
    .b (net24),
    .sel (net25),
    .out (net20)
  );
  mux_cell mux3 (
    .a (net26),
    .b (net27),
    .sel (net25),
    .out (net28)
  );
  mux_cell mux7 (
    .a (net29),
    .b (net30),
    .sel (net22),
    .out (net11)
  );
  mux_cell mux8 (
    .a (net31),
    .b (net32),
    .sel (net25),
    .out (net29)
  );
  mux_cell mux10 (
    .a (net33),
    .b (net34),
    .sel (net22),
    .out (net12)
  );
  mux_cell mux11 (
    .a (net35),
    .b (net36),
    .sel (net25),
    .out (net33)
  );
  mux_cell mux13 (
    .a (net37),
    .b (net38),
    .sel (net22),
    .out (net13)
  );
  mux_cell mux14 (
    .a (net39),
    .b (net40),
    .sel (net25),
    .out (net37)
  );
  mux_cell mux16 (
    .a (net41),
    .b (net42),
    .sel (net22),
    .out (net14)
  );
  mux_cell mux17 (
    .a (net43),
    .b (net44),
    .sel (net25),
    .out (net41)
  );
  mux_cell mux20 (
    .a (net45),
    .b (net46),
    .sel (net22),
    .out (net15)
  );
  mux_cell mux23 (
    .a (net47),
    .b (net48),
    .sel (net22),
    .out (net16)
  );
  not_cell not1 (
    .in (net49),
    .out (net22)
  );
  not_cell not2 (
    .in (net1),
    .out (net49)
  );
  not_cell not3 (
    .in (net50),
    .out (net25)
  );
  not_cell not4 (
    .in (net2),
    .out (net50)
  );
  dff_cell flop1 (
    .d (net3),
    .clk (net4),
    .q (net51)
  );
  dff_cell flop2 (
    .d (net51),
    .clk (net4),
    .q (net52)
  );
  dff_cell flop3 (
    .d (net52),
    .clk (net4),
    .q (net53)
  );
  dff_cell flop4 (
    .d (net53),
    .clk (net4),
    .q (net54)
  );
  dff_cell flop5 (
    .d (net54),
    .clk (net4),
    .q (net55)
  );
  dff_cell flop6 (
    .d (net55),
    .clk (net4),
    .q (net56)
  );
  dff_cell flop7 (
    .d (net56),
    .clk (net4),
    .q (net57)
  );
  dff_cell flop8 (
    .d (net57),
    .clk (net4),
    .q (net58)
  );
  dff_cell flop9 (
    .d (net51),
    .clk (net5),
    .q (net23)
  );
  dff_cell flop10 (
    .d (net52),
    .clk (net5),
    .q (net26)
  );
  dff_cell flop11 (
    .d (net53),
    .clk (net5),
    .q (net31)
  );
  dff_cell flop12 (
    .d (net54),
    .clk (net5),
    .q (net35)
  );
  dff_cell flop13 (
    .d (net55),
    .clk (net5),
    .q (net39)
  );
  dff_cell flop14 (
    .d (net56),
    .clk (net5),
    .q (net43)
  );
  dff_cell flop15 (
    .d (net57),
    .clk (net5),
    .q (net59)
  );
  dff_cell flop16 (
    .d (net58),
    .clk (net5),
    .q (net60)
  );
  and_cell and4 (
    .a (net61),
    .b (net62),
    .out (net63)
  );
  not_cell not9 (
    .in (net3),
    .out (net61)
  );
  not_cell not10 (
    .in (net4),
    .out (net62)
  );
  and_cell and5 (
    .a (net64),
    .b (net6),
    .out (net65)
  );
  not_cell not11 (
    .in (net5),
    .out (net64)
  );
  and_cell and6 (
    .a (net63),
    .b (net65),
    .out (net66)
  );
  and_cell and7 (
    .a (net67),
    .b (net68),
    .out (net69)
  );
  not_cell not12 (
    .in (net3),
    .out (net67)
  );
  not_cell not13 (
    .in (net4),
    .out (net68)
  );
  and_cell and8 (
    .a (net5),
    .b (net70),
    .out (net71)
  );
  not_cell not15 (
    .in (net6),
    .out (net70)
  );
  and_cell and9 (
    .a (net69),
    .b (net71),
    .out (net72)
  );
  and_cell and10 (
    .a (net73),
    .b (net74),
    .out (net75)
  );
  not_cell not14 (
    .in (net3),
    .out (net73)
  );
  not_cell not16 (
    .in (net4),
    .out (net74)
  );
  and_cell and11 (
    .a (net5),
    .b (net6),
    .out (net76)
  );
  and_cell and12 (
    .a (net75),
    .b (net76),
    .out (net77)
  );
  and_cell and13 (
    .a (net78),
    .b (net4),
    .out (net79)
  );
  not_cell not17 (
    .in (net3),
    .out (net78)
  );
  and_cell and14 (
    .a (net80),
    .b (net81),
    .out (net82)
  );
  not_cell not19 (
    .in (net5),
    .out (net80)
  );
  not_cell not20 (
    .in (net6),
    .out (net81)
  );
  and_cell and15 (
    .a (net79),
    .b (net82),
    .out (net83)
  );
  and_cell and16 (
    .a (net84),
    .b (net4),
    .out (net85)
  );
  not_cell not18 (
    .in (net3),
    .out (net84)
  );
  and_cell and17 (
    .a (net86),
    .b (net6),
    .out (net87)
  );
  not_cell not22 (
    .in (net5),
    .out (net86)
  );
  and_cell and18 (
    .a (net85),
    .b (net87),
    .out (net88)
  );
  and_cell and19 (
    .a (net89),
    .b (net4),
    .out (net90)
  );
  not_cell not21 (
    .in (net3),
    .out (net89)
  );
  and_cell and20 (
    .a (net5),
    .b (net91),
    .out (net92)
  );
  and_cell and21 (
    .a (net90),
    .b (net92),
    .out (net93)
  );
  and_cell and1 (
    .a (net94),
    .b (net95),
    .out (net96)
  );
  not_cell not5 (
    .in (net3),
    .out (net94)
  );
  not_cell not6 (
    .in (net4),
    .out (net95)
  );
  and_cell and2 (
    .a (net97),
    .b (net98),
    .out (net99)
  );
  not_cell not7 (
    .in (net5),
    .out (net97)
  );
  and_cell and3 (
    .a (net96),
    .b (net99),
    .out (net100)
  );
  not_cell not8 (
    .in (net6),
    .out (net98)
  );
  not_cell not24 (
    .in (net6),
    .out (net91)
  );
  and_cell and22 (
    .a (net101),
    .b (net4),
    .out (net102)
  );
  not_cell not23 (
    .in (net3),
    .out (net101)
  );
  and_cell and23 (
    .a (net5),
    .b (net6),
    .out (net103)
  );
  and_cell and24 (
    .a (net102),
    .b (net103),
    .out (net104)
  );
  and_cell and25 (
    .a (net3),
    .b (net105),
    .out (net106)
  );
  not_cell not26 (
    .in (net4),
    .out (net105)
  );
  and_cell and26 (
    .a (net107),
    .b (net108),
    .out (net109)
  );
  not_cell not27 (
    .in (net5),
    .out (net107)
  );
  and_cell and27 (
    .a (net106),
    .b (net109),
    .out (net110)
  );
  not_cell not28 (
    .in (net6),
    .out (net108)
  );
  and_cell and28 (
    .a (net3),
    .b (net111),
    .out (net112)
  );
  not_cell not29 (
    .in (net4),
    .out (net111)
  );
  and_cell and29 (
    .a (net113),
    .b (net6),
    .out (net114)
  );
  not_cell not30 (
    .in (net5),
    .out (net113)
  );
  and_cell and30 (
    .a (net112),
    .b (net114),
    .out (net115)
  );
  and_cell and31 (
    .a (net3),
    .b (net116),
    .out (net117)
  );
  not_cell not31 (
    .in (net4),
    .out (net116)
  );
  and_cell and32 (
    .a (net5),
    .b (net118),
    .out (net119)
  );
  and_cell and33 (
    .a (net117),
    .b (net119),
    .out (net120)
  );
  not_cell not33 (
    .in (net6),
    .out (net118)
  );
  and_cell and34 (
    .a (net3),
    .b (net121),
    .out (net122)
  );
  not_cell not35 (
    .in (net4),
    .out (net121)
  );
  and_cell and35 (
    .a (net5),
    .b (net6),
    .out (net123)
  );
  and_cell and36 (
    .a (net122),
    .b (net123),
    .out (net124)
  );
  and_cell and37 (
    .a (net3),
    .b (net4),
    .out (net125)
  );
  and_cell and38 (
    .a (net126),
    .b (net127),
    .out (net128)
  );
  not_cell not40 (
    .in (net5),
    .out (net126)
  );
  and_cell and39 (
    .a (net125),
    .b (net128),
    .out (net129)
  );
  not_cell not41 (
    .in (net6),
    .out (net127)
  );
  and_cell and40 (
    .a (net3),
    .b (net4),
    .out (net130)
  );
  and_cell and41 (
    .a (net131),
    .b (net6),
    .out (net132)
  );
  not_cell not34 (
    .in (net5),
    .out (net131)
  );
  and_cell and42 (
    .a (net130),
    .b (net132),
    .out (net133)
  );
  and_cell and43 (
    .a (net3),
    .b (net4),
    .out (net134)
  );
  and_cell and44 (
    .a (net5),
    .b (net135),
    .out (net136)
  );
  and_cell and45 (
    .a (net134),
    .b (net136),
    .out (net137)
  );
  not_cell not42 (
    .in (net6),
    .out (net135)
  );
  and_cell and46 (
    .a (net3),
    .b (net4),
    .out (net138)
  );
  and_cell and47 (
    .a (net5),
    .b (net6),
    .out (net139)
  );
  and_cell and48 (
    .a (net138),
    .b (net139),
    .out (net140)
  );
  or_cell or1 (
    .a (net141),
    .b (net142),
    .out (net143)
  );
  or_cell or2 (
    .a (net144),
    .b (net145),
    .out (net141)
  );
  or_cell or3 (
    .a (net146),
    .b (net147),
    .out (net142)
  );
  or_cell or4 (
    .a (net148),
    .b (net149),
    .out (net144)
  );
  or_cell or5 (
    .a (net150),
    .b (net151),
    .out (net145)
  );
  or_cell or6 (
    .a (net124),
    .b (net133),
    .out (net146)
  );
  or_cell or7 (
    .a (net137),
    .b (net140),
    .out (net147)
  );
  or_cell or8 (
    .a (net115),
    .b (net120),
    .out (net151)
  );
  or_cell or9 (
    .a (net93),
    .b (net110),
    .out (net150)
  );
  or_cell or10 (
    .a (net83),
    .b (net88),
    .out (net149)
  );
  or_cell or11 (
    .a (net72),
    .b (net77),
    .out (net148)
  );
  or_cell or12 (
    .a (net152),
    .b (net153),
    .out (net44)
  );
  or_cell or13 (
    .a (net154),
    .b (net155),
    .out (net152)
  );
  or_cell or14 (
    .a (net156),
    .b (net157),
    .out (net153)
  );
  or_cell or15 (
    .a (net158),
    .b (net159),
    .out (net154)
  );
  or_cell or16 (
    .a (net160),
    .b (net120),
    .out (net155)
  );
  or_cell or17 (
    .a (net124),
    .b (net129),
    .out (net156)
  );
  or_cell or18 (
    .a (net137),
    .b (net140),
    .out (net157)
  );
  or_cell or20 (
    .a (net110),
    .b (net115),
    .out (net160)
  );
  or_cell or21 (
    .a (net88),
    .b (net93),
    .out (net159)
  );
  or_cell or22 (
    .a (net100),
    .b (net83),
    .out (net158)
  );
  or_cell or19 (
    .a (net161),
    .b (net162),
    .out (net40)
  );
  or_cell or23 (
    .a (net163),
    .b (net164),
    .out (net161)
  );
  or_cell or24 (
    .a (net165),
    .b (net166),
    .out (net162)
  );
  or_cell or25 (
    .a (net167),
    .b (net168),
    .out (net163)
  );
  or_cell or26 (
    .a (net120),
    .b (net124),
    .out (net164)
  );
  or_cell or27 (
    .a (net129),
    .b (net133),
    .out (net165)
  );
  or_cell or28 (
    .a (net137),
    .b (net140),
    .out (net166)
  );
  or_cell or30 (
    .a (net93),
    .b (net110),
    .out (net168)
  );
  or_cell or31 (
    .a (net100),
    .b (net72),
    .out (net167)
  );
  or_cell or29 (
    .a (net169),
    .b (net170),
    .out (net36)
  );
  or_cell or32 (
    .a (net171),
    .b (net172),
    .out (net169)
  );
  or_cell or33 (
    .a (net173),
    .b (net174),
    .out (net170)
  );
  or_cell or34 (
    .a (net175),
    .b (net176),
    .out (net171)
  );
  or_cell or35 (
    .a (net93),
    .b (net110),
    .out (net172)
  );
  or_cell or36 (
    .a (net124),
    .b (net129),
    .out (net173)
  );
  or_cell or37 (
    .a (net133),
    .b (net137),
    .out (net174)
  );
  or_cell or38 (
    .a (net77),
    .b (net88),
    .out (net176)
  );
  or_cell or39 (
    .a (net100),
    .b (net72),
    .out (net175)
  );
  or_cell or40 (
    .a (net177),
    .b (net178),
    .out (net32)
  );
  or_cell or41 (
    .a (net179),
    .b (net180),
    .out (net177)
  );
  or_cell or42 (
    .a (net181),
    .b (net182),
    .out (net178)
  );
  or_cell or43 (
    .a (net183),
    .b (net184),
    .out (net179)
  );
  or_cell or44 (
    .a (net185),
    .b (net186),
    .out (net180)
  );
  or_cell or45 (
    .a (net115),
    .b (net120),
    .out (net181)
  );
  or_cell or46 (
    .a (net124),
    .b (net133),
    .out (net182)
  );
  or_cell or47 (
    .a (net104),
    .b (net110),
    .out (net186)
  );
  or_cell or48 (
    .a (net88),
    .b (net93),
    .out (net185)
  );
  or_cell or49 (
    .a (net77),
    .b (net83),
    .out (net184)
  );
  or_cell or50 (
    .a (net100),
    .b (net66),
    .out (net183)
  );
  or_cell or52 (
    .a (net187),
    .b (net188),
    .out (net27)
  );
  or_cell or53 (
    .a (net189),
    .b (net190),
    .out (net187)
  );
  or_cell or54 (
    .a (net191),
    .b (net192),
    .out (net188)
  );
  or_cell or55 (
    .a (net193),
    .b (net194),
    .out (net189)
  );
  or_cell or56 (
    .a (net83),
    .b (net104),
    .out (net190)
  );
  or_cell or57 (
    .a (net110),
    .b (net115),
    .out (net191)
  );
  or_cell or58 (
    .a (net120),
    .b (net133),
    .out (net192)
  );
  or_cell or59 (
    .a (net72),
    .b (net77),
    .out (net194)
  );
  or_cell or60 (
    .a (net100),
    .b (net66),
    .out (net193)
  );
  or_cell or61 (
    .a (net195),
    .b (net196),
    .out (net24)
  );
  or_cell or62 (
    .a (net197),
    .b (net198),
    .out (net195)
  );
  or_cell or63 (
    .a (net199),
    .b (net200),
    .out (net196)
  );
  or_cell or64 (
    .a (net201),
    .b (net202),
    .out (net197)
  );
  or_cell or65 (
    .a (net203),
    .b (net204),
    .out (net198)
  );
  or_cell or66 (
    .a (net120),
    .b (net129),
    .out (net199)
  );
  or_cell or67 (
    .a (net137),
    .b (net140),
    .out (net200)
  );
  or_cell or68 (
    .a (net110),
    .b (net115),
    .out (net204)
  );
  or_cell or69 (
    .a (net93),
    .b (net104),
    .out (net203)
  );
  or_cell or70 (
    .a (net77),
    .b (net88),
    .out (net202)
  );
  or_cell or71 (
    .a (net100),
    .b (net72),
    .out (net201)
  );
  mux_cell mux25 (
    .a (net206),
    .b (net207),
    .sel (net8),
    .out (net208)
  );
  mux_cell mux26 (
    .a (net209),
    .b (net210),
    .sel (net7),
    .out (net206)
  );
  mux_cell mux27 (
    .a (net211),
    .b (net212),
    .sel (net7),
    .out (net207)
  );
  xor_cell xor1 (
    .a (net3),
    .b (net4),
    .out (net213)
  );
  and_cell and49 (
    .a (net3),
    .b (net4),
    .out (net214)
  );
  or_cell or51 (
    .a (net3),
    .b (net4),
    .out (net215)
  );
  not_cell not25 (
    .in (net215),
    .out (net216)
  );
  xor_cell xor2 (
    .a (net3),
    .b (net4),
    .out (net217)
  );
  not_cell not32 (
    .in (net217),
    .out (net218)
  );
  or_cell or72 (
    .a (net3),
    .b (net4),
    .out (net219)
  );
  nand_cell nand1 (
    .a (net3),
    .b (net4),
    .out (net220)
  );
  mux_cell mux28 (
    .a (net213),
    .b (net218),
    .sel (net6),
    .out (net212)
  );
  mux_cell mux29 (
    .a (net219),
    .b (net216),
    .sel (net6),
    .out (net211)
  );
  mux_cell mux30 (
    .a (net214),
    .b (net220),
    .sel (net6),
    .out (net210)
  );
  mux_cell mux31 (
    .a (net221),
    .b (net222),
    .sel (net6),
    .out (net209)
  );
  xor_cell xor3 (
    .a (net3),
    .b (net4),
    .out (net223)
  );
  xor_cell xor4 (
    .a (net223),
    .b (net5),
    .out (net221)
  );
  and_cell and50 (
    .a (net5),
    .b (net223),
    .out (net224)
  );
  and_cell and51 (
    .a (net3),
    .b (net4),
    .out (net225)
  );
  or_cell or73 (
    .a (net224),
    .b (net225),
    .out (net222)
  );
  xor_cell xor6 (
    .a (net3),
    .b (net6),
    .out (net226)
  );
  and_cell and52 (
    .a (net3),
    .b (net6),
    .out (net227)
  );
  xor_cell xor7 (
    .a (net4),
    .b (net7),
    .out (net228)
  );
  xor_cell xor8 (
    .a (net228),
    .b (net227),
    .out (net229)
  );
  and_cell and54 (
    .a (net227),
    .b (net228),
    .out (net230)
  );
  and_cell and55 (
    .a (net4),
    .b (net7),
    .out (net231)
  );
  or_cell or75 (
    .a (net230),
    .b (net231),
    .out (net232)
  );
  xor_cell xor9 (
    .a (net5),
    .b (net8),
    .out (net233)
  );
  xor_cell xor10 (
    .a (net233),
    .b (net232),
    .out (net234)
  );
  and_cell and56 (
    .a (net232),
    .b (net233),
    .out (net235)
  );
  and_cell and57 (
    .a (net5),
    .b (net8),
    .out (net236)
  );
  or_cell or76 (
    .a (net235),
    .b (net236),
    .out (net237)
  );
  mux_cell mux2 (
    .a (net229),
    .b (net238),
    .sel (net25),
    .out (net30)
  );
  dffsr_cell flop17 (
    .d (net239),
    .clk (net240),
    .s (net241),
    .r (net242),
    .q (net243)
  );
  dff_cell flop18 (
    .d (net243),
    .clk (net240),
    .q (net244)
  );
  dff_cell flop19 (
    .d (net244),
    .clk (net240),
    .q (net245)
  );
  dff_cell flop20 (
    .d (net245),
    .clk (net240),
    .q (net246)
  );
  dff_cell flop21 (
    .d (net246),
    .clk (net240),
    .q (net247)
  );
  dff_cell flop22 (
    .d (net247),
    .clk (net240),
    .q (net239)
  );
  not_cell not36 (
    .in (net248),
    .out (net240)
  );
  not_cell not37 (
    .in (net5),
    .out (net248)
  );
  not_cell not38 (
    .in (net4),
    .out (net249)
  );
  not_cell not39 (
    .in (net249),
    .out (net242)
  );
  not_cell not43 (
    .in (net3),
    .out (net250)
  );
  not_cell not44 (
    .in (net250),
    .out (net241)
  );
  not_cell not45 (
    .in (net243),
    .out (net251)
  );
  not_cell not46 (
    .in (net251),
    .out (net252)
  );
  not_cell not47 (
    .in (net244),
    .out (net253)
  );
  not_cell not48 (
    .in (net253),
    .out (net254)
  );
  not_cell not49 (
    .in (net245),
    .out (net255)
  );
  not_cell not50 (
    .in (net255),
    .out (net238)
  );
  not_cell not51 (
    .in (net246),
    .out (net256)
  );
  not_cell not52 (
    .in (net256),
    .out (net257)
  );
  not_cell not53 (
    .in (net247),
    .out (net258)
  );
  not_cell not54 (
    .in (net258),
    .out (net259)
  );
  not_cell not55 (
    .in (net239),
    .out (net260)
  );
  not_cell not56 (
    .in (net260),
    .out (net261)
  );
  mux_cell mux4 (
    .a (net208),
    .b (net252),
    .sel (net25),
    .out (net21)
  );
  mux_cell mux6 (
    .a (net28),
    .b (net262),
    .sel (net22),
    .out (net10)
  );
  mux_cell mux9 (
    .a (net234),
    .b (net257),
    .sel (net25),
    .out (net34)
  );
  mux_cell mux12 (
    .a (net237),
    .b (net259),
    .sel (net25),
    .out (net38)
  );
  mux_cell mux18 (
    .a (net226),
    .b (net254),
    .sel (net25),
    .out (net262)
  );
  mux_cell mux15 (
    .a (net263),
    .b (net261),
    .sel (net25),
    .out (net42)
  );
  mux_cell mux19 (
    .a (net59),
    .b (net143),
    .sel (net25),
    .out (net45)
  );
  mux_cell mux21 (
    .a (net263),
    .b (net263),
    .sel (net25),
    .out (net46)
  );
  mux_cell mux22 (
    .a (net60),
    .b (net7),
    .sel (net25),
    .out (net47)
  );
  mux_cell mux24 (
    .a (net263),
    .b (net263),
    .sel (net25),
    .out (net48)
  );
endmodule
