magic
tech sky130A
magscale 1 2
timestamp 1682077834
<< obsli1 >>
rect 1104 1071 4876 22865
<< obsm1 >>
rect 382 1040 5598 22896
<< metal2 >>
rect 386 0 442 800
rect 1122 0 1178 800
rect 1858 0 1914 800
rect 2594 0 2650 800
rect 3330 0 3386 800
rect 4066 0 4122 800
rect 4802 0 4858 800
rect 5538 0 5594 800
<< obsm2 >>
rect 388 856 5594 23225
rect 498 711 1066 856
rect 1234 711 1802 856
rect 1970 711 2538 856
rect 2706 711 3274 856
rect 3442 711 4010 856
rect 4178 711 4746 856
rect 4914 711 5482 856
<< metal3 >>
rect 5200 23128 6000 23248
rect 5200 21632 6000 21752
rect 5200 20136 6000 20256
rect 5200 18640 6000 18760
rect 5200 17144 6000 17264
rect 5200 15648 6000 15768
rect 5200 14152 6000 14272
rect 5200 12656 6000 12776
rect 5200 11160 6000 11280
rect 5200 9664 6000 9784
rect 5200 8168 6000 8288
rect 5200 6672 6000 6792
rect 5200 5176 6000 5296
rect 5200 3680 6000 3800
rect 5200 2184 6000 2304
rect 5200 688 6000 808
<< obsm3 >>
rect 1417 23048 5120 23221
rect 1417 21832 5599 23048
rect 1417 21552 5120 21832
rect 1417 20336 5599 21552
rect 1417 20056 5120 20336
rect 1417 18840 5599 20056
rect 1417 18560 5120 18840
rect 1417 17344 5599 18560
rect 1417 17064 5120 17344
rect 1417 15848 5599 17064
rect 1417 15568 5120 15848
rect 1417 14352 5599 15568
rect 1417 14072 5120 14352
rect 1417 12856 5599 14072
rect 1417 12576 5120 12856
rect 1417 11360 5599 12576
rect 1417 11080 5120 11360
rect 1417 9864 5599 11080
rect 1417 9584 5120 9864
rect 1417 8368 5599 9584
rect 1417 8088 5120 8368
rect 1417 6872 5599 8088
rect 1417 6592 5120 6872
rect 1417 5376 5599 6592
rect 1417 5096 5120 5376
rect 1417 3880 5599 5096
rect 1417 3600 5120 3880
rect 1417 2384 5599 3600
rect 1417 2104 5120 2384
rect 1417 888 5599 2104
rect 1417 715 5120 888
<< metal4 >>
rect 1415 1040 1735 22896
rect 1886 1040 2206 22896
rect 2358 1040 2678 22896
rect 2829 1040 3149 22896
rect 3301 1040 3621 22896
rect 3772 1040 4092 22896
rect 4244 1040 4564 22896
rect 4715 1040 5035 22896
<< labels >>
rlabel metal2 s 386 0 442 800 6 clk_in
port 1 nsew signal input
rlabel metal2 s 5538 0 5594 800 6 clk_out
port 2 nsew signal output
rlabel metal2 s 1122 0 1178 800 6 data_in
port 3 nsew signal input
rlabel metal2 s 4802 0 4858 800 6 data_out
port 4 nsew signal output
rlabel metal2 s 2594 0 2650 800 6 latch_enable_in
port 5 nsew signal input
rlabel metal2 s 3330 0 3386 800 6 latch_enable_out
port 6 nsew signal output
rlabel metal3 s 5200 688 6000 808 6 module_data_in[0]
port 7 nsew signal output
rlabel metal3 s 5200 2184 6000 2304 6 module_data_in[1]
port 8 nsew signal output
rlabel metal3 s 5200 3680 6000 3800 6 module_data_in[2]
port 9 nsew signal output
rlabel metal3 s 5200 5176 6000 5296 6 module_data_in[3]
port 10 nsew signal output
rlabel metal3 s 5200 6672 6000 6792 6 module_data_in[4]
port 11 nsew signal output
rlabel metal3 s 5200 8168 6000 8288 6 module_data_in[5]
port 12 nsew signal output
rlabel metal3 s 5200 9664 6000 9784 6 module_data_in[6]
port 13 nsew signal output
rlabel metal3 s 5200 11160 6000 11280 6 module_data_in[7]
port 14 nsew signal output
rlabel metal3 s 5200 12656 6000 12776 6 module_data_out[0]
port 15 nsew signal input
rlabel metal3 s 5200 14152 6000 14272 6 module_data_out[1]
port 16 nsew signal input
rlabel metal3 s 5200 15648 6000 15768 6 module_data_out[2]
port 17 nsew signal input
rlabel metal3 s 5200 17144 6000 17264 6 module_data_out[3]
port 18 nsew signal input
rlabel metal3 s 5200 18640 6000 18760 6 module_data_out[4]
port 19 nsew signal input
rlabel metal3 s 5200 20136 6000 20256 6 module_data_out[5]
port 20 nsew signal input
rlabel metal3 s 5200 21632 6000 21752 6 module_data_out[6]
port 21 nsew signal input
rlabel metal3 s 5200 23128 6000 23248 6 module_data_out[7]
port 22 nsew signal input
rlabel metal2 s 1858 0 1914 800 6 scan_select_in
port 23 nsew signal input
rlabel metal2 s 4066 0 4122 800 6 scan_select_out
port 24 nsew signal output
rlabel metal4 s 1415 1040 1735 22896 6 vccd1
port 25 nsew power bidirectional
rlabel metal4 s 2358 1040 2678 22896 6 vccd1
port 25 nsew power bidirectional
rlabel metal4 s 3301 1040 3621 22896 6 vccd1
port 25 nsew power bidirectional
rlabel metal4 s 4244 1040 4564 22896 6 vccd1
port 25 nsew power bidirectional
rlabel metal4 s 1886 1040 2206 22896 6 vssd1
port 26 nsew ground bidirectional
rlabel metal4 s 2829 1040 3149 22896 6 vssd1
port 26 nsew ground bidirectional
rlabel metal4 s 3772 1040 4092 22896 6 vssd1
port 26 nsew ground bidirectional
rlabel metal4 s 4715 1040 5035 22896 6 vssd1
port 26 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 6000 24000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 342136
string GDS_FILE /home/matt/work/asic-workshop/shuttle9/tinytapeout-03/openlane/scanchain/runs/23_04_21_13_50/results/signoff/scanchain.magic.gds
string GDS_START 82636
<< end >>

