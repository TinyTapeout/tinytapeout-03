VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO scanchain
  CLASS BLOCK ;
  FOREIGN scanchain ;
  ORIGIN 0.000 0.000 ;
  SIZE 30.000 BY 120.000 ;
  PIN clk_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 6.840 4.000 7.440 ;
    END
  END clk_in
  PIN clk_out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 111.560 4.000 112.160 ;
    END
  END clk_out
  PIN data_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 21.800 4.000 22.400 ;
    END
  END data_in
  PIN data_out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 96.600 4.000 97.200 ;
    END
  END data_out
  PIN latch_enable_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 51.720 4.000 52.320 ;
    END
  END latch_enable_in
  PIN latch_enable_out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 66.680 4.000 67.280 ;
    END
  END latch_enable_out
  PIN module_data_in[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 26.000 3.440 30.000 4.040 ;
    END
  END module_data_in[0]
  PIN module_data_in[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 26.000 10.920 30.000 11.520 ;
    END
  END module_data_in[1]
  PIN module_data_in[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 26.000 18.400 30.000 19.000 ;
    END
  END module_data_in[2]
  PIN module_data_in[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 26.000 25.880 30.000 26.480 ;
    END
  END module_data_in[3]
  PIN module_data_in[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 26.000 33.360 30.000 33.960 ;
    END
  END module_data_in[4]
  PIN module_data_in[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 26.000 40.840 30.000 41.440 ;
    END
  END module_data_in[5]
  PIN module_data_in[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 26.000 48.320 30.000 48.920 ;
    END
  END module_data_in[6]
  PIN module_data_in[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 26.000 55.800 30.000 56.400 ;
    END
  END module_data_in[7]
  PIN module_data_out[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 26.000 63.280 30.000 63.880 ;
    END
  END module_data_out[0]
  PIN module_data_out[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 26.000 70.760 30.000 71.360 ;
    END
  END module_data_out[1]
  PIN module_data_out[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 26.000 78.240 30.000 78.840 ;
    END
  END module_data_out[2]
  PIN module_data_out[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 26.000 85.720 30.000 86.320 ;
    END
  END module_data_out[3]
  PIN module_data_out[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 26.000 93.200 30.000 93.800 ;
    END
  END module_data_out[4]
  PIN module_data_out[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 26.000 100.680 30.000 101.280 ;
    END
  END module_data_out[5]
  PIN module_data_out[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 26.000 108.160 30.000 108.760 ;
    END
  END module_data_out[6]
  PIN module_data_out[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 26.000 115.640 30.000 116.240 ;
    END
  END module_data_out[7]
  PIN scan_select_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 36.760 4.000 37.360 ;
    END
  END scan_select_in
  PIN scan_select_out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 81.640 4.000 82.240 ;
    END
  END scan_select_out
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 7.075 5.200 8.675 114.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 11.790 5.200 13.390 114.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 16.505 5.200 18.105 114.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 21.220 5.200 22.820 114.480 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 9.430 5.200 11.030 114.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 14.145 5.200 15.745 114.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 18.860 5.200 20.460 114.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 23.575 5.200 25.175 114.480 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 5.355 24.380 114.325 ;
      LAYER met1 ;
        RECT 4.670 5.200 27.070 114.480 ;
      LAYER met2 ;
        RECT 4.690 3.555 27.040 116.125 ;
      LAYER met3 ;
        RECT 4.000 115.240 25.600 116.105 ;
        RECT 4.000 112.560 27.290 115.240 ;
        RECT 4.400 111.160 27.290 112.560 ;
        RECT 4.000 109.160 27.290 111.160 ;
        RECT 4.000 107.760 25.600 109.160 ;
        RECT 4.000 101.680 27.290 107.760 ;
        RECT 4.000 100.280 25.600 101.680 ;
        RECT 4.000 97.600 27.290 100.280 ;
        RECT 4.400 96.200 27.290 97.600 ;
        RECT 4.000 94.200 27.290 96.200 ;
        RECT 4.000 92.800 25.600 94.200 ;
        RECT 4.000 86.720 27.290 92.800 ;
        RECT 4.000 85.320 25.600 86.720 ;
        RECT 4.000 82.640 27.290 85.320 ;
        RECT 4.400 81.240 27.290 82.640 ;
        RECT 4.000 79.240 27.290 81.240 ;
        RECT 4.000 77.840 25.600 79.240 ;
        RECT 4.000 71.760 27.290 77.840 ;
        RECT 4.000 70.360 25.600 71.760 ;
        RECT 4.000 67.680 27.290 70.360 ;
        RECT 4.400 66.280 27.290 67.680 ;
        RECT 4.000 64.280 27.290 66.280 ;
        RECT 4.000 62.880 25.600 64.280 ;
        RECT 4.000 56.800 27.290 62.880 ;
        RECT 4.000 55.400 25.600 56.800 ;
        RECT 4.000 52.720 27.290 55.400 ;
        RECT 4.400 51.320 27.290 52.720 ;
        RECT 4.000 49.320 27.290 51.320 ;
        RECT 4.000 47.920 25.600 49.320 ;
        RECT 4.000 41.840 27.290 47.920 ;
        RECT 4.000 40.440 25.600 41.840 ;
        RECT 4.000 37.760 27.290 40.440 ;
        RECT 4.400 36.360 27.290 37.760 ;
        RECT 4.000 34.360 27.290 36.360 ;
        RECT 4.000 32.960 25.600 34.360 ;
        RECT 4.000 26.880 27.290 32.960 ;
        RECT 4.000 25.480 25.600 26.880 ;
        RECT 4.000 22.800 27.290 25.480 ;
        RECT 4.400 21.400 27.290 22.800 ;
        RECT 4.000 19.400 27.290 21.400 ;
        RECT 4.000 18.000 25.600 19.400 ;
        RECT 4.000 11.920 27.290 18.000 ;
        RECT 4.000 10.520 25.600 11.920 ;
        RECT 4.000 7.840 27.290 10.520 ;
        RECT 4.400 6.440 27.290 7.840 ;
        RECT 4.000 4.440 27.290 6.440 ;
        RECT 4.000 3.575 25.600 4.440 ;
  END
END scanchain
END LIBRARY

