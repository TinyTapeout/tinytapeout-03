* NGSPICE file created from user_project_wrapper.ext - technology: sky130A

* Black-box entry subcircuit for psychogenic_neptuneprop abstract view
.subckt psychogenic_neptuneprop io_in[0] io_in[1] io_in[2] io_in[3] io_in[4] io_in[5]
+ io_in[6] io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5] io_out[6]
+ io_out[7] vccd1 vssd1
.ends

* Black-box entry subcircuit for scanchain abstract view
.subckt scanchain clk_in clk_out data_in data_out latch_enable_in latch_enable_out
+ module_data_in[0] module_data_in[1] module_data_in[2] module_data_in[3] module_data_in[4]
+ module_data_in[5] module_data_in[6] module_data_in[7] module_data_out[0] module_data_out[1]
+ module_data_out[2] module_data_out[3] module_data_out[4] module_data_out[5] module_data_out[6]
+ module_data_out[7] scan_select_in scan_select_out vccd1 vssd1
.ends

* Black-box entry subcircuit for top_tt03 abstract view
.subckt top_tt03 io_in[0] io_in[1] io_in[2] io_in[3] io_in[4] io_in[5] io_in[6] io_in[7]
+ io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7]
+ vccd1 vssd1
.ends

* Black-box entry subcircuit for user_module_361728533238569985 abstract view
.subckt user_module_361728533238569985 io_in[0] io_in[1] io_in[2] io_in[3] io_in[4]
+ io_in[5] io_in[6] io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5]
+ io_out[6] io_out[7] vccd1 vssd1
.ends

* Black-box entry subcircuit for diferential_muxpga abstract view
.subckt diferential_muxpga io_in[0] io_in[1] io_in[2] io_in[3] io_in[4] io_in[5] io_in[6]
+ io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7]
+ vccd1 vssd1
.ends

* Black-box entry subcircuit for user_module_360295047631610881 abstract view
.subckt user_module_360295047631610881 io_in[0] io_in[1] io_in[2] io_in[3] io_in[4]
+ io_in[5] io_in[6] io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5]
+ io_out[6] io_out[7] vccd1 vssd1
.ends

* Black-box entry subcircuit for aidan_mcnay_PrimeDetector abstract view
.subckt aidan_mcnay_PrimeDetector io_in[0] io_in[1] io_in[2] io_in[3] io_in[4] io_in[5]
+ io_in[6] io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5] io_out[6]
+ io_out[7] vccd1 vssd1
.ends

* Black-box entry subcircuit for s4ga abstract view
.subckt s4ga io_in[0] io_in[1] io_in[2] io_in[3] io_in[4] io_in[5] io_in[6] io_in[7]
+ io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7]
+ vccd1 vssd1
.ends

* Black-box entry subcircuit for user_module_347140425276981843 abstract view
.subckt user_module_347140425276981843 io_in[0] io_in[1] io_in[2] io_in[3] io_in[4]
+ io_in[5] io_in[6] io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5]
+ io_out[6] io_out[7] vccd1 vssd1
.ends

* Black-box entry subcircuit for user_module_357106633951414273 abstract view
.subckt user_module_357106633951414273 io_in[0] io_in[1] io_in[2] io_in[3] io_in[4]
+ io_in[5] io_in[6] io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5]
+ io_out[6] io_out[7] vccd1 vssd1
.ends

* Black-box entry subcircuit for diferential_rvb3 abstract view
.subckt diferential_rvb3 io_in[0] io_in[1] io_in[2] io_in[3] io_in[4] io_in[5] io_in[6]
+ io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7]
+ vccd1 vssd1
.ends

* Black-box entry subcircuit for kiwih_tt_top abstract view
.subckt kiwih_tt_top io_in[0] io_in[1] io_in[2] io_in[3] io_in[4] io_in[5] io_in[6]
+ io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7]
+ vccd1 vssd1
.ends

* Black-box entry subcircuit for morningjava_top abstract view
.subckt morningjava_top io_in[0] io_in[1] io_in[2] io_in[3] io_in[4] io_in[5] io_in[6]
+ io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7]
+ vccd1 vssd1
.ends

* Black-box entry subcircuit for user_module_357897381919942657 abstract view
.subckt user_module_357897381919942657 io_in[0] io_in[1] io_in[2] io_in[3] io_in[4]
+ io_in[5] io_in[6] io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5]
+ io_out[6] io_out[7] vccd1 vssd1
.ends

* Black-box entry subcircuit for psychogenic_neptunefixed abstract view
.subckt psychogenic_neptunefixed io_in[0] io_in[1] io_in[2] io_in[3] io_in[4] io_in[5]
+ io_in[6] io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5] io_out[6]
+ io_out[7] vccd1 vssd1
.ends

* Black-box entry subcircuit for user_module_354091612057990145 abstract view
.subckt user_module_354091612057990145 io_in[0] io_in[1] io_in[2] io_in[3] io_in[4]
+ io_in[5] io_in[6] io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5]
+ io_out[6] io_out[7] vccd1 vssd1
.ends

* Black-box entry subcircuit for user_module_362371515213982721 abstract view
.subckt user_module_362371515213982721 io_in[0] io_in[1] io_in[2] io_in[3] io_in[4]
+ io_in[5] io_in[6] io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5]
+ io_out[6] io_out[7] vccd1 vssd1
.ends

* Black-box entry subcircuit for user_module_361728681519813633 abstract view
.subckt user_module_361728681519813633 io_in[0] io_in[1] io_in[2] io_in[3] io_in[4]
+ io_in[5] io_in[6] io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5]
+ io_out[6] io_out[7] vccd1 vssd1
.ends

* Black-box entry subcircuit for maheredia_arbiter_game abstract view
.subckt maheredia_arbiter_game io_in[0] io_in[1] io_in[2] io_in[3] io_in[4] io_in[5]
+ io_in[6] io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5] io_out[6]
+ io_out[7] vccd1 vssd1
.ends

* Black-box entry subcircuit for my_design abstract view
.subckt my_design io_in[0] io_in[1] io_in[2] io_in[3] io_in[4] io_in[5] io_in[6] io_in[7]
+ io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7]
+ vccd1 vssd1
.ends

* Black-box entry subcircuit for user_module_360014965627378689 abstract view
.subckt user_module_360014965627378689 io_in[0] io_in[1] io_in[2] io_in[3] io_in[4]
+ io_in[5] io_in[6] io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5]
+ io_out[6] io_out[7] vccd1 vssd1
.ends

* Black-box entry subcircuit for user_module_357917324056483841 abstract view
.subckt user_module_357917324056483841 io_in[0] io_in[1] io_in[2] io_in[3] io_in[4]
+ io_in[5] io_in[6] io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5]
+ io_out[6] io_out[7] vccd1 vssd1
.ends

* Black-box entry subcircuit for moonbase_pdp8 abstract view
.subckt moonbase_pdp8 io_in[0] io_in[1] io_in[2] io_in[3] io_in[4] io_in[5] io_in[6]
+ io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7]
+ vccd1 vssd1
.ends

* Black-box entry subcircuit for user_module_359353377078748161 abstract view
.subckt user_module_359353377078748161 io_in[0] io_in[1] io_in[2] io_in[3] io_in[4]
+ io_in[5] io_in[6] io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5]
+ io_out[6] io_out[7] vccd1 vssd1
.ends

* Black-box entry subcircuit for BenAtUvu_combo abstract view
.subckt BenAtUvu_combo io_in[0] io_in[1] io_in[2] io_in[3] io_in[4] io_in[5] io_in[6]
+ io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7]
+ vccd1 vssd1
.ends

* Black-box entry subcircuit for user_module_359372419264319489 abstract view
.subckt user_module_359372419264319489 io_in[0] io_in[1] io_in[2] io_in[3] io_in[4]
+ io_in[5] io_in[6] io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5]
+ io_out[6] io_out[7] vccd1 vssd1
.ends

* Black-box entry subcircuit for dwisehart_top abstract view
.subckt dwisehart_top io_in[0] io_in[1] io_in[2] io_in[3] io_in[4] io_in[5] io_in[6]
+ io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7]
+ vccd1 vssd1
.ends

* Black-box entry subcircuit for user_module_362336485347742721 abstract view
.subckt user_module_362336485347742721 io_in[0] io_in[1] io_in[2] io_in[3] io_in[4]
+ io_in[5] io_in[6] io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5]
+ io_out[6] io_out[7] vccd1 vssd1
.ends

* Black-box entry subcircuit for kevinwguan_tiny_tapeout abstract view
.subckt kevinwguan_tiny_tapeout io_in[0] io_in[1] io_in[2] io_in[3] io_in[4] io_in[5]
+ io_in[6] io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5] io_out[6]
+ io_out[7] vccd1 vssd1
.ends

* Black-box entry subcircuit for MichaelBell_6bit_fifo abstract view
.subckt MichaelBell_6bit_fifo io_in[0] io_in[1] io_in[2] io_in[3] io_in[4] io_in[5]
+ io_in[6] io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5] io_out[6]
+ io_out[7] vccd1 vssd1
.ends

* Black-box entry subcircuit for jblocklove_cgpt_benchmark_wrapper abstract view
.subckt jblocklove_cgpt_benchmark_wrapper io_in[0] io_in[1] io_in[2] io_in[3] io_in[4]
+ io_in[5] io_in[6] io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5]
+ io_out[6] io_out[7] vccd1 vssd1
.ends

* Black-box entry subcircuit for user_module_347497504164545108 abstract view
.subckt user_module_347497504164545108 io_in[0] io_in[1] io_in[2] io_in[3] io_in[4]
+ io_in[5] io_in[6] io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5]
+ io_out[6] io_out[7] vccd1 vssd1
.ends

* Black-box entry subcircuit for MichaelBell_hovalaag abstract view
.subckt MichaelBell_hovalaag io_in[0] io_in[1] io_in[2] io_in[3] io_in[4] io_in[5]
+ io_in[6] io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5] io_out[6]
+ io_out[7] vccd1 vssd1
.ends

* Black-box entry subcircuit for robbertvanginkel_hamming74 abstract view
.subckt robbertvanginkel_hamming74 io_in[0] io_in[1] io_in[2] io_in[3] io_in[4] io_in[5]
+ io_in[6] io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5] io_out[6]
+ io_out[7] vccd1 vssd1
.ends

* Black-box entry subcircuit for dratini0_fsk_modem_top abstract view
.subckt dratini0_fsk_modem_top io_in[0] io_in[1] io_in[2] io_in[3] io_in[4] io_in[5]
+ io_in[6] io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5] io_out[6]
+ io_out[7] vccd1 vssd1
.ends

* Black-box entry subcircuit for shadow1229_player abstract view
.subckt shadow1229_player io_in[0] io_in[1] io_in[2] io_in[3] io_in[4] io_in[5] io_in[6]
+ io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7]
+ vccd1 vssd1
.ends

* Black-box entry subcircuit for gbsha_ttfir_top abstract view
.subckt gbsha_ttfir_top io_in[0] io_in[1] io_in[2] io_in[3] io_in[4] io_in[5] io_in[6]
+ io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7]
+ vccd1 vssd1
.ends

* Black-box entry subcircuit for diferential_rvb2 abstract view
.subckt diferential_rvb2 io_in[0] io_in[1] io_in[2] io_in[3] io_in[4] io_in[5] io_in[6]
+ io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7]
+ vccd1 vssd1
.ends

* Black-box entry subcircuit for greenstyle_lfsr abstract view
.subckt greenstyle_lfsr io_in[0] io_in[1] io_in[2] io_in[3] io_in[4] io_in[5] io_in[6]
+ io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7]
+ vccd1 vssd1
.ends

* Black-box entry subcircuit for HiddenRoom_HiddenCPU abstract view
.subckt HiddenRoom_HiddenCPU io_in[0] io_in[1] io_in[2] io_in[3] io_in[4] io_in[5]
+ io_in[6] io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5] io_out[6]
+ io_out[7] vccd1 vssd1
.ends

* Black-box entry subcircuit for dratini0_pov_display_top abstract view
.subckt dratini0_pov_display_top io_in[0] io_in[1] io_in[2] io_in[3] io_in[4] io_in[5]
+ io_in[6] io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5] io_out[6]
+ io_out[7] vccd1 vssd1
.ends

* Black-box entry subcircuit for wormy_top abstract view
.subckt wormy_top io_in[0] io_in[1] io_in[2] io_in[3] io_in[4] io_in[5] io_in[6] io_in[7]
+ io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7]
+ vccd1 vssd1
.ends

* Black-box entry subcircuit for bat52_pwm_ddpm_top abstract view
.subckt bat52_pwm_ddpm_top io_in[0] io_in[1] io_in[2] io_in[3] io_in[4] io_in[5] io_in[6]
+ io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7]
+ vccd1 vssd1
.ends

* Black-box entry subcircuit for user_module_340805072482992722 abstract view
.subckt user_module_340805072482992722 io_in[0] io_in[1] io_in[2] io_in[3] io_in[4]
+ io_in[5] io_in[6] io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5]
+ io_out[6] io_out[7] vccd1 vssd1
.ends

* Black-box entry subcircuit for clemensnasenberg_top abstract view
.subckt clemensnasenberg_top io_in[0] io_in[1] io_in[2] io_in[3] io_in[4] io_in[5]
+ io_in[6] io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5] io_out[6]
+ io_out[7] vccd1 vssd1
.ends

* Black-box entry subcircuit for blueintegral_mat_mult abstract view
.subckt blueintegral_mat_mult io_in[0] io_in[1] io_in[2] io_in[3] io_in[4] io_in[5]
+ io_in[6] io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5] io_out[6]
+ io_out[7] vccd1 vssd1
.ends

* Black-box entry subcircuit for wokwi_tt03_simon_top abstract view
.subckt wokwi_tt03_simon_top io_in[0] io_in[1] io_in[2] io_in[3] io_in[4] io_in[5]
+ io_in[6] io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5] io_out[6]
+ io_out[7] vccd1 vssd1
.ends

* Black-box entry subcircuit for user_module_362867354023533569 abstract view
.subckt user_module_362867354023533569 io_in[0] io_in[1] io_in[2] io_in[3] io_in[4]
+ io_in[5] io_in[6] io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5]
+ io_out[6] io_out[7] vccd1 vssd1
.ends

* Black-box entry subcircuit for user_module_362249236392794113 abstract view
.subckt user_module_362249236392794113 io_in[0] io_in[1] io_in[2] io_in[3] io_in[4]
+ io_in[5] io_in[6] io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5]
+ io_out[6] io_out[7] vccd1 vssd1
.ends

* Black-box entry subcircuit for user_module_362441918332875777 abstract view
.subckt user_module_362441918332875777 io_in[0] io_in[1] io_in[2] io_in[3] io_in[4]
+ io_in[5] io_in[6] io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5]
+ io_out[6] io_out[7] vccd1 vssd1
.ends

* Black-box entry subcircuit for htfab_microtapeout abstract view
.subckt htfab_microtapeout io_in[0] io_in[1] io_in[2] io_in[3] io_in[4] io_in[5] io_in[6]
+ io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7]
+ vccd1 vssd1
.ends

* Black-box entry subcircuit for hpretl_tt03_temperature_sensor abstract view
.subckt hpretl_tt03_temperature_sensor io_in[0] io_in[1] io_in[2] io_in[3] io_in[4]
+ io_in[5] io_in[6] io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5]
+ io_out[6] io_out[7] vccd1 vssd1
.ends

* Black-box entry subcircuit for zl_uart abstract view
.subckt zl_uart io_in[0] io_in[1] io_in[2] io_in[3] io_in[4] io_in[5] io_in[6] io_in[7]
+ io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7]
+ vccd1 vssd1
.ends

* Black-box entry subcircuit for tinysat abstract view
.subckt tinysat io_in[0] io_in[1] io_in[2] io_in[3] io_in[4] io_in[5] io_in[6] io_in[7]
+ io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7]
+ vccd1 vssd1
.ends

* Black-box entry subcircuit for dwisehart_ring_top abstract view
.subckt dwisehart_ring_top io_in[0] io_in[1] io_in[2] io_in[3] io_in[4] io_in[5] io_in[6]
+ io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7]
+ vccd1 vssd1
.ends

* Black-box entry subcircuit for jmw95_top abstract view
.subckt jmw95_top io_in[0] io_in[1] io_in[2] io_in[3] io_in[4] io_in[5] io_in[6] io_in[7]
+ io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7]
+ vccd1 vssd1
.ends

* Black-box entry subcircuit for user_module_361684719151591425 abstract view
.subckt user_module_361684719151591425 io_in[0] io_in[1] io_in[2] io_in[3] io_in[4]
+ io_in[5] io_in[6] io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5]
+ io_out[6] io_out[7] vccd1 vssd1
.ends

* Black-box entry subcircuit for dsp_4bits_seq_alu abstract view
.subckt dsp_4bits_seq_alu io_in[0] io_in[1] io_in[2] io_in[3] io_in[4] io_in[5] io_in[6]
+ io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7]
+ vccd1 vssd1
.ends

* Black-box entry subcircuit for guianmonezm_ezmcpu abstract view
.subckt guianmonezm_ezmcpu io_in[0] io_in[1] io_in[2] io_in[3] io_in[4] io_in[5] io_in[6]
+ io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7]
+ vccd1 vssd1
.ends

* Black-box entry subcircuit for lukevassallo_xor_cipher abstract view
.subckt lukevassallo_xor_cipher io_in[0] io_in[1] io_in[2] io_in[3] io_in[4] io_in[5]
+ io_in[6] io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5] io_out[6]
+ io_out[7] vccd1 vssd1
.ends

* Black-box entry subcircuit for user_module_360745091952588801 abstract view
.subckt user_module_360745091952588801 io_in[0] io_in[1] io_in[2] io_in[3] io_in[4]
+ io_in[5] io_in[6] io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5]
+ io_out[6] io_out[7] vccd1 vssd1
.ends

* Black-box entry subcircuit for user_module_358370685977079809 abstract view
.subckt user_module_358370685977079809 io_in[0] io_in[1] io_in[2] io_in[3] io_in[4]
+ io_in[5] io_in[6] io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5]
+ io_out[6] io_out[7] vccd1 vssd1
.ends

* Black-box entry subcircuit for user_module_362675777226104833 abstract view
.subckt user_module_362675777226104833 io_in[0] io_in[1] io_in[2] io_in[3] io_in[4]
+ io_in[5] io_in[6] io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5]
+ io_out[6] io_out[7] vccd1 vssd1
.ends

* Black-box entry subcircuit for meiniki_pi abstract view
.subckt meiniki_pi io_in[0] io_in[1] io_in[2] io_in[3] io_in[4] io_in[5] io_in[6]
+ io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7]
+ vccd1 vssd1
.ends

* Black-box entry subcircuit for user_module_347417602591556180 abstract view
.subckt user_module_347417602591556180 io_in[0] io_in[1] io_in[2] io_in[3] io_in[4]
+ io_in[5] io_in[6] io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5]
+ io_out[6] io_out[7] vccd1 vssd1
.ends

* Black-box entry subcircuit for seven_segment_seconds abstract view
.subckt seven_segment_seconds io_in[0] io_in[1] io_in[2] io_in[3] io_in[4] io_in[5]
+ io_in[6] io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5] io_out[6]
+ io_out[7] vccd1 vssd1
.ends

* Black-box entry subcircuit for tomkeddie_top_tto_a abstract view
.subckt tomkeddie_top_tto_a io_in[0] io_in[1] io_in[2] io_in[3] io_in[4] io_in[5]
+ io_in[6] io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5] io_out[6]
+ io_out[7] vccd1 vssd1
.ends

* Black-box entry subcircuit for diferential_rvb1 abstract view
.subckt diferential_rvb1 io_in[0] io_in[1] io_in[2] io_in[3] io_in[4] io_in[5] io_in[6]
+ io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7]
+ vccd1 vssd1
.ends

* Black-box entry subcircuit for jordan336_toy_cpu abstract view
.subckt jordan336_toy_cpu io_in[0] io_in[1] io_in[2] io_in[3] io_in[4] io_in[5] io_in[6]
+ io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7]
+ vccd1 vssd1
.ends

* Black-box entry subcircuit for knight_rider_KolosKoblasz abstract view
.subckt knight_rider_KolosKoblasz io_in[0] io_in[1] io_in[2] io_in[3] io_in[4] io_in[5]
+ io_in[6] io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5] io_out[6]
+ io_out[7] vccd1 vssd1
.ends

* Black-box entry subcircuit for user_module_357752736742764545 abstract view
.subckt user_module_357752736742764545 io_in[0] io_in[1] io_in[2] io_in[3] io_in[4]
+ io_in[5] io_in[6] io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5]
+ io_out[6] io_out[7] vccd1 vssd1
.ends

* Black-box entry subcircuit for user_module_362208154278843393 abstract view
.subckt user_module_362208154278843393 io_in[0] io_in[1] io_in[2] io_in[3] io_in[4]
+ io_in[5] io_in[6] io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5]
+ io_out[6] io_out[7] vccd1 vssd1
.ends

* Black-box entry subcircuit for user_module_359357227471086593 abstract view
.subckt user_module_359357227471086593 io_in[0] io_in[1] io_in[2] io_in[3] io_in[4]
+ io_in[5] io_in[6] io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5]
+ io_out[6] io_out[7] vccd1 vssd1
.ends

* Black-box entry subcircuit for user_module_362592986761938945 abstract view
.subckt user_module_362592986761938945 io_in[0] io_in[1] io_in[2] io_in[3] io_in[4]
+ io_in[5] io_in[6] io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5]
+ io_out[6] io_out[7] vccd1 vssd1
.ends

* Black-box entry subcircuit for diferential_rvb4 abstract view
.subckt diferential_rvb4 io_in[0] io_in[1] io_in[2] io_in[3] io_in[4] io_in[5] io_in[6]
+ io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7]
+ vccd1 vssd1
.ends

* Black-box entry subcircuit for tiny_bnn abstract view
.subckt tiny_bnn io_in[0] io_in[1] io_in[2] io_in[3] io_in[4] io_in[5] io_in[6] io_in[7]
+ io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7]
+ vccd1 vssd1
.ends

* Black-box entry subcircuit for user_module_358970514554149889 abstract view
.subckt user_module_358970514554149889 io_in[0] io_in[1] io_in[2] io_in[3] io_in[4]
+ io_in[5] io_in[6] io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5]
+ io_out[6] io_out[7] vccd1 vssd1
.ends

* Black-box entry subcircuit for FSM_LAT abstract view
.subckt FSM_LAT io_in[0] io_in[1] io_in[2] io_in[3] io_in[4] io_in[5] io_in[6] io_in[7]
+ io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7]
+ vccd1 vssd1
.ends

* Black-box entry subcircuit for pwm abstract view
.subckt pwm io_in[0] io_in[1] io_in[2] io_in[3] io_in[4] io_in[5] io_in[6] io_in[7]
+ io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7]
+ vccd1 vssd1
.ends

* Black-box entry subcircuit for scan_controller abstract view
.subckt scan_controller active_select[0] active_select[1] active_select[2] active_select[3]
+ active_select[4] active_select[5] active_select[6] active_select[7] active_select[8]
+ clk driver_sel[0] driver_sel[1] inputs[0] inputs[1] inputs[2] inputs[3] inputs[4]
+ inputs[5] inputs[6] inputs[7] la_scan_clk_in la_scan_data_in la_scan_data_out la_scan_latch_en
+ la_scan_select oeb[0] oeb[10] oeb[11] oeb[12] oeb[13] oeb[14] oeb[15] oeb[16] oeb[17]
+ oeb[18] oeb[19] oeb[1] oeb[20] oeb[21] oeb[22] oeb[23] oeb[24] oeb[25] oeb[26] oeb[27]
+ oeb[28] oeb[29] oeb[2] oeb[30] oeb[31] oeb[32] oeb[33] oeb[34] oeb[35] oeb[36] oeb[37]
+ oeb[3] oeb[4] oeb[5] oeb[6] oeb[7] oeb[8] oeb[9] outputs[0] outputs[1] outputs[2]
+ outputs[3] outputs[4] outputs[5] outputs[6] outputs[7] ready reset scan_clk_in scan_clk_out
+ scan_data_in scan_data_out scan_latch_en scan_select set_clk_div slow_clk vccd1
+ vssd1
.ends

* Black-box entry subcircuit for user_module_362379207695863809 abstract view
.subckt user_module_362379207695863809 io_in[0] io_in[1] io_in[2] io_in[3] io_in[4]
+ io_in[5] io_in[6] io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5]
+ io_out[6] io_out[7] vccd1 vssd1
.ends

* Black-box entry subcircuit for user_module_359387860730498049 abstract view
.subckt user_module_359387860730498049 io_in[0] io_in[1] io_in[2] io_in[3] io_in[4]
+ io_in[5] io_in[6] io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5]
+ io_out[6] io_out[7] vccd1 vssd1
.ends

* Black-box entry subcircuit for nikor_clock abstract view
.subckt nikor_clock io_in[0] io_in[1] io_in[2] io_in[3] io_in[4] io_in[5] io_in[6]
+ io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7]
+ vccd1 vssd1
.ends

* Black-box entry subcircuit for granth_crc_decelerator abstract view
.subckt granth_crc_decelerator io_in[0] io_in[1] io_in[2] io_in[3] io_in[4] io_in[5]
+ io_in[6] io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5] io_out[6]
+ io_out[7] vccd1 vssd1
.ends

* Black-box entry subcircuit for user_module_359360834113498113 abstract view
.subckt user_module_359360834113498113 io_in[0] io_in[1] io_in[2] io_in[3] io_in[4]
+ io_in[5] io_in[6] io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5]
+ io_out[6] io_out[7] vccd1 vssd1
.ends

* Black-box entry subcircuit for yannickreiss_dot_op abstract view
.subckt yannickreiss_dot_op io_in[0] io_in[1] io_in[2] io_in[3] io_in[4] io_in[5]
+ io_in[6] io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5] io_out[6]
+ io_out[7] vccd1 vssd1
.ends

* Black-box entry subcircuit for lucaz97_tt_top abstract view
.subckt lucaz97_tt_top io_in[0] io_in[1] io_in[2] io_in[3] io_in[4] io_in[5] io_in[6]
+ io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7]
+ vccd1 vssd1
.ends

* Black-box entry subcircuit for yubex_tiny_logic_analyzer abstract view
.subckt yubex_tiny_logic_analyzer io_in[0] io_in[1] io_in[2] io_in[3] io_in[4] io_in[5]
+ io_in[6] io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5] io_out[6]
+ io_out[7] vccd1 vssd1
.ends

* Black-box entry subcircuit for user_module_339501025136214612 abstract view
.subckt user_module_339501025136214612 io_in[0] io_in[1] io_in[2] io_in[3] io_in[4]
+ io_in[5] io_in[6] io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5]
+ io_out[6] io_out[7] vccd1 vssd1
.ends

* Black-box entry subcircuit for user_module_347144898258928211 abstract view
.subckt user_module_347144898258928211 io_in[0] io_in[1] io_in[2] io_in[3] io_in[4]
+ io_in[5] io_in[6] io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5]
+ io_out[6] io_out[7] vccd1 vssd1
.ends

.subckt user_project_wrapper analog_io[0] analog_io[10] analog_io[11] analog_io[12]
+ analog_io[13] analog_io[14] analog_io[15] analog_io[16] analog_io[17] analog_io[18]
+ analog_io[19] analog_io[1] analog_io[20] analog_io[21] analog_io[22] analog_io[23]
+ analog_io[24] analog_io[25] analog_io[26] analog_io[27] analog_io[28] analog_io[2]
+ analog_io[3] analog_io[4] analog_io[5] analog_io[6] analog_io[7] analog_io[8] analog_io[9]
+ io_in[0] io_in[10] io_in[11] io_in[12] io_in[13] io_in[14] io_in[15] io_in[16] io_in[17]
+ io_in[18] io_in[19] io_in[1] io_in[20] io_in[21] io_in[22] io_in[23] io_in[24] io_in[25]
+ io_in[26] io_in[27] io_in[28] io_in[29] io_in[2] io_in[30] io_in[31] io_in[32] io_in[33]
+ io_in[34] io_in[35] io_in[36] io_in[37] io_in[3] io_in[4] io_in[5] io_in[6] io_in[7]
+ io_in[8] io_in[9] io_oeb[0] io_oeb[10] io_oeb[11] io_oeb[12] io_oeb[13] io_oeb[14]
+ io_oeb[15] io_oeb[16] io_oeb[17] io_oeb[18] io_oeb[19] io_oeb[1] io_oeb[20] io_oeb[21]
+ io_oeb[22] io_oeb[23] io_oeb[24] io_oeb[25] io_oeb[26] io_oeb[27] io_oeb[28] io_oeb[29]
+ io_oeb[2] io_oeb[30] io_oeb[31] io_oeb[32] io_oeb[33] io_oeb[34] io_oeb[35] io_oeb[36]
+ io_oeb[37] io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7] io_oeb[8] io_oeb[9]
+ io_out[0] io_out[10] io_out[11] io_out[12] io_out[13] io_out[14] io_out[15] io_out[16]
+ io_out[17] io_out[18] io_out[19] io_out[1] io_out[20] io_out[21] io_out[22] io_out[23]
+ io_out[24] io_out[25] io_out[26] io_out[27] io_out[28] io_out[29] io_out[2] io_out[30]
+ io_out[31] io_out[32] io_out[33] io_out[34] io_out[35] io_out[36] io_out[37] io_out[3]
+ io_out[4] io_out[5] io_out[6] io_out[7] io_out[8] io_out[9] la_data_in[0] la_data_in[100]
+ la_data_in[101] la_data_in[102] la_data_in[103] la_data_in[104] la_data_in[105]
+ la_data_in[106] la_data_in[107] la_data_in[108] la_data_in[109] la_data_in[10] la_data_in[110]
+ la_data_in[111] la_data_in[112] la_data_in[113] la_data_in[114] la_data_in[115]
+ la_data_in[116] la_data_in[117] la_data_in[118] la_data_in[119] la_data_in[11] la_data_in[120]
+ la_data_in[121] la_data_in[122] la_data_in[123] la_data_in[124] la_data_in[125]
+ la_data_in[126] la_data_in[127] la_data_in[12] la_data_in[13] la_data_in[14] la_data_in[15]
+ la_data_in[16] la_data_in[17] la_data_in[18] la_data_in[19] la_data_in[1] la_data_in[20]
+ la_data_in[21] la_data_in[22] la_data_in[23] la_data_in[24] la_data_in[25] la_data_in[26]
+ la_data_in[27] la_data_in[28] la_data_in[29] la_data_in[2] la_data_in[30] la_data_in[31]
+ la_data_in[32] la_data_in[33] la_data_in[34] la_data_in[35] la_data_in[36] la_data_in[37]
+ la_data_in[38] la_data_in[39] la_data_in[3] la_data_in[40] la_data_in[41] la_data_in[42]
+ la_data_in[43] la_data_in[44] la_data_in[45] la_data_in[46] la_data_in[47] la_data_in[48]
+ la_data_in[49] la_data_in[4] la_data_in[50] la_data_in[51] la_data_in[52] la_data_in[53]
+ la_data_in[54] la_data_in[55] la_data_in[56] la_data_in[57] la_data_in[58] la_data_in[59]
+ la_data_in[5] la_data_in[60] la_data_in[61] la_data_in[62] la_data_in[63] la_data_in[64]
+ la_data_in[65] la_data_in[66] la_data_in[67] la_data_in[68] la_data_in[69] la_data_in[6]
+ la_data_in[70] la_data_in[71] la_data_in[72] la_data_in[73] la_data_in[74] la_data_in[75]
+ la_data_in[76] la_data_in[77] la_data_in[78] la_data_in[79] la_data_in[7] la_data_in[80]
+ la_data_in[81] la_data_in[82] la_data_in[83] la_data_in[84] la_data_in[85] la_data_in[86]
+ la_data_in[87] la_data_in[88] la_data_in[89] la_data_in[8] la_data_in[90] la_data_in[91]
+ la_data_in[92] la_data_in[93] la_data_in[94] la_data_in[95] la_data_in[96] la_data_in[97]
+ la_data_in[98] la_data_in[99] la_data_in[9] la_data_out[0] la_data_out[100] la_data_out[101]
+ la_data_out[102] la_data_out[103] la_data_out[104] la_data_out[105] la_data_out[106]
+ la_data_out[107] la_data_out[108] la_data_out[109] la_data_out[10] la_data_out[110]
+ la_data_out[111] la_data_out[112] la_data_out[113] la_data_out[114] la_data_out[115]
+ la_data_out[116] la_data_out[117] la_data_out[118] la_data_out[119] la_data_out[11]
+ la_data_out[120] la_data_out[121] la_data_out[122] la_data_out[123] la_data_out[124]
+ la_data_out[125] la_data_out[126] la_data_out[127] la_data_out[12] la_data_out[13]
+ la_data_out[14] la_data_out[15] la_data_out[16] la_data_out[17] la_data_out[18]
+ la_data_out[19] la_data_out[1] la_data_out[20] la_data_out[21] la_data_out[22] la_data_out[23]
+ la_data_out[24] la_data_out[25] la_data_out[26] la_data_out[27] la_data_out[28]
+ la_data_out[29] la_data_out[2] la_data_out[30] la_data_out[31] la_data_out[32] la_data_out[33]
+ la_data_out[34] la_data_out[35] la_data_out[36] la_data_out[37] la_data_out[38]
+ la_data_out[39] la_data_out[3] la_data_out[40] la_data_out[41] la_data_out[42] la_data_out[43]
+ la_data_out[44] la_data_out[45] la_data_out[46] la_data_out[47] la_data_out[48]
+ la_data_out[49] la_data_out[4] la_data_out[50] la_data_out[51] la_data_out[52] la_data_out[53]
+ la_data_out[54] la_data_out[55] la_data_out[56] la_data_out[57] la_data_out[58]
+ la_data_out[59] la_data_out[5] la_data_out[60] la_data_out[61] la_data_out[62] la_data_out[63]
+ la_data_out[64] la_data_out[65] la_data_out[66] la_data_out[67] la_data_out[68]
+ la_data_out[69] la_data_out[6] la_data_out[70] la_data_out[71] la_data_out[72] la_data_out[73]
+ la_data_out[74] la_data_out[75] la_data_out[76] la_data_out[77] la_data_out[78]
+ la_data_out[79] la_data_out[7] la_data_out[80] la_data_out[81] la_data_out[82] la_data_out[83]
+ la_data_out[84] la_data_out[85] la_data_out[86] la_data_out[87] la_data_out[88]
+ la_data_out[89] la_data_out[8] la_data_out[90] la_data_out[91] la_data_out[92] la_data_out[93]
+ la_data_out[94] la_data_out[95] la_data_out[96] la_data_out[97] la_data_out[98]
+ la_data_out[99] la_data_out[9] la_oenb[0] la_oenb[100] la_oenb[101] la_oenb[102]
+ la_oenb[103] la_oenb[104] la_oenb[105] la_oenb[106] la_oenb[107] la_oenb[108] la_oenb[109]
+ la_oenb[10] la_oenb[110] la_oenb[111] la_oenb[112] la_oenb[113] la_oenb[114] la_oenb[115]
+ la_oenb[116] la_oenb[117] la_oenb[118] la_oenb[119] la_oenb[11] la_oenb[120] la_oenb[121]
+ la_oenb[122] la_oenb[123] la_oenb[124] la_oenb[125] la_oenb[126] la_oenb[127] la_oenb[12]
+ la_oenb[13] la_oenb[14] la_oenb[15] la_oenb[16] la_oenb[17] la_oenb[18] la_oenb[19]
+ la_oenb[1] la_oenb[20] la_oenb[21] la_oenb[22] la_oenb[23] la_oenb[24] la_oenb[25]
+ la_oenb[26] la_oenb[27] la_oenb[28] la_oenb[29] la_oenb[2] la_oenb[30] la_oenb[31]
+ la_oenb[32] la_oenb[33] la_oenb[34] la_oenb[35] la_oenb[36] la_oenb[37] la_oenb[38]
+ la_oenb[39] la_oenb[3] la_oenb[40] la_oenb[41] la_oenb[42] la_oenb[43] la_oenb[44]
+ la_oenb[45] la_oenb[46] la_oenb[47] la_oenb[48] la_oenb[49] la_oenb[4] la_oenb[50]
+ la_oenb[51] la_oenb[52] la_oenb[53] la_oenb[54] la_oenb[55] la_oenb[56] la_oenb[57]
+ la_oenb[58] la_oenb[59] la_oenb[5] la_oenb[60] la_oenb[61] la_oenb[62] la_oenb[63]
+ la_oenb[64] la_oenb[65] la_oenb[66] la_oenb[67] la_oenb[68] la_oenb[69] la_oenb[6]
+ la_oenb[70] la_oenb[71] la_oenb[72] la_oenb[73] la_oenb[74] la_oenb[75] la_oenb[76]
+ la_oenb[77] la_oenb[78] la_oenb[79] la_oenb[7] la_oenb[80] la_oenb[81] la_oenb[82]
+ la_oenb[83] la_oenb[84] la_oenb[85] la_oenb[86] la_oenb[87] la_oenb[88] la_oenb[89]
+ la_oenb[8] la_oenb[90] la_oenb[91] la_oenb[92] la_oenb[93] la_oenb[94] la_oenb[95]
+ la_oenb[96] la_oenb[97] la_oenb[98] la_oenb[99] la_oenb[9] user_clock2 user_irq[0]
+ user_irq[1] user_irq[2] vccd1 vccd2 vdda1 vdda2 vssa1 vssa2 vssd1 vssd2 wb_clk_i
+ wb_rst_i wbs_ack_o wbs_adr_i[0] wbs_adr_i[10] wbs_adr_i[11] wbs_adr_i[12] wbs_adr_i[13]
+ wbs_adr_i[14] wbs_adr_i[15] wbs_adr_i[16] wbs_adr_i[17] wbs_adr_i[18] wbs_adr_i[19]
+ wbs_adr_i[1] wbs_adr_i[20] wbs_adr_i[21] wbs_adr_i[22] wbs_adr_i[23] wbs_adr_i[24]
+ wbs_adr_i[25] wbs_adr_i[26] wbs_adr_i[27] wbs_adr_i[28] wbs_adr_i[29] wbs_adr_i[2]
+ wbs_adr_i[30] wbs_adr_i[31] wbs_adr_i[3] wbs_adr_i[4] wbs_adr_i[5] wbs_adr_i[6]
+ wbs_adr_i[7] wbs_adr_i[8] wbs_adr_i[9] wbs_cyc_i wbs_dat_i[0] wbs_dat_i[10] wbs_dat_i[11]
+ wbs_dat_i[12] wbs_dat_i[13] wbs_dat_i[14] wbs_dat_i[15] wbs_dat_i[16] wbs_dat_i[17]
+ wbs_dat_i[18] wbs_dat_i[19] wbs_dat_i[1] wbs_dat_i[20] wbs_dat_i[21] wbs_dat_i[22]
+ wbs_dat_i[23] wbs_dat_i[24] wbs_dat_i[25] wbs_dat_i[26] wbs_dat_i[27] wbs_dat_i[28]
+ wbs_dat_i[29] wbs_dat_i[2] wbs_dat_i[30] wbs_dat_i[31] wbs_dat_i[3] wbs_dat_i[4]
+ wbs_dat_i[5] wbs_dat_i[6] wbs_dat_i[7] wbs_dat_i[8] wbs_dat_i[9] wbs_dat_o[0] wbs_dat_o[10]
+ wbs_dat_o[11] wbs_dat_o[12] wbs_dat_o[13] wbs_dat_o[14] wbs_dat_o[15] wbs_dat_o[16]
+ wbs_dat_o[17] wbs_dat_o[18] wbs_dat_o[19] wbs_dat_o[1] wbs_dat_o[20] wbs_dat_o[21]
+ wbs_dat_o[22] wbs_dat_o[23] wbs_dat_o[24] wbs_dat_o[25] wbs_dat_o[26] wbs_dat_o[27]
+ wbs_dat_o[28] wbs_dat_o[29] wbs_dat_o[2] wbs_dat_o[30] wbs_dat_o[31] wbs_dat_o[3]
+ wbs_dat_o[4] wbs_dat_o[5] wbs_dat_o[6] wbs_dat_o[7] wbs_dat_o[8] wbs_dat_o[9] wbs_sel_i[0]
+ wbs_sel_i[1] wbs_sel_i[2] wbs_sel_i[3] wbs_stb_i wbs_we_i
Xpsychogenic_neptuneprop_053 scanchain_053/module_data_in[0] scanchain_053/module_data_in[1]
+ scanchain_053/module_data_in[2] scanchain_053/module_data_in[3] scanchain_053/module_data_in[4]
+ scanchain_053/module_data_in[5] scanchain_053/module_data_in[6] scanchain_053/module_data_in[7]
+ scanchain_053/module_data_out[0] scanchain_053/module_data_out[1] scanchain_053/module_data_out[2]
+ scanchain_053/module_data_out[3] scanchain_053/module_data_out[4] scanchain_053/module_data_out[5]
+ scanchain_053/module_data_out[6] scanchain_053/module_data_out[7] vccd1 vssd1 psychogenic_neptuneprop
Xscanchain_150 scanchain_150/clk_in scanchain_151/clk_in scanchain_150/data_in scanchain_151/data_in
+ scanchain_150/latch_enable_in scanchain_151/latch_enable_in scanchain_150/module_data_in[0]
+ scanchain_150/module_data_in[1] scanchain_150/module_data_in[2] scanchain_150/module_data_in[3]
+ scanchain_150/module_data_in[4] scanchain_150/module_data_in[5] scanchain_150/module_data_in[6]
+ scanchain_150/module_data_in[7] scanchain_150/module_data_out[0] scanchain_150/module_data_out[1]
+ scanchain_150/module_data_out[2] scanchain_150/module_data_out[3] scanchain_150/module_data_out[4]
+ scanchain_150/module_data_out[5] scanchain_150/module_data_out[6] scanchain_150/module_data_out[7]
+ scanchain_150/scan_select_in scanchain_151/scan_select_in vccd1 vssd1 scanchain
Xscanchain_161 scanchain_161/clk_in scanchain_162/clk_in scanchain_161/data_in scanchain_162/data_in
+ scanchain_161/latch_enable_in scanchain_162/latch_enable_in scanchain_161/module_data_in[0]
+ scanchain_161/module_data_in[1] scanchain_161/module_data_in[2] scanchain_161/module_data_in[3]
+ scanchain_161/module_data_in[4] scanchain_161/module_data_in[5] scanchain_161/module_data_in[6]
+ scanchain_161/module_data_in[7] scanchain_161/module_data_out[0] scanchain_161/module_data_out[1]
+ scanchain_161/module_data_out[2] scanchain_161/module_data_out[3] scanchain_161/module_data_out[4]
+ scanchain_161/module_data_out[5] scanchain_161/module_data_out[6] scanchain_161/module_data_out[7]
+ scanchain_161/scan_select_in scanchain_162/scan_select_in vccd1 vssd1 scanchain
Xscanchain_194 scanchain_194/clk_in scanchain_195/clk_in scanchain_194/data_in scanchain_195/data_in
+ scanchain_194/latch_enable_in scanchain_195/latch_enable_in scanchain_194/module_data_in[0]
+ scanchain_194/module_data_in[1] scanchain_194/module_data_in[2] scanchain_194/module_data_in[3]
+ scanchain_194/module_data_in[4] scanchain_194/module_data_in[5] scanchain_194/module_data_in[6]
+ scanchain_194/module_data_in[7] scanchain_194/module_data_out[0] scanchain_194/module_data_out[1]
+ scanchain_194/module_data_out[2] scanchain_194/module_data_out[3] scanchain_194/module_data_out[4]
+ scanchain_194/module_data_out[5] scanchain_194/module_data_out[6] scanchain_194/module_data_out[7]
+ scanchain_194/scan_select_in scanchain_195/scan_select_in vccd1 vssd1 scanchain
Xscanchain_183 scanchain_183/clk_in scanchain_184/clk_in scanchain_183/data_in scanchain_184/data_in
+ scanchain_183/latch_enable_in scanchain_184/latch_enable_in scanchain_183/module_data_in[0]
+ scanchain_183/module_data_in[1] scanchain_183/module_data_in[2] scanchain_183/module_data_in[3]
+ scanchain_183/module_data_in[4] scanchain_183/module_data_in[5] scanchain_183/module_data_in[6]
+ scanchain_183/module_data_in[7] scanchain_183/module_data_out[0] scanchain_183/module_data_out[1]
+ scanchain_183/module_data_out[2] scanchain_183/module_data_out[3] scanchain_183/module_data_out[4]
+ scanchain_183/module_data_out[5] scanchain_183/module_data_out[6] scanchain_183/module_data_out[7]
+ scanchain_183/scan_select_in scanchain_184/scan_select_in vccd1 vssd1 scanchain
Xscanchain_172 scanchain_172/clk_in scanchain_173/clk_in scanchain_172/data_in scanchain_173/data_in
+ scanchain_172/latch_enable_in scanchain_173/latch_enable_in scanchain_172/module_data_in[0]
+ scanchain_172/module_data_in[1] scanchain_172/module_data_in[2] scanchain_172/module_data_in[3]
+ scanchain_172/module_data_in[4] scanchain_172/module_data_in[5] scanchain_172/module_data_in[6]
+ scanchain_172/module_data_in[7] scanchain_172/module_data_out[0] scanchain_172/module_data_out[1]
+ scanchain_172/module_data_out[2] scanchain_172/module_data_out[3] scanchain_172/module_data_out[4]
+ scanchain_172/module_data_out[5] scanchain_172/module_data_out[6] scanchain_172/module_data_out[7]
+ scanchain_172/scan_select_in scanchain_173/scan_select_in vccd1 vssd1 scanchain
Xtop_tt03_059 top_tt03_059/io_in[0] top_tt03_059/io_in[1] top_tt03_059/io_in[2] top_tt03_059/io_in[3]
+ top_tt03_059/io_in[4] top_tt03_059/io_in[5] top_tt03_059/io_in[6] top_tt03_059/io_in[7]
+ top_tt03_059/io_out[0] top_tt03_059/io_out[1] top_tt03_059/io_out[2] top_tt03_059/io_out[3]
+ top_tt03_059/io_out[4] top_tt03_059/io_out[5] top_tt03_059/io_out[6] top_tt03_059/io_out[7]
+ vccd1 vssd1 top_tt03
Xuser_module_361728533238569985_128 scanchain_128/module_data_in[0] scanchain_128/module_data_in[1]
+ scanchain_128/module_data_in[2] scanchain_128/module_data_in[3] scanchain_128/module_data_in[4]
+ scanchain_128/module_data_in[5] scanchain_128/module_data_in[6] scanchain_128/module_data_in[7]
+ scanchain_128/module_data_out[0] scanchain_128/module_data_out[1] scanchain_128/module_data_out[2]
+ scanchain_128/module_data_out[3] scanchain_128/module_data_out[4] scanchain_128/module_data_out[5]
+ scanchain_128/module_data_out[6] scanchain_128/module_data_out[7] vccd1 vssd1 user_module_361728533238569985
Xuser_module_361728533238569985_117 scanchain_117/module_data_in[0] scanchain_117/module_data_in[1]
+ scanchain_117/module_data_in[2] scanchain_117/module_data_in[3] scanchain_117/module_data_in[4]
+ scanchain_117/module_data_in[5] scanchain_117/module_data_in[6] scanchain_117/module_data_in[7]
+ scanchain_117/module_data_out[0] scanchain_117/module_data_out[1] scanchain_117/module_data_out[2]
+ scanchain_117/module_data_out[3] scanchain_117/module_data_out[4] scanchain_117/module_data_out[5]
+ scanchain_117/module_data_out[6] scanchain_117/module_data_out[7] vccd1 vssd1 user_module_361728533238569985
Xuser_module_361728533238569985_106 scanchain_106/module_data_in[0] scanchain_106/module_data_in[1]
+ scanchain_106/module_data_in[2] scanchain_106/module_data_in[3] scanchain_106/module_data_in[4]
+ scanchain_106/module_data_in[5] scanchain_106/module_data_in[6] scanchain_106/module_data_in[7]
+ scanchain_106/module_data_out[0] scanchain_106/module_data_out[1] scanchain_106/module_data_out[2]
+ scanchain_106/module_data_out[3] scanchain_106/module_data_out[4] scanchain_106/module_data_out[5]
+ scanchain_106/module_data_out[6] scanchain_106/module_data_out[7] vccd1 vssd1 user_module_361728533238569985
Xuser_module_361728533238569985_139 scanchain_139/module_data_in[0] scanchain_139/module_data_in[1]
+ scanchain_139/module_data_in[2] scanchain_139/module_data_in[3] scanchain_139/module_data_in[4]
+ scanchain_139/module_data_in[5] scanchain_139/module_data_in[6] scanchain_139/module_data_in[7]
+ scanchain_139/module_data_out[0] scanchain_139/module_data_out[1] scanchain_139/module_data_out[2]
+ scanchain_139/module_data_out[3] scanchain_139/module_data_out[4] scanchain_139/module_data_out[5]
+ scanchain_139/module_data_out[6] scanchain_139/module_data_out[7] vccd1 vssd1 user_module_361728533238569985
Xdiferential_muxpga_017 scanchain_017/module_data_in[0] scanchain_017/module_data_in[1]
+ scanchain_017/module_data_in[2] scanchain_017/module_data_in[3] scanchain_017/module_data_in[4]
+ scanchain_017/module_data_in[5] scanchain_017/module_data_in[6] scanchain_017/module_data_in[7]
+ scanchain_017/module_data_out[0] scanchain_017/module_data_out[1] scanchain_017/module_data_out[2]
+ scanchain_017/module_data_out[3] scanchain_017/module_data_out[4] scanchain_017/module_data_out[5]
+ scanchain_017/module_data_out[6] scanchain_017/module_data_out[7] vccd1 vssd1 diferential_muxpga
Xscanchain_140 scanchain_140/clk_in scanchain_141/clk_in scanchain_140/data_in scanchain_141/data_in
+ scanchain_140/latch_enable_in scanchain_141/latch_enable_in scanchain_140/module_data_in[0]
+ scanchain_140/module_data_in[1] scanchain_140/module_data_in[2] scanchain_140/module_data_in[3]
+ scanchain_140/module_data_in[4] scanchain_140/module_data_in[5] scanchain_140/module_data_in[6]
+ scanchain_140/module_data_in[7] scanchain_140/module_data_out[0] scanchain_140/module_data_out[1]
+ scanchain_140/module_data_out[2] scanchain_140/module_data_out[3] scanchain_140/module_data_out[4]
+ scanchain_140/module_data_out[5] scanchain_140/module_data_out[6] scanchain_140/module_data_out[7]
+ scanchain_140/scan_select_in scanchain_141/scan_select_in vccd1 vssd1 scanchain
Xscanchain_151 scanchain_151/clk_in scanchain_152/clk_in scanchain_151/data_in scanchain_152/data_in
+ scanchain_151/latch_enable_in scanchain_152/latch_enable_in scanchain_151/module_data_in[0]
+ scanchain_151/module_data_in[1] scanchain_151/module_data_in[2] scanchain_151/module_data_in[3]
+ scanchain_151/module_data_in[4] scanchain_151/module_data_in[5] scanchain_151/module_data_in[6]
+ scanchain_151/module_data_in[7] scanchain_151/module_data_out[0] scanchain_151/module_data_out[1]
+ scanchain_151/module_data_out[2] scanchain_151/module_data_out[3] scanchain_151/module_data_out[4]
+ scanchain_151/module_data_out[5] scanchain_151/module_data_out[6] scanchain_151/module_data_out[7]
+ scanchain_151/scan_select_in scanchain_152/scan_select_in vccd1 vssd1 scanchain
Xscanchain_195 scanchain_195/clk_in scanchain_196/clk_in scanchain_195/data_in scanchain_196/data_in
+ scanchain_195/latch_enable_in scanchain_196/latch_enable_in scanchain_195/module_data_in[0]
+ scanchain_195/module_data_in[1] scanchain_195/module_data_in[2] scanchain_195/module_data_in[3]
+ scanchain_195/module_data_in[4] scanchain_195/module_data_in[5] scanchain_195/module_data_in[6]
+ scanchain_195/module_data_in[7] scanchain_195/module_data_out[0] scanchain_195/module_data_out[1]
+ scanchain_195/module_data_out[2] scanchain_195/module_data_out[3] scanchain_195/module_data_out[4]
+ scanchain_195/module_data_out[5] scanchain_195/module_data_out[6] scanchain_195/module_data_out[7]
+ scanchain_195/scan_select_in scanchain_196/scan_select_in vccd1 vssd1 scanchain
Xscanchain_184 scanchain_184/clk_in scanchain_185/clk_in scanchain_184/data_in scanchain_185/data_in
+ scanchain_184/latch_enable_in scanchain_185/latch_enable_in scanchain_184/module_data_in[0]
+ scanchain_184/module_data_in[1] scanchain_184/module_data_in[2] scanchain_184/module_data_in[3]
+ scanchain_184/module_data_in[4] scanchain_184/module_data_in[5] scanchain_184/module_data_in[6]
+ scanchain_184/module_data_in[7] scanchain_184/module_data_out[0] scanchain_184/module_data_out[1]
+ scanchain_184/module_data_out[2] scanchain_184/module_data_out[3] scanchain_184/module_data_out[4]
+ scanchain_184/module_data_out[5] scanchain_184/module_data_out[6] scanchain_184/module_data_out[7]
+ scanchain_184/scan_select_in scanchain_185/scan_select_in vccd1 vssd1 scanchain
Xscanchain_173 scanchain_173/clk_in scanchain_174/clk_in scanchain_173/data_in scanchain_174/data_in
+ scanchain_173/latch_enable_in scanchain_174/latch_enable_in scanchain_173/module_data_in[0]
+ scanchain_173/module_data_in[1] scanchain_173/module_data_in[2] scanchain_173/module_data_in[3]
+ scanchain_173/module_data_in[4] scanchain_173/module_data_in[5] scanchain_173/module_data_in[6]
+ scanchain_173/module_data_in[7] scanchain_173/module_data_out[0] scanchain_173/module_data_out[1]
+ scanchain_173/module_data_out[2] scanchain_173/module_data_out[3] scanchain_173/module_data_out[4]
+ scanchain_173/module_data_out[5] scanchain_173/module_data_out[6] scanchain_173/module_data_out[7]
+ scanchain_173/scan_select_in scanchain_174/scan_select_in vccd1 vssd1 scanchain
Xscanchain_162 scanchain_162/clk_in scanchain_163/clk_in scanchain_162/data_in scanchain_163/data_in
+ scanchain_162/latch_enable_in scanchain_163/latch_enable_in scanchain_162/module_data_in[0]
+ scanchain_162/module_data_in[1] scanchain_162/module_data_in[2] scanchain_162/module_data_in[3]
+ scanchain_162/module_data_in[4] scanchain_162/module_data_in[5] scanchain_162/module_data_in[6]
+ scanchain_162/module_data_in[7] scanchain_162/module_data_out[0] scanchain_162/module_data_out[1]
+ scanchain_162/module_data_out[2] scanchain_162/module_data_out[3] scanchain_162/module_data_out[4]
+ scanchain_162/module_data_out[5] scanchain_162/module_data_out[6] scanchain_162/module_data_out[7]
+ scanchain_162/scan_select_in scanchain_163/scan_select_in vccd1 vssd1 scanchain
Xuser_module_360295047631610881_038 scanchain_038/module_data_in[0] scanchain_038/module_data_in[1]
+ scanchain_038/module_data_in[2] scanchain_038/module_data_in[3] scanchain_038/module_data_in[4]
+ scanchain_038/module_data_in[5] scanchain_038/module_data_in[6] scanchain_038/module_data_in[7]
+ scanchain_038/module_data_out[0] scanchain_038/module_data_out[1] scanchain_038/module_data_out[2]
+ scanchain_038/module_data_out[3] scanchain_038/module_data_out[4] scanchain_038/module_data_out[5]
+ scanchain_038/module_data_out[6] scanchain_038/module_data_out[7] vccd1 vssd1 user_module_360295047631610881
Xuser_module_361728533238569985_118 scanchain_118/module_data_in[0] scanchain_118/module_data_in[1]
+ scanchain_118/module_data_in[2] scanchain_118/module_data_in[3] scanchain_118/module_data_in[4]
+ scanchain_118/module_data_in[5] scanchain_118/module_data_in[6] scanchain_118/module_data_in[7]
+ scanchain_118/module_data_out[0] scanchain_118/module_data_out[1] scanchain_118/module_data_out[2]
+ scanchain_118/module_data_out[3] scanchain_118/module_data_out[4] scanchain_118/module_data_out[5]
+ scanchain_118/module_data_out[6] scanchain_118/module_data_out[7] vccd1 vssd1 user_module_361728533238569985
Xuser_module_361728533238569985_129 scanchain_129/module_data_in[0] scanchain_129/module_data_in[1]
+ scanchain_129/module_data_in[2] scanchain_129/module_data_in[3] scanchain_129/module_data_in[4]
+ scanchain_129/module_data_in[5] scanchain_129/module_data_in[6] scanchain_129/module_data_in[7]
+ scanchain_129/module_data_out[0] scanchain_129/module_data_out[1] scanchain_129/module_data_out[2]
+ scanchain_129/module_data_out[3] scanchain_129/module_data_out[4] scanchain_129/module_data_out[5]
+ scanchain_129/module_data_out[6] scanchain_129/module_data_out[7] vccd1 vssd1 user_module_361728533238569985
Xuser_module_361728533238569985_107 scanchain_107/module_data_in[0] scanchain_107/module_data_in[1]
+ scanchain_107/module_data_in[2] scanchain_107/module_data_in[3] scanchain_107/module_data_in[4]
+ scanchain_107/module_data_in[5] scanchain_107/module_data_in[6] scanchain_107/module_data_in[7]
+ scanchain_107/module_data_out[0] scanchain_107/module_data_out[1] scanchain_107/module_data_out[2]
+ scanchain_107/module_data_out[3] scanchain_107/module_data_out[4] scanchain_107/module_data_out[5]
+ scanchain_107/module_data_out[6] scanchain_107/module_data_out[7] vccd1 vssd1 user_module_361728533238569985
Xaidan_mcnay_PrimeDetector_026 scanchain_026/module_data_in[0] scanchain_026/module_data_in[1]
+ scanchain_026/module_data_in[2] scanchain_026/module_data_in[3] scanchain_026/module_data_in[4]
+ scanchain_026/module_data_in[5] scanchain_026/module_data_in[6] scanchain_026/module_data_in[7]
+ scanchain_026/module_data_out[0] scanchain_026/module_data_out[1] scanchain_026/module_data_out[2]
+ scanchain_026/module_data_out[3] scanchain_026/module_data_out[4] scanchain_026/module_data_out[5]
+ scanchain_026/module_data_out[6] scanchain_026/module_data_out[7] vccd1 vssd1 aidan_mcnay_PrimeDetector
Xs4ga_070 s4ga_070/io_in[0] s4ga_070/io_in[1] s4ga_070/io_in[2] s4ga_070/io_in[3]
+ s4ga_070/io_in[4] s4ga_070/io_in[5] s4ga_070/io_in[6] s4ga_070/io_in[7] s4ga_070/io_out[0]
+ s4ga_070/io_out[1] s4ga_070/io_out[2] s4ga_070/io_out[3] s4ga_070/io_out[4] s4ga_070/io_out[5]
+ s4ga_070/io_out[6] s4ga_070/io_out[7] vccd1 vssd1 s4ga
Xscanchain_130 scanchain_130/clk_in scanchain_131/clk_in scanchain_130/data_in scanchain_131/data_in
+ scanchain_130/latch_enable_in scanchain_131/latch_enable_in scanchain_130/module_data_in[0]
+ scanchain_130/module_data_in[1] scanchain_130/module_data_in[2] scanchain_130/module_data_in[3]
+ scanchain_130/module_data_in[4] scanchain_130/module_data_in[5] scanchain_130/module_data_in[6]
+ scanchain_130/module_data_in[7] scanchain_130/module_data_out[0] scanchain_130/module_data_out[1]
+ scanchain_130/module_data_out[2] scanchain_130/module_data_out[3] scanchain_130/module_data_out[4]
+ scanchain_130/module_data_out[5] scanchain_130/module_data_out[6] scanchain_130/module_data_out[7]
+ scanchain_130/scan_select_in scanchain_131/scan_select_in vccd1 vssd1 scanchain
Xscanchain_141 scanchain_141/clk_in scanchain_142/clk_in scanchain_141/data_in scanchain_142/data_in
+ scanchain_141/latch_enable_in scanchain_142/latch_enable_in scanchain_141/module_data_in[0]
+ scanchain_141/module_data_in[1] scanchain_141/module_data_in[2] scanchain_141/module_data_in[3]
+ scanchain_141/module_data_in[4] scanchain_141/module_data_in[5] scanchain_141/module_data_in[6]
+ scanchain_141/module_data_in[7] scanchain_141/module_data_out[0] scanchain_141/module_data_out[1]
+ scanchain_141/module_data_out[2] scanchain_141/module_data_out[3] scanchain_141/module_data_out[4]
+ scanchain_141/module_data_out[5] scanchain_141/module_data_out[6] scanchain_141/module_data_out[7]
+ scanchain_141/scan_select_in scanchain_142/scan_select_in vccd1 vssd1 scanchain
Xscanchain_152 scanchain_152/clk_in scanchain_153/clk_in scanchain_152/data_in scanchain_153/data_in
+ scanchain_152/latch_enable_in scanchain_153/latch_enable_in scanchain_152/module_data_in[0]
+ scanchain_152/module_data_in[1] scanchain_152/module_data_in[2] scanchain_152/module_data_in[3]
+ scanchain_152/module_data_in[4] scanchain_152/module_data_in[5] scanchain_152/module_data_in[6]
+ scanchain_152/module_data_in[7] scanchain_152/module_data_out[0] scanchain_152/module_data_out[1]
+ scanchain_152/module_data_out[2] scanchain_152/module_data_out[3] scanchain_152/module_data_out[4]
+ scanchain_152/module_data_out[5] scanchain_152/module_data_out[6] scanchain_152/module_data_out[7]
+ scanchain_152/scan_select_in scanchain_153/scan_select_in vccd1 vssd1 scanchain
Xscanchain_196 scanchain_196/clk_in scanchain_197/clk_in scanchain_196/data_in scanchain_197/data_in
+ scanchain_196/latch_enable_in scanchain_197/latch_enable_in scanchain_196/module_data_in[0]
+ scanchain_196/module_data_in[1] scanchain_196/module_data_in[2] scanchain_196/module_data_in[3]
+ scanchain_196/module_data_in[4] scanchain_196/module_data_in[5] scanchain_196/module_data_in[6]
+ scanchain_196/module_data_in[7] scanchain_196/module_data_out[0] scanchain_196/module_data_out[1]
+ scanchain_196/module_data_out[2] scanchain_196/module_data_out[3] scanchain_196/module_data_out[4]
+ scanchain_196/module_data_out[5] scanchain_196/module_data_out[6] scanchain_196/module_data_out[7]
+ scanchain_196/scan_select_in scanchain_197/scan_select_in vccd1 vssd1 scanchain
Xscanchain_185 scanchain_185/clk_in scanchain_186/clk_in scanchain_185/data_in scanchain_186/data_in
+ scanchain_185/latch_enable_in scanchain_186/latch_enable_in scanchain_185/module_data_in[0]
+ scanchain_185/module_data_in[1] scanchain_185/module_data_in[2] scanchain_185/module_data_in[3]
+ scanchain_185/module_data_in[4] scanchain_185/module_data_in[5] scanchain_185/module_data_in[6]
+ scanchain_185/module_data_in[7] scanchain_185/module_data_out[0] scanchain_185/module_data_out[1]
+ scanchain_185/module_data_out[2] scanchain_185/module_data_out[3] scanchain_185/module_data_out[4]
+ scanchain_185/module_data_out[5] scanchain_185/module_data_out[6] scanchain_185/module_data_out[7]
+ scanchain_185/scan_select_in scanchain_186/scan_select_in vccd1 vssd1 scanchain
Xscanchain_174 scanchain_174/clk_in scanchain_175/clk_in scanchain_174/data_in scanchain_175/data_in
+ scanchain_174/latch_enable_in scanchain_175/latch_enable_in scanchain_174/module_data_in[0]
+ scanchain_174/module_data_in[1] scanchain_174/module_data_in[2] scanchain_174/module_data_in[3]
+ scanchain_174/module_data_in[4] scanchain_174/module_data_in[5] scanchain_174/module_data_in[6]
+ scanchain_174/module_data_in[7] scanchain_174/module_data_out[0] scanchain_174/module_data_out[1]
+ scanchain_174/module_data_out[2] scanchain_174/module_data_out[3] scanchain_174/module_data_out[4]
+ scanchain_174/module_data_out[5] scanchain_174/module_data_out[6] scanchain_174/module_data_out[7]
+ scanchain_174/scan_select_in scanchain_175/scan_select_in vccd1 vssd1 scanchain
Xscanchain_163 scanchain_163/clk_in scanchain_164/clk_in scanchain_163/data_in scanchain_164/data_in
+ scanchain_163/latch_enable_in scanchain_164/latch_enable_in scanchain_163/module_data_in[0]
+ scanchain_163/module_data_in[1] scanchain_163/module_data_in[2] scanchain_163/module_data_in[3]
+ scanchain_163/module_data_in[4] scanchain_163/module_data_in[5] scanchain_163/module_data_in[6]
+ scanchain_163/module_data_in[7] scanchain_163/module_data_out[0] scanchain_163/module_data_out[1]
+ scanchain_163/module_data_out[2] scanchain_163/module_data_out[3] scanchain_163/module_data_out[4]
+ scanchain_163/module_data_out[5] scanchain_163/module_data_out[6] scanchain_163/module_data_out[7]
+ scanchain_163/scan_select_in scanchain_164/scan_select_in vccd1 vssd1 scanchain
Xuser_module_347140425276981843_087 scanchain_087/module_data_in[0] scanchain_087/module_data_in[1]
+ scanchain_087/module_data_in[2] scanchain_087/module_data_in[3] scanchain_087/module_data_in[4]
+ scanchain_087/module_data_in[5] scanchain_087/module_data_in[6] scanchain_087/module_data_in[7]
+ scanchain_087/module_data_out[0] scanchain_087/module_data_out[1] scanchain_087/module_data_out[2]
+ scanchain_087/module_data_out[3] scanchain_087/module_data_out[4] scanchain_087/module_data_out[5]
+ scanchain_087/module_data_out[6] scanchain_087/module_data_out[7] vccd1 vssd1 user_module_347140425276981843
Xuser_module_357106633951414273_008 scanchain_008/module_data_in[0] scanchain_008/module_data_in[1]
+ scanchain_008/module_data_in[2] scanchain_008/module_data_in[3] scanchain_008/module_data_in[4]
+ scanchain_008/module_data_in[5] scanchain_008/module_data_in[6] scanchain_008/module_data_in[7]
+ scanchain_008/module_data_out[0] scanchain_008/module_data_out[1] scanchain_008/module_data_out[2]
+ scanchain_008/module_data_out[3] scanchain_008/module_data_out[4] scanchain_008/module_data_out[5]
+ scanchain_008/module_data_out[6] scanchain_008/module_data_out[7] vccd1 vssd1 user_module_357106633951414273
Xuser_module_361728533238569985_119 scanchain_119/module_data_in[0] scanchain_119/module_data_in[1]
+ scanchain_119/module_data_in[2] scanchain_119/module_data_in[3] scanchain_119/module_data_in[4]
+ scanchain_119/module_data_in[5] scanchain_119/module_data_in[6] scanchain_119/module_data_in[7]
+ scanchain_119/module_data_out[0] scanchain_119/module_data_out[1] scanchain_119/module_data_out[2]
+ scanchain_119/module_data_out[3] scanchain_119/module_data_out[4] scanchain_119/module_data_out[5]
+ scanchain_119/module_data_out[6] scanchain_119/module_data_out[7] vccd1 vssd1 user_module_361728533238569985
Xuser_module_361728533238569985_108 scanchain_108/module_data_in[0] scanchain_108/module_data_in[1]
+ scanchain_108/module_data_in[2] scanchain_108/module_data_in[3] scanchain_108/module_data_in[4]
+ scanchain_108/module_data_in[5] scanchain_108/module_data_in[6] scanchain_108/module_data_in[7]
+ scanchain_108/module_data_out[0] scanchain_108/module_data_out[1] scanchain_108/module_data_out[2]
+ scanchain_108/module_data_out[3] scanchain_108/module_data_out[4] scanchain_108/module_data_out[5]
+ scanchain_108/module_data_out[6] scanchain_108/module_data_out[7] vccd1 vssd1 user_module_361728533238569985
Xscanchain_131 scanchain_131/clk_in scanchain_132/clk_in scanchain_131/data_in scanchain_132/data_in
+ scanchain_131/latch_enable_in scanchain_132/latch_enable_in scanchain_131/module_data_in[0]
+ scanchain_131/module_data_in[1] scanchain_131/module_data_in[2] scanchain_131/module_data_in[3]
+ scanchain_131/module_data_in[4] scanchain_131/module_data_in[5] scanchain_131/module_data_in[6]
+ scanchain_131/module_data_in[7] scanchain_131/module_data_out[0] scanchain_131/module_data_out[1]
+ scanchain_131/module_data_out[2] scanchain_131/module_data_out[3] scanchain_131/module_data_out[4]
+ scanchain_131/module_data_out[5] scanchain_131/module_data_out[6] scanchain_131/module_data_out[7]
+ scanchain_131/scan_select_in scanchain_132/scan_select_in vccd1 vssd1 scanchain
Xscanchain_120 scanchain_120/clk_in scanchain_121/clk_in scanchain_120/data_in scanchain_121/data_in
+ scanchain_120/latch_enable_in scanchain_121/latch_enable_in scanchain_120/module_data_in[0]
+ scanchain_120/module_data_in[1] scanchain_120/module_data_in[2] scanchain_120/module_data_in[3]
+ scanchain_120/module_data_in[4] scanchain_120/module_data_in[5] scanchain_120/module_data_in[6]
+ scanchain_120/module_data_in[7] scanchain_120/module_data_out[0] scanchain_120/module_data_out[1]
+ scanchain_120/module_data_out[2] scanchain_120/module_data_out[3] scanchain_120/module_data_out[4]
+ scanchain_120/module_data_out[5] scanchain_120/module_data_out[6] scanchain_120/module_data_out[7]
+ scanchain_120/scan_select_in scanchain_121/scan_select_in vccd1 vssd1 scanchain
Xscanchain_142 scanchain_142/clk_in scanchain_143/clk_in scanchain_142/data_in scanchain_143/data_in
+ scanchain_142/latch_enable_in scanchain_143/latch_enable_in scanchain_142/module_data_in[0]
+ scanchain_142/module_data_in[1] scanchain_142/module_data_in[2] scanchain_142/module_data_in[3]
+ scanchain_142/module_data_in[4] scanchain_142/module_data_in[5] scanchain_142/module_data_in[6]
+ scanchain_142/module_data_in[7] scanchain_142/module_data_out[0] scanchain_142/module_data_out[1]
+ scanchain_142/module_data_out[2] scanchain_142/module_data_out[3] scanchain_142/module_data_out[4]
+ scanchain_142/module_data_out[5] scanchain_142/module_data_out[6] scanchain_142/module_data_out[7]
+ scanchain_142/scan_select_in scanchain_143/scan_select_in vccd1 vssd1 scanchain
Xscanchain_197 scanchain_197/clk_in scanchain_198/clk_in scanchain_197/data_in scanchain_198/data_in
+ scanchain_197/latch_enable_in scanchain_198/latch_enable_in scanchain_197/module_data_in[0]
+ scanchain_197/module_data_in[1] scanchain_197/module_data_in[2] scanchain_197/module_data_in[3]
+ scanchain_197/module_data_in[4] scanchain_197/module_data_in[5] scanchain_197/module_data_in[6]
+ scanchain_197/module_data_in[7] scanchain_197/module_data_out[0] scanchain_197/module_data_out[1]
+ scanchain_197/module_data_out[2] scanchain_197/module_data_out[3] scanchain_197/module_data_out[4]
+ scanchain_197/module_data_out[5] scanchain_197/module_data_out[6] scanchain_197/module_data_out[7]
+ scanchain_197/scan_select_in scanchain_198/scan_select_in vccd1 vssd1 scanchain
Xscanchain_186 scanchain_186/clk_in scanchain_187/clk_in scanchain_186/data_in scanchain_187/data_in
+ scanchain_186/latch_enable_in scanchain_187/latch_enable_in scanchain_186/module_data_in[0]
+ scanchain_186/module_data_in[1] scanchain_186/module_data_in[2] scanchain_186/module_data_in[3]
+ scanchain_186/module_data_in[4] scanchain_186/module_data_in[5] scanchain_186/module_data_in[6]
+ scanchain_186/module_data_in[7] scanchain_186/module_data_out[0] scanchain_186/module_data_out[1]
+ scanchain_186/module_data_out[2] scanchain_186/module_data_out[3] scanchain_186/module_data_out[4]
+ scanchain_186/module_data_out[5] scanchain_186/module_data_out[6] scanchain_186/module_data_out[7]
+ scanchain_186/scan_select_in scanchain_187/scan_select_in vccd1 vssd1 scanchain
Xscanchain_175 scanchain_175/clk_in scanchain_176/clk_in scanchain_175/data_in scanchain_176/data_in
+ scanchain_175/latch_enable_in scanchain_176/latch_enable_in scanchain_175/module_data_in[0]
+ scanchain_175/module_data_in[1] scanchain_175/module_data_in[2] scanchain_175/module_data_in[3]
+ scanchain_175/module_data_in[4] scanchain_175/module_data_in[5] scanchain_175/module_data_in[6]
+ scanchain_175/module_data_in[7] scanchain_175/module_data_out[0] scanchain_175/module_data_out[1]
+ scanchain_175/module_data_out[2] scanchain_175/module_data_out[3] scanchain_175/module_data_out[4]
+ scanchain_175/module_data_out[5] scanchain_175/module_data_out[6] scanchain_175/module_data_out[7]
+ scanchain_175/scan_select_in scanchain_176/scan_select_in vccd1 vssd1 scanchain
Xscanchain_164 scanchain_164/clk_in scanchain_165/clk_in scanchain_164/data_in scanchain_165/data_in
+ scanchain_164/latch_enable_in scanchain_165/latch_enable_in scanchain_164/module_data_in[0]
+ scanchain_164/module_data_in[1] scanchain_164/module_data_in[2] scanchain_164/module_data_in[3]
+ scanchain_164/module_data_in[4] scanchain_164/module_data_in[5] scanchain_164/module_data_in[6]
+ scanchain_164/module_data_in[7] scanchain_164/module_data_out[0] scanchain_164/module_data_out[1]
+ scanchain_164/module_data_out[2] scanchain_164/module_data_out[3] scanchain_164/module_data_out[4]
+ scanchain_164/module_data_out[5] scanchain_164/module_data_out[6] scanchain_164/module_data_out[7]
+ scanchain_164/scan_select_in scanchain_165/scan_select_in vccd1 vssd1 scanchain
Xscanchain_153 scanchain_153/clk_in scanchain_154/clk_in scanchain_153/data_in scanchain_154/data_in
+ scanchain_153/latch_enable_in scanchain_154/latch_enable_in scanchain_153/module_data_in[0]
+ scanchain_153/module_data_in[1] scanchain_153/module_data_in[2] scanchain_153/module_data_in[3]
+ scanchain_153/module_data_in[4] scanchain_153/module_data_in[5] scanchain_153/module_data_in[6]
+ scanchain_153/module_data_in[7] scanchain_153/module_data_out[0] scanchain_153/module_data_out[1]
+ scanchain_153/module_data_out[2] scanchain_153/module_data_out[3] scanchain_153/module_data_out[4]
+ scanchain_153/module_data_out[5] scanchain_153/module_data_out[6] scanchain_153/module_data_out[7]
+ scanchain_153/scan_select_in scanchain_154/scan_select_in vccd1 vssd1 scanchain
Xdiferential_rvb3_024 diferential_rvb3_024/io_in[0] diferential_rvb3_024/io_in[1]
+ diferential_rvb3_024/io_in[2] diferential_rvb3_024/io_in[3] diferential_rvb3_024/io_in[4]
+ diferential_rvb3_024/io_in[5] diferential_rvb3_024/io_in[6] diferential_rvb3_024/io_in[7]
+ diferential_rvb3_024/io_out[0] diferential_rvb3_024/io_out[1] diferential_rvb3_024/io_out[2]
+ diferential_rvb3_024/io_out[3] diferential_rvb3_024/io_out[4] diferential_rvb3_024/io_out[5]
+ diferential_rvb3_024/io_out[6] diferential_rvb3_024/io_out[7] vccd1 vssd1 diferential_rvb3
Xkiwih_tt_top_045 kiwih_tt_top_045/io_in[0] kiwih_tt_top_045/io_in[1] kiwih_tt_top_045/io_in[2]
+ kiwih_tt_top_045/io_in[3] kiwih_tt_top_045/io_in[4] kiwih_tt_top_045/io_in[5] kiwih_tt_top_045/io_in[6]
+ kiwih_tt_top_045/io_in[7] kiwih_tt_top_045/io_out[0] kiwih_tt_top_045/io_out[1]
+ kiwih_tt_top_045/io_out[2] kiwih_tt_top_045/io_out[3] kiwih_tt_top_045/io_out[4]
+ kiwih_tt_top_045/io_out[5] kiwih_tt_top_045/io_out[6] kiwih_tt_top_045/io_out[7]
+ vccd1 vssd1 kiwih_tt_top
Xuser_module_361728533238569985_109 scanchain_109/module_data_in[0] scanchain_109/module_data_in[1]
+ scanchain_109/module_data_in[2] scanchain_109/module_data_in[3] scanchain_109/module_data_in[4]
+ scanchain_109/module_data_in[5] scanchain_109/module_data_in[6] scanchain_109/module_data_in[7]
+ scanchain_109/module_data_out[0] scanchain_109/module_data_out[1] scanchain_109/module_data_out[2]
+ scanchain_109/module_data_out[3] scanchain_109/module_data_out[4] scanchain_109/module_data_out[5]
+ scanchain_109/module_data_out[6] scanchain_109/module_data_out[7] vccd1 vssd1 user_module_361728533238569985
Xmorningjava_top_001 morningjava_top_001/io_in[0] morningjava_top_001/io_in[1] morningjava_top_001/io_in[2]
+ morningjava_top_001/io_in[3] morningjava_top_001/io_in[4] morningjava_top_001/io_in[5]
+ morningjava_top_001/io_in[6] morningjava_top_001/io_in[7] morningjava_top_001/io_out[0]
+ morningjava_top_001/io_out[1] morningjava_top_001/io_out[2] morningjava_top_001/io_out[3]
+ morningjava_top_001/io_out[4] morningjava_top_001/io_out[5] morningjava_top_001/io_out[6]
+ morningjava_top_001/io_out[7] vccd1 vssd1 morningjava_top
Xscanchain_121 scanchain_121/clk_in scanchain_122/clk_in scanchain_121/data_in scanchain_122/data_in
+ scanchain_121/latch_enable_in scanchain_122/latch_enable_in scanchain_121/module_data_in[0]
+ scanchain_121/module_data_in[1] scanchain_121/module_data_in[2] scanchain_121/module_data_in[3]
+ scanchain_121/module_data_in[4] scanchain_121/module_data_in[5] scanchain_121/module_data_in[6]
+ scanchain_121/module_data_in[7] scanchain_121/module_data_out[0] scanchain_121/module_data_out[1]
+ scanchain_121/module_data_out[2] scanchain_121/module_data_out[3] scanchain_121/module_data_out[4]
+ scanchain_121/module_data_out[5] scanchain_121/module_data_out[6] scanchain_121/module_data_out[7]
+ scanchain_121/scan_select_in scanchain_122/scan_select_in vccd1 vssd1 scanchain
Xscanchain_132 scanchain_132/clk_in scanchain_133/clk_in scanchain_132/data_in scanchain_133/data_in
+ scanchain_132/latch_enable_in scanchain_133/latch_enable_in scanchain_132/module_data_in[0]
+ scanchain_132/module_data_in[1] scanchain_132/module_data_in[2] scanchain_132/module_data_in[3]
+ scanchain_132/module_data_in[4] scanchain_132/module_data_in[5] scanchain_132/module_data_in[6]
+ scanchain_132/module_data_in[7] scanchain_132/module_data_out[0] scanchain_132/module_data_out[1]
+ scanchain_132/module_data_out[2] scanchain_132/module_data_out[3] scanchain_132/module_data_out[4]
+ scanchain_132/module_data_out[5] scanchain_132/module_data_out[6] scanchain_132/module_data_out[7]
+ scanchain_132/scan_select_in scanchain_133/scan_select_in vccd1 vssd1 scanchain
Xscanchain_143 scanchain_143/clk_in scanchain_144/clk_in scanchain_143/data_in scanchain_144/data_in
+ scanchain_143/latch_enable_in scanchain_144/latch_enable_in scanchain_143/module_data_in[0]
+ scanchain_143/module_data_in[1] scanchain_143/module_data_in[2] scanchain_143/module_data_in[3]
+ scanchain_143/module_data_in[4] scanchain_143/module_data_in[5] scanchain_143/module_data_in[6]
+ scanchain_143/module_data_in[7] scanchain_143/module_data_out[0] scanchain_143/module_data_out[1]
+ scanchain_143/module_data_out[2] scanchain_143/module_data_out[3] scanchain_143/module_data_out[4]
+ scanchain_143/module_data_out[5] scanchain_143/module_data_out[6] scanchain_143/module_data_out[7]
+ scanchain_143/scan_select_in scanchain_144/scan_select_in vccd1 vssd1 scanchain
Xscanchain_110 scanchain_110/clk_in scanchain_111/clk_in scanchain_110/data_in scanchain_111/data_in
+ scanchain_110/latch_enable_in scanchain_111/latch_enable_in scanchain_110/module_data_in[0]
+ scanchain_110/module_data_in[1] scanchain_110/module_data_in[2] scanchain_110/module_data_in[3]
+ scanchain_110/module_data_in[4] scanchain_110/module_data_in[5] scanchain_110/module_data_in[6]
+ scanchain_110/module_data_in[7] scanchain_110/module_data_out[0] scanchain_110/module_data_out[1]
+ scanchain_110/module_data_out[2] scanchain_110/module_data_out[3] scanchain_110/module_data_out[4]
+ scanchain_110/module_data_out[5] scanchain_110/module_data_out[6] scanchain_110/module_data_out[7]
+ scanchain_110/scan_select_in scanchain_111/scan_select_in vccd1 vssd1 scanchain
Xuser_module_357897381919942657_007 scanchain_007/module_data_in[0] scanchain_007/module_data_in[1]
+ scanchain_007/module_data_in[2] scanchain_007/module_data_in[3] scanchain_007/module_data_in[4]
+ scanchain_007/module_data_in[5] scanchain_007/module_data_in[6] scanchain_007/module_data_in[7]
+ scanchain_007/module_data_out[0] scanchain_007/module_data_out[1] scanchain_007/module_data_out[2]
+ scanchain_007/module_data_out[3] scanchain_007/module_data_out[4] scanchain_007/module_data_out[5]
+ scanchain_007/module_data_out[6] scanchain_007/module_data_out[7] vccd1 vssd1 user_module_357897381919942657
Xscanchain_198 scanchain_198/clk_in scanchain_199/clk_in scanchain_198/data_in scanchain_199/data_in
+ scanchain_198/latch_enable_in scanchain_199/latch_enable_in scanchain_198/module_data_in[0]
+ scanchain_198/module_data_in[1] scanchain_198/module_data_in[2] scanchain_198/module_data_in[3]
+ scanchain_198/module_data_in[4] scanchain_198/module_data_in[5] scanchain_198/module_data_in[6]
+ scanchain_198/module_data_in[7] scanchain_198/module_data_out[0] scanchain_198/module_data_out[1]
+ scanchain_198/module_data_out[2] scanchain_198/module_data_out[3] scanchain_198/module_data_out[4]
+ scanchain_198/module_data_out[5] scanchain_198/module_data_out[6] scanchain_198/module_data_out[7]
+ scanchain_198/scan_select_in scanchain_199/scan_select_in vccd1 vssd1 scanchain
Xscanchain_187 scanchain_187/clk_in scanchain_188/clk_in scanchain_187/data_in scanchain_188/data_in
+ scanchain_187/latch_enable_in scanchain_188/latch_enable_in scanchain_187/module_data_in[0]
+ scanchain_187/module_data_in[1] scanchain_187/module_data_in[2] scanchain_187/module_data_in[3]
+ scanchain_187/module_data_in[4] scanchain_187/module_data_in[5] scanchain_187/module_data_in[6]
+ scanchain_187/module_data_in[7] scanchain_187/module_data_out[0] scanchain_187/module_data_out[1]
+ scanchain_187/module_data_out[2] scanchain_187/module_data_out[3] scanchain_187/module_data_out[4]
+ scanchain_187/module_data_out[5] scanchain_187/module_data_out[6] scanchain_187/module_data_out[7]
+ scanchain_187/scan_select_in scanchain_188/scan_select_in vccd1 vssd1 scanchain
Xscanchain_176 scanchain_176/clk_in scanchain_177/clk_in scanchain_176/data_in scanchain_177/data_in
+ scanchain_176/latch_enable_in scanchain_177/latch_enable_in scanchain_176/module_data_in[0]
+ scanchain_176/module_data_in[1] scanchain_176/module_data_in[2] scanchain_176/module_data_in[3]
+ scanchain_176/module_data_in[4] scanchain_176/module_data_in[5] scanchain_176/module_data_in[6]
+ scanchain_176/module_data_in[7] scanchain_176/module_data_out[0] scanchain_176/module_data_out[1]
+ scanchain_176/module_data_out[2] scanchain_176/module_data_out[3] scanchain_176/module_data_out[4]
+ scanchain_176/module_data_out[5] scanchain_176/module_data_out[6] scanchain_176/module_data_out[7]
+ scanchain_176/scan_select_in scanchain_177/scan_select_in vccd1 vssd1 scanchain
Xscanchain_165 scanchain_165/clk_in scanchain_166/clk_in scanchain_165/data_in scanchain_166/data_in
+ scanchain_165/latch_enable_in scanchain_166/latch_enable_in scanchain_165/module_data_in[0]
+ scanchain_165/module_data_in[1] scanchain_165/module_data_in[2] scanchain_165/module_data_in[3]
+ scanchain_165/module_data_in[4] scanchain_165/module_data_in[5] scanchain_165/module_data_in[6]
+ scanchain_165/module_data_in[7] scanchain_165/module_data_out[0] scanchain_165/module_data_out[1]
+ scanchain_165/module_data_out[2] scanchain_165/module_data_out[3] scanchain_165/module_data_out[4]
+ scanchain_165/module_data_out[5] scanchain_165/module_data_out[6] scanchain_165/module_data_out[7]
+ scanchain_165/scan_select_in scanchain_166/scan_select_in vccd1 vssd1 scanchain
Xscanchain_154 scanchain_154/clk_in scanchain_155/clk_in scanchain_154/data_in scanchain_155/data_in
+ scanchain_154/latch_enable_in scanchain_155/latch_enable_in scanchain_154/module_data_in[0]
+ scanchain_154/module_data_in[1] scanchain_154/module_data_in[2] scanchain_154/module_data_in[3]
+ scanchain_154/module_data_in[4] scanchain_154/module_data_in[5] scanchain_154/module_data_in[6]
+ scanchain_154/module_data_in[7] scanchain_154/module_data_out[0] scanchain_154/module_data_out[1]
+ scanchain_154/module_data_out[2] scanchain_154/module_data_out[3] scanchain_154/module_data_out[4]
+ scanchain_154/module_data_out[5] scanchain_154/module_data_out[6] scanchain_154/module_data_out[7]
+ scanchain_154/scan_select_in scanchain_155/scan_select_in vccd1 vssd1 scanchain
Xpsychogenic_neptunefixed_052 scanchain_052/module_data_in[0] scanchain_052/module_data_in[1]
+ scanchain_052/module_data_in[2] scanchain_052/module_data_in[3] scanchain_052/module_data_in[4]
+ scanchain_052/module_data_in[5] scanchain_052/module_data_in[6] scanchain_052/module_data_in[7]
+ scanchain_052/module_data_out[0] scanchain_052/module_data_out[1] scanchain_052/module_data_out[2]
+ scanchain_052/module_data_out[3] scanchain_052/module_data_out[4] scanchain_052/module_data_out[5]
+ scanchain_052/module_data_out[6] scanchain_052/module_data_out[7] vccd1 vssd1 psychogenic_neptunefixed
Xuser_module_354091612057990145_018 scanchain_018/module_data_in[0] scanchain_018/module_data_in[1]
+ scanchain_018/module_data_in[2] scanchain_018/module_data_in[3] scanchain_018/module_data_in[4]
+ scanchain_018/module_data_in[5] scanchain_018/module_data_in[6] scanchain_018/module_data_in[7]
+ scanchain_018/module_data_out[0] scanchain_018/module_data_out[1] scanchain_018/module_data_out[2]
+ scanchain_018/module_data_out[3] scanchain_018/module_data_out[4] scanchain_018/module_data_out[5]
+ scanchain_018/module_data_out[6] scanchain_018/module_data_out[7] vccd1 vssd1 user_module_354091612057990145
Xscanchain_122 scanchain_122/clk_in scanchain_123/clk_in scanchain_122/data_in scanchain_123/data_in
+ scanchain_122/latch_enable_in scanchain_123/latch_enable_in scanchain_122/module_data_in[0]
+ scanchain_122/module_data_in[1] scanchain_122/module_data_in[2] scanchain_122/module_data_in[3]
+ scanchain_122/module_data_in[4] scanchain_122/module_data_in[5] scanchain_122/module_data_in[6]
+ scanchain_122/module_data_in[7] scanchain_122/module_data_out[0] scanchain_122/module_data_out[1]
+ scanchain_122/module_data_out[2] scanchain_122/module_data_out[3] scanchain_122/module_data_out[4]
+ scanchain_122/module_data_out[5] scanchain_122/module_data_out[6] scanchain_122/module_data_out[7]
+ scanchain_122/scan_select_in scanchain_123/scan_select_in vccd1 vssd1 scanchain
Xscanchain_133 scanchain_133/clk_in scanchain_134/clk_in scanchain_133/data_in scanchain_134/data_in
+ scanchain_133/latch_enable_in scanchain_134/latch_enable_in scanchain_133/module_data_in[0]
+ scanchain_133/module_data_in[1] scanchain_133/module_data_in[2] scanchain_133/module_data_in[3]
+ scanchain_133/module_data_in[4] scanchain_133/module_data_in[5] scanchain_133/module_data_in[6]
+ scanchain_133/module_data_in[7] scanchain_133/module_data_out[0] scanchain_133/module_data_out[1]
+ scanchain_133/module_data_out[2] scanchain_133/module_data_out[3] scanchain_133/module_data_out[4]
+ scanchain_133/module_data_out[5] scanchain_133/module_data_out[6] scanchain_133/module_data_out[7]
+ scanchain_133/scan_select_in scanchain_134/scan_select_in vccd1 vssd1 scanchain
Xscanchain_111 scanchain_111/clk_in scanchain_112/clk_in scanchain_111/data_in scanchain_112/data_in
+ scanchain_111/latch_enable_in scanchain_112/latch_enable_in scanchain_111/module_data_in[0]
+ scanchain_111/module_data_in[1] scanchain_111/module_data_in[2] scanchain_111/module_data_in[3]
+ scanchain_111/module_data_in[4] scanchain_111/module_data_in[5] scanchain_111/module_data_in[6]
+ scanchain_111/module_data_in[7] scanchain_111/module_data_out[0] scanchain_111/module_data_out[1]
+ scanchain_111/module_data_out[2] scanchain_111/module_data_out[3] scanchain_111/module_data_out[4]
+ scanchain_111/module_data_out[5] scanchain_111/module_data_out[6] scanchain_111/module_data_out[7]
+ scanchain_111/scan_select_in scanchain_112/scan_select_in vccd1 vssd1 scanchain
Xscanchain_144 scanchain_144/clk_in scanchain_145/clk_in scanchain_144/data_in scanchain_145/data_in
+ scanchain_144/latch_enable_in scanchain_145/latch_enable_in scanchain_144/module_data_in[0]
+ scanchain_144/module_data_in[1] scanchain_144/module_data_in[2] scanchain_144/module_data_in[3]
+ scanchain_144/module_data_in[4] scanchain_144/module_data_in[5] scanchain_144/module_data_in[6]
+ scanchain_144/module_data_in[7] scanchain_144/module_data_out[0] scanchain_144/module_data_out[1]
+ scanchain_144/module_data_out[2] scanchain_144/module_data_out[3] scanchain_144/module_data_out[4]
+ scanchain_144/module_data_out[5] scanchain_144/module_data_out[6] scanchain_144/module_data_out[7]
+ scanchain_144/scan_select_in scanchain_145/scan_select_in vccd1 vssd1 scanchain
Xscanchain_100 scanchain_100/clk_in scanchain_101/clk_in scanchain_100/data_in scanchain_101/data_in
+ scanchain_100/latch_enable_in scanchain_101/latch_enable_in scanchain_100/module_data_in[0]
+ scanchain_100/module_data_in[1] scanchain_100/module_data_in[2] scanchain_100/module_data_in[3]
+ scanchain_100/module_data_in[4] scanchain_100/module_data_in[5] scanchain_100/module_data_in[6]
+ scanchain_100/module_data_in[7] scanchain_100/module_data_out[0] scanchain_100/module_data_out[1]
+ scanchain_100/module_data_out[2] scanchain_100/module_data_out[3] scanchain_100/module_data_out[4]
+ scanchain_100/module_data_out[5] scanchain_100/module_data_out[6] scanchain_100/module_data_out[7]
+ scanchain_100/scan_select_in scanchain_101/scan_select_in vccd1 vssd1 scanchain
Xscanchain_166 scanchain_166/clk_in scanchain_167/clk_in scanchain_166/data_in scanchain_167/data_in
+ scanchain_166/latch_enable_in scanchain_167/latch_enable_in scanchain_166/module_data_in[0]
+ scanchain_166/module_data_in[1] scanchain_166/module_data_in[2] scanchain_166/module_data_in[3]
+ scanchain_166/module_data_in[4] scanchain_166/module_data_in[5] scanchain_166/module_data_in[6]
+ scanchain_166/module_data_in[7] scanchain_166/module_data_out[0] scanchain_166/module_data_out[1]
+ scanchain_166/module_data_out[2] scanchain_166/module_data_out[3] scanchain_166/module_data_out[4]
+ scanchain_166/module_data_out[5] scanchain_166/module_data_out[6] scanchain_166/module_data_out[7]
+ scanchain_166/scan_select_in scanchain_167/scan_select_in vccd1 vssd1 scanchain
Xscanchain_155 scanchain_155/clk_in scanchain_156/clk_in scanchain_155/data_in scanchain_156/data_in
+ scanchain_155/latch_enable_in scanchain_156/latch_enable_in scanchain_155/module_data_in[0]
+ scanchain_155/module_data_in[1] scanchain_155/module_data_in[2] scanchain_155/module_data_in[3]
+ scanchain_155/module_data_in[4] scanchain_155/module_data_in[5] scanchain_155/module_data_in[6]
+ scanchain_155/module_data_in[7] scanchain_155/module_data_out[0] scanchain_155/module_data_out[1]
+ scanchain_155/module_data_out[2] scanchain_155/module_data_out[3] scanchain_155/module_data_out[4]
+ scanchain_155/module_data_out[5] scanchain_155/module_data_out[6] scanchain_155/module_data_out[7]
+ scanchain_155/scan_select_in scanchain_156/scan_select_in vccd1 vssd1 scanchain
Xscanchain_199 scanchain_199/clk_in scanchain_200/clk_in scanchain_199/data_in scanchain_200/data_in
+ scanchain_199/latch_enable_in scanchain_200/latch_enable_in scanchain_199/module_data_in[0]
+ scanchain_199/module_data_in[1] scanchain_199/module_data_in[2] scanchain_199/module_data_in[3]
+ scanchain_199/module_data_in[4] scanchain_199/module_data_in[5] scanchain_199/module_data_in[6]
+ scanchain_199/module_data_in[7] scanchain_199/module_data_out[0] scanchain_199/module_data_out[1]
+ scanchain_199/module_data_out[2] scanchain_199/module_data_out[3] scanchain_199/module_data_out[4]
+ scanchain_199/module_data_out[5] scanchain_199/module_data_out[6] scanchain_199/module_data_out[7]
+ scanchain_199/scan_select_in scanchain_200/scan_select_in vccd1 vssd1 scanchain
Xscanchain_188 scanchain_188/clk_in scanchain_189/clk_in scanchain_188/data_in scanchain_189/data_in
+ scanchain_188/latch_enable_in scanchain_189/latch_enable_in scanchain_188/module_data_in[0]
+ scanchain_188/module_data_in[1] scanchain_188/module_data_in[2] scanchain_188/module_data_in[3]
+ scanchain_188/module_data_in[4] scanchain_188/module_data_in[5] scanchain_188/module_data_in[6]
+ scanchain_188/module_data_in[7] scanchain_188/module_data_out[0] scanchain_188/module_data_out[1]
+ scanchain_188/module_data_out[2] scanchain_188/module_data_out[3] scanchain_188/module_data_out[4]
+ scanchain_188/module_data_out[5] scanchain_188/module_data_out[6] scanchain_188/module_data_out[7]
+ scanchain_188/scan_select_in scanchain_189/scan_select_in vccd1 vssd1 scanchain
Xscanchain_177 scanchain_177/clk_in scanchain_178/clk_in scanchain_177/data_in scanchain_178/data_in
+ scanchain_177/latch_enable_in scanchain_178/latch_enable_in scanchain_177/module_data_in[0]
+ scanchain_177/module_data_in[1] scanchain_177/module_data_in[2] scanchain_177/module_data_in[3]
+ scanchain_177/module_data_in[4] scanchain_177/module_data_in[5] scanchain_177/module_data_in[6]
+ scanchain_177/module_data_in[7] scanchain_177/module_data_out[0] scanchain_177/module_data_out[1]
+ scanchain_177/module_data_out[2] scanchain_177/module_data_out[3] scanchain_177/module_data_out[4]
+ scanchain_177/module_data_out[5] scanchain_177/module_data_out[6] scanchain_177/module_data_out[7]
+ scanchain_177/scan_select_in scanchain_178/scan_select_in vccd1 vssd1 scanchain
Xuser_module_362371515213982721_077 scanchain_077/module_data_in[0] scanchain_077/module_data_in[1]
+ scanchain_077/module_data_in[2] scanchain_077/module_data_in[3] scanchain_077/module_data_in[4]
+ scanchain_077/module_data_in[5] scanchain_077/module_data_in[6] scanchain_077/module_data_in[7]
+ scanchain_077/module_data_out[0] scanchain_077/module_data_out[1] scanchain_077/module_data_out[2]
+ scanchain_077/module_data_out[3] scanchain_077/module_data_out[4] scanchain_077/module_data_out[5]
+ scanchain_077/module_data_out[6] scanchain_077/module_data_out[7] vccd1 vssd1 user_module_362371515213982721
Xuser_module_361728533238569985_090 scanchain_090/module_data_in[0] scanchain_090/module_data_in[1]
+ scanchain_090/module_data_in[2] scanchain_090/module_data_in[3] scanchain_090/module_data_in[4]
+ scanchain_090/module_data_in[5] scanchain_090/module_data_in[6] scanchain_090/module_data_in[7]
+ scanchain_090/module_data_out[0] scanchain_090/module_data_out[1] scanchain_090/module_data_out[2]
+ scanchain_090/module_data_out[3] scanchain_090/module_data_out[4] scanchain_090/module_data_out[5]
+ scanchain_090/module_data_out[6] scanchain_090/module_data_out[7] vccd1 vssd1 user_module_361728533238569985
Xuser_module_361728681519813633_071 scanchain_071/module_data_in[0] scanchain_071/module_data_in[1]
+ scanchain_071/module_data_in[2] scanchain_071/module_data_in[3] scanchain_071/module_data_in[4]
+ scanchain_071/module_data_in[5] scanchain_071/module_data_in[6] scanchain_071/module_data_in[7]
+ scanchain_071/module_data_out[0] scanchain_071/module_data_out[1] scanchain_071/module_data_out[2]
+ scanchain_071/module_data_out[3] scanchain_071/module_data_out[4] scanchain_071/module_data_out[5]
+ scanchain_071/module_data_out[6] scanchain_071/module_data_out[7] vccd1 vssd1 user_module_361728681519813633
Xmaheredia_arbiter_game_074 scanchain_074/module_data_in[0] scanchain_074/module_data_in[1]
+ scanchain_074/module_data_in[2] scanchain_074/module_data_in[3] scanchain_074/module_data_in[4]
+ scanchain_074/module_data_in[5] scanchain_074/module_data_in[6] scanchain_074/module_data_in[7]
+ scanchain_074/module_data_out[0] scanchain_074/module_data_out[1] scanchain_074/module_data_out[2]
+ scanchain_074/module_data_out[3] scanchain_074/module_data_out[4] scanchain_074/module_data_out[5]
+ scanchain_074/module_data_out[6] scanchain_074/module_data_out[7] vccd1 vssd1 maheredia_arbiter_game
Xmy_design_047 my_design_047/io_in[0] my_design_047/io_in[1] my_design_047/io_in[2]
+ my_design_047/io_in[3] my_design_047/io_in[4] my_design_047/io_in[5] my_design_047/io_in[6]
+ my_design_047/io_in[7] my_design_047/io_out[0] my_design_047/io_out[1] my_design_047/io_out[2]
+ my_design_047/io_out[3] my_design_047/io_out[4] my_design_047/io_out[5] my_design_047/io_out[6]
+ my_design_047/io_out[7] vccd1 vssd1 my_design
Xscanchain_123 scanchain_123/clk_in scanchain_124/clk_in scanchain_123/data_in scanchain_124/data_in
+ scanchain_123/latch_enable_in scanchain_124/latch_enable_in scanchain_123/module_data_in[0]
+ scanchain_123/module_data_in[1] scanchain_123/module_data_in[2] scanchain_123/module_data_in[3]
+ scanchain_123/module_data_in[4] scanchain_123/module_data_in[5] scanchain_123/module_data_in[6]
+ scanchain_123/module_data_in[7] scanchain_123/module_data_out[0] scanchain_123/module_data_out[1]
+ scanchain_123/module_data_out[2] scanchain_123/module_data_out[3] scanchain_123/module_data_out[4]
+ scanchain_123/module_data_out[5] scanchain_123/module_data_out[6] scanchain_123/module_data_out[7]
+ scanchain_123/scan_select_in scanchain_124/scan_select_in vccd1 vssd1 scanchain
Xscanchain_134 scanchain_134/clk_in scanchain_135/clk_in scanchain_134/data_in scanchain_135/data_in
+ scanchain_134/latch_enable_in scanchain_135/latch_enable_in scanchain_134/module_data_in[0]
+ scanchain_134/module_data_in[1] scanchain_134/module_data_in[2] scanchain_134/module_data_in[3]
+ scanchain_134/module_data_in[4] scanchain_134/module_data_in[5] scanchain_134/module_data_in[6]
+ scanchain_134/module_data_in[7] scanchain_134/module_data_out[0] scanchain_134/module_data_out[1]
+ scanchain_134/module_data_out[2] scanchain_134/module_data_out[3] scanchain_134/module_data_out[4]
+ scanchain_134/module_data_out[5] scanchain_134/module_data_out[6] scanchain_134/module_data_out[7]
+ scanchain_134/scan_select_in scanchain_135/scan_select_in vccd1 vssd1 scanchain
Xscanchain_112 scanchain_112/clk_in scanchain_113/clk_in scanchain_112/data_in scanchain_113/data_in
+ scanchain_112/latch_enable_in scanchain_113/latch_enable_in scanchain_112/module_data_in[0]
+ scanchain_112/module_data_in[1] scanchain_112/module_data_in[2] scanchain_112/module_data_in[3]
+ scanchain_112/module_data_in[4] scanchain_112/module_data_in[5] scanchain_112/module_data_in[6]
+ scanchain_112/module_data_in[7] scanchain_112/module_data_out[0] scanchain_112/module_data_out[1]
+ scanchain_112/module_data_out[2] scanchain_112/module_data_out[3] scanchain_112/module_data_out[4]
+ scanchain_112/module_data_out[5] scanchain_112/module_data_out[6] scanchain_112/module_data_out[7]
+ scanchain_112/scan_select_in scanchain_113/scan_select_in vccd1 vssd1 scanchain
Xscanchain_145 scanchain_145/clk_in scanchain_146/clk_in scanchain_145/data_in scanchain_146/data_in
+ scanchain_145/latch_enable_in scanchain_146/latch_enable_in scanchain_145/module_data_in[0]
+ scanchain_145/module_data_in[1] scanchain_145/module_data_in[2] scanchain_145/module_data_in[3]
+ scanchain_145/module_data_in[4] scanchain_145/module_data_in[5] scanchain_145/module_data_in[6]
+ scanchain_145/module_data_in[7] scanchain_145/module_data_out[0] scanchain_145/module_data_out[1]
+ scanchain_145/module_data_out[2] scanchain_145/module_data_out[3] scanchain_145/module_data_out[4]
+ scanchain_145/module_data_out[5] scanchain_145/module_data_out[6] scanchain_145/module_data_out[7]
+ scanchain_145/scan_select_in scanchain_146/scan_select_in vccd1 vssd1 scanchain
Xscanchain_101 scanchain_101/clk_in scanchain_102/clk_in scanchain_101/data_in scanchain_102/data_in
+ scanchain_101/latch_enable_in scanchain_102/latch_enable_in scanchain_101/module_data_in[0]
+ scanchain_101/module_data_in[1] scanchain_101/module_data_in[2] scanchain_101/module_data_in[3]
+ scanchain_101/module_data_in[4] scanchain_101/module_data_in[5] scanchain_101/module_data_in[6]
+ scanchain_101/module_data_in[7] scanchain_101/module_data_out[0] scanchain_101/module_data_out[1]
+ scanchain_101/module_data_out[2] scanchain_101/module_data_out[3] scanchain_101/module_data_out[4]
+ scanchain_101/module_data_out[5] scanchain_101/module_data_out[6] scanchain_101/module_data_out[7]
+ scanchain_101/scan_select_in scanchain_102/scan_select_in vccd1 vssd1 scanchain
Xscanchain_189 scanchain_189/clk_in scanchain_190/clk_in scanchain_189/data_in scanchain_190/data_in
+ scanchain_189/latch_enable_in scanchain_190/latch_enable_in scanchain_189/module_data_in[0]
+ scanchain_189/module_data_in[1] scanchain_189/module_data_in[2] scanchain_189/module_data_in[3]
+ scanchain_189/module_data_in[4] scanchain_189/module_data_in[5] scanchain_189/module_data_in[6]
+ scanchain_189/module_data_in[7] scanchain_189/module_data_out[0] scanchain_189/module_data_out[1]
+ scanchain_189/module_data_out[2] scanchain_189/module_data_out[3] scanchain_189/module_data_out[4]
+ scanchain_189/module_data_out[5] scanchain_189/module_data_out[6] scanchain_189/module_data_out[7]
+ scanchain_189/scan_select_in scanchain_190/scan_select_in vccd1 vssd1 scanchain
Xscanchain_167 scanchain_167/clk_in scanchain_168/clk_in scanchain_167/data_in scanchain_168/data_in
+ scanchain_167/latch_enable_in scanchain_168/latch_enable_in scanchain_167/module_data_in[0]
+ scanchain_167/module_data_in[1] scanchain_167/module_data_in[2] scanchain_167/module_data_in[3]
+ scanchain_167/module_data_in[4] scanchain_167/module_data_in[5] scanchain_167/module_data_in[6]
+ scanchain_167/module_data_in[7] scanchain_167/module_data_out[0] scanchain_167/module_data_out[1]
+ scanchain_167/module_data_out[2] scanchain_167/module_data_out[3] scanchain_167/module_data_out[4]
+ scanchain_167/module_data_out[5] scanchain_167/module_data_out[6] scanchain_167/module_data_out[7]
+ scanchain_167/scan_select_in scanchain_168/scan_select_in vccd1 vssd1 scanchain
Xscanchain_178 scanchain_178/clk_in scanchain_179/clk_in scanchain_178/data_in scanchain_179/data_in
+ scanchain_178/latch_enable_in scanchain_179/latch_enable_in scanchain_178/module_data_in[0]
+ scanchain_178/module_data_in[1] scanchain_178/module_data_in[2] scanchain_178/module_data_in[3]
+ scanchain_178/module_data_in[4] scanchain_178/module_data_in[5] scanchain_178/module_data_in[6]
+ scanchain_178/module_data_in[7] scanchain_178/module_data_out[0] scanchain_178/module_data_out[1]
+ scanchain_178/module_data_out[2] scanchain_178/module_data_out[3] scanchain_178/module_data_out[4]
+ scanchain_178/module_data_out[5] scanchain_178/module_data_out[6] scanchain_178/module_data_out[7]
+ scanchain_178/scan_select_in scanchain_179/scan_select_in vccd1 vssd1 scanchain
Xscanchain_156 scanchain_156/clk_in scanchain_157/clk_in scanchain_156/data_in scanchain_157/data_in
+ scanchain_156/latch_enable_in scanchain_157/latch_enable_in scanchain_156/module_data_in[0]
+ scanchain_156/module_data_in[1] scanchain_156/module_data_in[2] scanchain_156/module_data_in[3]
+ scanchain_156/module_data_in[4] scanchain_156/module_data_in[5] scanchain_156/module_data_in[6]
+ scanchain_156/module_data_in[7] scanchain_156/module_data_out[0] scanchain_156/module_data_out[1]
+ scanchain_156/module_data_out[2] scanchain_156/module_data_out[3] scanchain_156/module_data_out[4]
+ scanchain_156/module_data_out[5] scanchain_156/module_data_out[6] scanchain_156/module_data_out[7]
+ scanchain_156/scan_select_in scanchain_157/scan_select_in vccd1 vssd1 scanchain
Xuser_module_360014965627378689_020 scanchain_020/module_data_in[0] scanchain_020/module_data_in[1]
+ scanchain_020/module_data_in[2] scanchain_020/module_data_in[3] scanchain_020/module_data_in[4]
+ scanchain_020/module_data_in[5] scanchain_020/module_data_in[6] scanchain_020/module_data_in[7]
+ scanchain_020/module_data_out[0] scanchain_020/module_data_out[1] scanchain_020/module_data_out[2]
+ scanchain_020/module_data_out[3] scanchain_020/module_data_out[4] scanchain_020/module_data_out[5]
+ scanchain_020/module_data_out[6] scanchain_020/module_data_out[7] vccd1 vssd1 user_module_360014965627378689
Xuser_module_361728533238569985_091 scanchain_091/module_data_in[0] scanchain_091/module_data_in[1]
+ scanchain_091/module_data_in[2] scanchain_091/module_data_in[3] scanchain_091/module_data_in[4]
+ scanchain_091/module_data_in[5] scanchain_091/module_data_in[6] scanchain_091/module_data_in[7]
+ scanchain_091/module_data_out[0] scanchain_091/module_data_out[1] scanchain_091/module_data_out[2]
+ scanchain_091/module_data_out[3] scanchain_091/module_data_out[4] scanchain_091/module_data_out[5]
+ scanchain_091/module_data_out[6] scanchain_091/module_data_out[7] vccd1 vssd1 user_module_361728533238569985
Xuser_module_357917324056483841_054 scanchain_054/module_data_in[0] scanchain_054/module_data_in[1]
+ scanchain_054/module_data_in[2] scanchain_054/module_data_in[3] scanchain_054/module_data_in[4]
+ scanchain_054/module_data_in[5] scanchain_054/module_data_in[6] scanchain_054/module_data_in[7]
+ scanchain_054/module_data_out[0] scanchain_054/module_data_out[1] scanchain_054/module_data_out[2]
+ scanchain_054/module_data_out[3] scanchain_054/module_data_out[4] scanchain_054/module_data_out[5]
+ scanchain_054/module_data_out[6] scanchain_054/module_data_out[7] vccd1 vssd1 user_module_357917324056483841
Xmoonbase_pdp8_019 moonbase_pdp8_019/io_in[0] moonbase_pdp8_019/io_in[1] moonbase_pdp8_019/io_in[2]
+ moonbase_pdp8_019/io_in[3] moonbase_pdp8_019/io_in[4] moonbase_pdp8_019/io_in[5]
+ moonbase_pdp8_019/io_in[6] moonbase_pdp8_019/io_in[7] moonbase_pdp8_019/io_out[0]
+ moonbase_pdp8_019/io_out[1] moonbase_pdp8_019/io_out[2] moonbase_pdp8_019/io_out[3]
+ moonbase_pdp8_019/io_out[4] moonbase_pdp8_019/io_out[5] moonbase_pdp8_019/io_out[6]
+ moonbase_pdp8_019/io_out[7] vccd1 vssd1 moonbase_pdp8
Xuser_module_359353377078748161_010 scanchain_010/module_data_in[0] scanchain_010/module_data_in[1]
+ scanchain_010/module_data_in[2] scanchain_010/module_data_in[3] scanchain_010/module_data_in[4]
+ scanchain_010/module_data_in[5] scanchain_010/module_data_in[6] scanchain_010/module_data_in[7]
+ scanchain_010/module_data_out[0] scanchain_010/module_data_out[1] scanchain_010/module_data_out[2]
+ scanchain_010/module_data_out[3] scanchain_010/module_data_out[4] scanchain_010/module_data_out[5]
+ scanchain_010/module_data_out[6] scanchain_010/module_data_out[7] vccd1 vssd1 user_module_359353377078748161
Xscanchain_124 scanchain_124/clk_in scanchain_125/clk_in scanchain_124/data_in scanchain_125/data_in
+ scanchain_124/latch_enable_in scanchain_125/latch_enable_in scanchain_124/module_data_in[0]
+ scanchain_124/module_data_in[1] scanchain_124/module_data_in[2] scanchain_124/module_data_in[3]
+ scanchain_124/module_data_in[4] scanchain_124/module_data_in[5] scanchain_124/module_data_in[6]
+ scanchain_124/module_data_in[7] scanchain_124/module_data_out[0] scanchain_124/module_data_out[1]
+ scanchain_124/module_data_out[2] scanchain_124/module_data_out[3] scanchain_124/module_data_out[4]
+ scanchain_124/module_data_out[5] scanchain_124/module_data_out[6] scanchain_124/module_data_out[7]
+ scanchain_124/scan_select_in scanchain_125/scan_select_in vccd1 vssd1 scanchain
Xscanchain_135 scanchain_135/clk_in scanchain_136/clk_in scanchain_135/data_in scanchain_136/data_in
+ scanchain_135/latch_enable_in scanchain_136/latch_enable_in scanchain_135/module_data_in[0]
+ scanchain_135/module_data_in[1] scanchain_135/module_data_in[2] scanchain_135/module_data_in[3]
+ scanchain_135/module_data_in[4] scanchain_135/module_data_in[5] scanchain_135/module_data_in[6]
+ scanchain_135/module_data_in[7] scanchain_135/module_data_out[0] scanchain_135/module_data_out[1]
+ scanchain_135/module_data_out[2] scanchain_135/module_data_out[3] scanchain_135/module_data_out[4]
+ scanchain_135/module_data_out[5] scanchain_135/module_data_out[6] scanchain_135/module_data_out[7]
+ scanchain_135/scan_select_in scanchain_136/scan_select_in vccd1 vssd1 scanchain
Xscanchain_113 scanchain_113/clk_in scanchain_114/clk_in scanchain_113/data_in scanchain_114/data_in
+ scanchain_113/latch_enable_in scanchain_114/latch_enable_in scanchain_113/module_data_in[0]
+ scanchain_113/module_data_in[1] scanchain_113/module_data_in[2] scanchain_113/module_data_in[3]
+ scanchain_113/module_data_in[4] scanchain_113/module_data_in[5] scanchain_113/module_data_in[6]
+ scanchain_113/module_data_in[7] scanchain_113/module_data_out[0] scanchain_113/module_data_out[1]
+ scanchain_113/module_data_out[2] scanchain_113/module_data_out[3] scanchain_113/module_data_out[4]
+ scanchain_113/module_data_out[5] scanchain_113/module_data_out[6] scanchain_113/module_data_out[7]
+ scanchain_113/scan_select_in scanchain_114/scan_select_in vccd1 vssd1 scanchain
Xscanchain_146 scanchain_146/clk_in scanchain_147/clk_in scanchain_146/data_in scanchain_147/data_in
+ scanchain_146/latch_enable_in scanchain_147/latch_enable_in scanchain_146/module_data_in[0]
+ scanchain_146/module_data_in[1] scanchain_146/module_data_in[2] scanchain_146/module_data_in[3]
+ scanchain_146/module_data_in[4] scanchain_146/module_data_in[5] scanchain_146/module_data_in[6]
+ scanchain_146/module_data_in[7] scanchain_146/module_data_out[0] scanchain_146/module_data_out[1]
+ scanchain_146/module_data_out[2] scanchain_146/module_data_out[3] scanchain_146/module_data_out[4]
+ scanchain_146/module_data_out[5] scanchain_146/module_data_out[6] scanchain_146/module_data_out[7]
+ scanchain_146/scan_select_in scanchain_147/scan_select_in vccd1 vssd1 scanchain
Xscanchain_102 scanchain_102/clk_in scanchain_103/clk_in scanchain_102/data_in scanchain_103/data_in
+ scanchain_102/latch_enable_in scanchain_103/latch_enable_in scanchain_102/module_data_in[0]
+ scanchain_102/module_data_in[1] scanchain_102/module_data_in[2] scanchain_102/module_data_in[3]
+ scanchain_102/module_data_in[4] scanchain_102/module_data_in[5] scanchain_102/module_data_in[6]
+ scanchain_102/module_data_in[7] scanchain_102/module_data_out[0] scanchain_102/module_data_out[1]
+ scanchain_102/module_data_out[2] scanchain_102/module_data_out[3] scanchain_102/module_data_out[4]
+ scanchain_102/module_data_out[5] scanchain_102/module_data_out[6] scanchain_102/module_data_out[7]
+ scanchain_102/scan_select_in scanchain_103/scan_select_in vccd1 vssd1 scanchain
Xuser_module_361728533238569985_240 scanchain_240/module_data_in[0] scanchain_240/module_data_in[1]
+ scanchain_240/module_data_in[2] scanchain_240/module_data_in[3] scanchain_240/module_data_in[4]
+ scanchain_240/module_data_in[5] scanchain_240/module_data_in[6] scanchain_240/module_data_in[7]
+ scanchain_240/module_data_out[0] scanchain_240/module_data_out[1] scanchain_240/module_data_out[2]
+ scanchain_240/module_data_out[3] scanchain_240/module_data_out[4] scanchain_240/module_data_out[5]
+ scanchain_240/module_data_out[6] scanchain_240/module_data_out[7] vccd1 vssd1 user_module_361728533238569985
Xscanchain_168 scanchain_168/clk_in scanchain_169/clk_in scanchain_168/data_in scanchain_169/data_in
+ scanchain_168/latch_enable_in scanchain_169/latch_enable_in scanchain_168/module_data_in[0]
+ scanchain_168/module_data_in[1] scanchain_168/module_data_in[2] scanchain_168/module_data_in[3]
+ scanchain_168/module_data_in[4] scanchain_168/module_data_in[5] scanchain_168/module_data_in[6]
+ scanchain_168/module_data_in[7] scanchain_168/module_data_out[0] scanchain_168/module_data_out[1]
+ scanchain_168/module_data_out[2] scanchain_168/module_data_out[3] scanchain_168/module_data_out[4]
+ scanchain_168/module_data_out[5] scanchain_168/module_data_out[6] scanchain_168/module_data_out[7]
+ scanchain_168/scan_select_in scanchain_169/scan_select_in vccd1 vssd1 scanchain
Xscanchain_179 scanchain_179/clk_in scanchain_180/clk_in scanchain_179/data_in scanchain_180/data_in
+ scanchain_179/latch_enable_in scanchain_180/latch_enable_in scanchain_179/module_data_in[0]
+ scanchain_179/module_data_in[1] scanchain_179/module_data_in[2] scanchain_179/module_data_in[3]
+ scanchain_179/module_data_in[4] scanchain_179/module_data_in[5] scanchain_179/module_data_in[6]
+ scanchain_179/module_data_in[7] scanchain_179/module_data_out[0] scanchain_179/module_data_out[1]
+ scanchain_179/module_data_out[2] scanchain_179/module_data_out[3] scanchain_179/module_data_out[4]
+ scanchain_179/module_data_out[5] scanchain_179/module_data_out[6] scanchain_179/module_data_out[7]
+ scanchain_179/scan_select_in scanchain_180/scan_select_in vccd1 vssd1 scanchain
Xscanchain_157 scanchain_157/clk_in scanchain_158/clk_in scanchain_157/data_in scanchain_158/data_in
+ scanchain_157/latch_enable_in scanchain_158/latch_enable_in scanchain_157/module_data_in[0]
+ scanchain_157/module_data_in[1] scanchain_157/module_data_in[2] scanchain_157/module_data_in[3]
+ scanchain_157/module_data_in[4] scanchain_157/module_data_in[5] scanchain_157/module_data_in[6]
+ scanchain_157/module_data_in[7] scanchain_157/module_data_out[0] scanchain_157/module_data_out[1]
+ scanchain_157/module_data_out[2] scanchain_157/module_data_out[3] scanchain_157/module_data_out[4]
+ scanchain_157/module_data_out[5] scanchain_157/module_data_out[6] scanchain_157/module_data_out[7]
+ scanchain_157/scan_select_in scanchain_158/scan_select_in vccd1 vssd1 scanchain
Xuser_module_361728533238569985_092 scanchain_092/module_data_in[0] scanchain_092/module_data_in[1]
+ scanchain_092/module_data_in[2] scanchain_092/module_data_in[3] scanchain_092/module_data_in[4]
+ scanchain_092/module_data_in[5] scanchain_092/module_data_in[6] scanchain_092/module_data_in[7]
+ scanchain_092/module_data_out[0] scanchain_092/module_data_out[1] scanchain_092/module_data_out[2]
+ scanchain_092/module_data_out[3] scanchain_092/module_data_out[4] scanchain_092/module_data_out[5]
+ scanchain_092/module_data_out[6] scanchain_092/module_data_out[7] vccd1 vssd1 user_module_361728533238569985
XBenAtUvu_combo_058 BenAtUvu_combo_058/io_in[0] BenAtUvu_combo_058/io_in[1] BenAtUvu_combo_058/io_in[2]
+ BenAtUvu_combo_058/io_in[3] BenAtUvu_combo_058/io_in[4] BenAtUvu_combo_058/io_in[5]
+ BenAtUvu_combo_058/io_in[6] BenAtUvu_combo_058/io_in[7] BenAtUvu_combo_058/io_out[0]
+ BenAtUvu_combo_058/io_out[1] BenAtUvu_combo_058/io_out[2] BenAtUvu_combo_058/io_out[3]
+ BenAtUvu_combo_058/io_out[4] BenAtUvu_combo_058/io_out[5] BenAtUvu_combo_058/io_out[6]
+ BenAtUvu_combo_058/io_out[7] vccd1 vssd1 BenAtUvu_combo
Xscanchain_125 scanchain_125/clk_in scanchain_126/clk_in scanchain_125/data_in scanchain_126/data_in
+ scanchain_125/latch_enable_in scanchain_126/latch_enable_in scanchain_125/module_data_in[0]
+ scanchain_125/module_data_in[1] scanchain_125/module_data_in[2] scanchain_125/module_data_in[3]
+ scanchain_125/module_data_in[4] scanchain_125/module_data_in[5] scanchain_125/module_data_in[6]
+ scanchain_125/module_data_in[7] scanchain_125/module_data_out[0] scanchain_125/module_data_out[1]
+ scanchain_125/module_data_out[2] scanchain_125/module_data_out[3] scanchain_125/module_data_out[4]
+ scanchain_125/module_data_out[5] scanchain_125/module_data_out[6] scanchain_125/module_data_out[7]
+ scanchain_125/scan_select_in scanchain_126/scan_select_in vccd1 vssd1 scanchain
Xscanchain_136 scanchain_136/clk_in scanchain_137/clk_in scanchain_136/data_in scanchain_137/data_in
+ scanchain_136/latch_enable_in scanchain_137/latch_enable_in scanchain_136/module_data_in[0]
+ scanchain_136/module_data_in[1] scanchain_136/module_data_in[2] scanchain_136/module_data_in[3]
+ scanchain_136/module_data_in[4] scanchain_136/module_data_in[5] scanchain_136/module_data_in[6]
+ scanchain_136/module_data_in[7] scanchain_136/module_data_out[0] scanchain_136/module_data_out[1]
+ scanchain_136/module_data_out[2] scanchain_136/module_data_out[3] scanchain_136/module_data_out[4]
+ scanchain_136/module_data_out[5] scanchain_136/module_data_out[6] scanchain_136/module_data_out[7]
+ scanchain_136/scan_select_in scanchain_137/scan_select_in vccd1 vssd1 scanchain
Xscanchain_114 scanchain_114/clk_in scanchain_115/clk_in scanchain_114/data_in scanchain_115/data_in
+ scanchain_114/latch_enable_in scanchain_115/latch_enable_in scanchain_114/module_data_in[0]
+ scanchain_114/module_data_in[1] scanchain_114/module_data_in[2] scanchain_114/module_data_in[3]
+ scanchain_114/module_data_in[4] scanchain_114/module_data_in[5] scanchain_114/module_data_in[6]
+ scanchain_114/module_data_in[7] scanchain_114/module_data_out[0] scanchain_114/module_data_out[1]
+ scanchain_114/module_data_out[2] scanchain_114/module_data_out[3] scanchain_114/module_data_out[4]
+ scanchain_114/module_data_out[5] scanchain_114/module_data_out[6] scanchain_114/module_data_out[7]
+ scanchain_114/scan_select_in scanchain_115/scan_select_in vccd1 vssd1 scanchain
Xscanchain_147 scanchain_147/clk_in scanchain_148/clk_in scanchain_147/data_in scanchain_148/data_in
+ scanchain_147/latch_enable_in scanchain_148/latch_enable_in scanchain_147/module_data_in[0]
+ scanchain_147/module_data_in[1] scanchain_147/module_data_in[2] scanchain_147/module_data_in[3]
+ scanchain_147/module_data_in[4] scanchain_147/module_data_in[5] scanchain_147/module_data_in[6]
+ scanchain_147/module_data_in[7] scanchain_147/module_data_out[0] scanchain_147/module_data_out[1]
+ scanchain_147/module_data_out[2] scanchain_147/module_data_out[3] scanchain_147/module_data_out[4]
+ scanchain_147/module_data_out[5] scanchain_147/module_data_out[6] scanchain_147/module_data_out[7]
+ scanchain_147/scan_select_in scanchain_148/scan_select_in vccd1 vssd1 scanchain
Xscanchain_103 scanchain_103/clk_in scanchain_104/clk_in scanchain_103/data_in scanchain_104/data_in
+ scanchain_103/latch_enable_in scanchain_104/latch_enable_in scanchain_103/module_data_in[0]
+ scanchain_103/module_data_in[1] scanchain_103/module_data_in[2] scanchain_103/module_data_in[3]
+ scanchain_103/module_data_in[4] scanchain_103/module_data_in[5] scanchain_103/module_data_in[6]
+ scanchain_103/module_data_in[7] scanchain_103/module_data_out[0] scanchain_103/module_data_out[1]
+ scanchain_103/module_data_out[2] scanchain_103/module_data_out[3] scanchain_103/module_data_out[4]
+ scanchain_103/module_data_out[5] scanchain_103/module_data_out[6] scanchain_103/module_data_out[7]
+ scanchain_103/scan_select_in scanchain_104/scan_select_in vccd1 vssd1 scanchain
Xuser_module_361728533238569985_230 scanchain_230/module_data_in[0] scanchain_230/module_data_in[1]
+ scanchain_230/module_data_in[2] scanchain_230/module_data_in[3] scanchain_230/module_data_in[4]
+ scanchain_230/module_data_in[5] scanchain_230/module_data_in[6] scanchain_230/module_data_in[7]
+ scanchain_230/module_data_out[0] scanchain_230/module_data_out[1] scanchain_230/module_data_out[2]
+ scanchain_230/module_data_out[3] scanchain_230/module_data_out[4] scanchain_230/module_data_out[5]
+ scanchain_230/module_data_out[6] scanchain_230/module_data_out[7] vccd1 vssd1 user_module_361728533238569985
Xuser_module_361728533238569985_241 scanchain_241/module_data_in[0] scanchain_241/module_data_in[1]
+ scanchain_241/module_data_in[2] scanchain_241/module_data_in[3] scanchain_241/module_data_in[4]
+ scanchain_241/module_data_in[5] scanchain_241/module_data_in[6] scanchain_241/module_data_in[7]
+ scanchain_241/module_data_out[0] scanchain_241/module_data_out[1] scanchain_241/module_data_out[2]
+ scanchain_241/module_data_out[3] scanchain_241/module_data_out[4] scanchain_241/module_data_out[5]
+ scanchain_241/module_data_out[6] scanchain_241/module_data_out[7] vccd1 vssd1 user_module_361728533238569985
Xscanchain_169 scanchain_169/clk_in scanchain_170/clk_in scanchain_169/data_in scanchain_170/data_in
+ scanchain_169/latch_enable_in scanchain_170/latch_enable_in scanchain_169/module_data_in[0]
+ scanchain_169/module_data_in[1] scanchain_169/module_data_in[2] scanchain_169/module_data_in[3]
+ scanchain_169/module_data_in[4] scanchain_169/module_data_in[5] scanchain_169/module_data_in[6]
+ scanchain_169/module_data_in[7] scanchain_169/module_data_out[0] scanchain_169/module_data_out[1]
+ scanchain_169/module_data_out[2] scanchain_169/module_data_out[3] scanchain_169/module_data_out[4]
+ scanchain_169/module_data_out[5] scanchain_169/module_data_out[6] scanchain_169/module_data_out[7]
+ scanchain_169/scan_select_in scanchain_170/scan_select_in vccd1 vssd1 scanchain
Xscanchain_158 scanchain_158/clk_in scanchain_159/clk_in scanchain_158/data_in scanchain_159/data_in
+ scanchain_158/latch_enable_in scanchain_159/latch_enable_in scanchain_158/module_data_in[0]
+ scanchain_158/module_data_in[1] scanchain_158/module_data_in[2] scanchain_158/module_data_in[3]
+ scanchain_158/module_data_in[4] scanchain_158/module_data_in[5] scanchain_158/module_data_in[6]
+ scanchain_158/module_data_in[7] scanchain_158/module_data_out[0] scanchain_158/module_data_out[1]
+ scanchain_158/module_data_out[2] scanchain_158/module_data_out[3] scanchain_158/module_data_out[4]
+ scanchain_158/module_data_out[5] scanchain_158/module_data_out[6] scanchain_158/module_data_out[7]
+ scanchain_158/scan_select_in scanchain_159/scan_select_in vccd1 vssd1 scanchain
Xuser_module_361728533238569985_093 scanchain_093/module_data_in[0] scanchain_093/module_data_in[1]
+ scanchain_093/module_data_in[2] scanchain_093/module_data_in[3] scanchain_093/module_data_in[4]
+ scanchain_093/module_data_in[5] scanchain_093/module_data_in[6] scanchain_093/module_data_in[7]
+ scanchain_093/module_data_out[0] scanchain_093/module_data_out[1] scanchain_093/module_data_out[2]
+ scanchain_093/module_data_out[3] scanchain_093/module_data_out[4] scanchain_093/module_data_out[5]
+ scanchain_093/module_data_out[6] scanchain_093/module_data_out[7] vccd1 vssd1 user_module_361728533238569985
Xscanchain_126 scanchain_126/clk_in scanchain_127/clk_in scanchain_126/data_in scanchain_127/data_in
+ scanchain_126/latch_enable_in scanchain_127/latch_enable_in scanchain_126/module_data_in[0]
+ scanchain_126/module_data_in[1] scanchain_126/module_data_in[2] scanchain_126/module_data_in[3]
+ scanchain_126/module_data_in[4] scanchain_126/module_data_in[5] scanchain_126/module_data_in[6]
+ scanchain_126/module_data_in[7] scanchain_126/module_data_out[0] scanchain_126/module_data_out[1]
+ scanchain_126/module_data_out[2] scanchain_126/module_data_out[3] scanchain_126/module_data_out[4]
+ scanchain_126/module_data_out[5] scanchain_126/module_data_out[6] scanchain_126/module_data_out[7]
+ scanchain_126/scan_select_in scanchain_127/scan_select_in vccd1 vssd1 scanchain
Xscanchain_115 scanchain_115/clk_in scanchain_116/clk_in scanchain_115/data_in scanchain_116/data_in
+ scanchain_115/latch_enable_in scanchain_116/latch_enable_in scanchain_115/module_data_in[0]
+ scanchain_115/module_data_in[1] scanchain_115/module_data_in[2] scanchain_115/module_data_in[3]
+ scanchain_115/module_data_in[4] scanchain_115/module_data_in[5] scanchain_115/module_data_in[6]
+ scanchain_115/module_data_in[7] scanchain_115/module_data_out[0] scanchain_115/module_data_out[1]
+ scanchain_115/module_data_out[2] scanchain_115/module_data_out[3] scanchain_115/module_data_out[4]
+ scanchain_115/module_data_out[5] scanchain_115/module_data_out[6] scanchain_115/module_data_out[7]
+ scanchain_115/scan_select_in scanchain_116/scan_select_in vccd1 vssd1 scanchain
Xscanchain_137 scanchain_137/clk_in scanchain_138/clk_in scanchain_137/data_in scanchain_138/data_in
+ scanchain_137/latch_enable_in scanchain_138/latch_enable_in scanchain_137/module_data_in[0]
+ scanchain_137/module_data_in[1] scanchain_137/module_data_in[2] scanchain_137/module_data_in[3]
+ scanchain_137/module_data_in[4] scanchain_137/module_data_in[5] scanchain_137/module_data_in[6]
+ scanchain_137/module_data_in[7] scanchain_137/module_data_out[0] scanchain_137/module_data_out[1]
+ scanchain_137/module_data_out[2] scanchain_137/module_data_out[3] scanchain_137/module_data_out[4]
+ scanchain_137/module_data_out[5] scanchain_137/module_data_out[6] scanchain_137/module_data_out[7]
+ scanchain_137/scan_select_in scanchain_138/scan_select_in vccd1 vssd1 scanchain
Xscanchain_104 scanchain_104/clk_in scanchain_105/clk_in scanchain_104/data_in scanchain_105/data_in
+ scanchain_104/latch_enable_in scanchain_105/latch_enable_in scanchain_104/module_data_in[0]
+ scanchain_104/module_data_in[1] scanchain_104/module_data_in[2] scanchain_104/module_data_in[3]
+ scanchain_104/module_data_in[4] scanchain_104/module_data_in[5] scanchain_104/module_data_in[6]
+ scanchain_104/module_data_in[7] scanchain_104/module_data_out[0] scanchain_104/module_data_out[1]
+ scanchain_104/module_data_out[2] scanchain_104/module_data_out[3] scanchain_104/module_data_out[4]
+ scanchain_104/module_data_out[5] scanchain_104/module_data_out[6] scanchain_104/module_data_out[7]
+ scanchain_104/scan_select_in scanchain_105/scan_select_in vccd1 vssd1 scanchain
Xscanchain_148 scanchain_148/clk_in scanchain_149/clk_in scanchain_148/data_in scanchain_149/data_in
+ scanchain_148/latch_enable_in scanchain_149/latch_enable_in scanchain_148/module_data_in[0]
+ scanchain_148/module_data_in[1] scanchain_148/module_data_in[2] scanchain_148/module_data_in[3]
+ scanchain_148/module_data_in[4] scanchain_148/module_data_in[5] scanchain_148/module_data_in[6]
+ scanchain_148/module_data_in[7] scanchain_148/module_data_out[0] scanchain_148/module_data_out[1]
+ scanchain_148/module_data_out[2] scanchain_148/module_data_out[3] scanchain_148/module_data_out[4]
+ scanchain_148/module_data_out[5] scanchain_148/module_data_out[6] scanchain_148/module_data_out[7]
+ scanchain_148/scan_select_in scanchain_149/scan_select_in vccd1 vssd1 scanchain
Xscanchain_159 scanchain_159/clk_in scanchain_160/clk_in scanchain_159/data_in scanchain_160/data_in
+ scanchain_159/latch_enable_in scanchain_160/latch_enable_in scanchain_159/module_data_in[0]
+ scanchain_159/module_data_in[1] scanchain_159/module_data_in[2] scanchain_159/module_data_in[3]
+ scanchain_159/module_data_in[4] scanchain_159/module_data_in[5] scanchain_159/module_data_in[6]
+ scanchain_159/module_data_in[7] scanchain_159/module_data_out[0] scanchain_159/module_data_out[1]
+ scanchain_159/module_data_out[2] scanchain_159/module_data_out[3] scanchain_159/module_data_out[4]
+ scanchain_159/module_data_out[5] scanchain_159/module_data_out[6] scanchain_159/module_data_out[7]
+ scanchain_159/scan_select_in scanchain_160/scan_select_in vccd1 vssd1 scanchain
Xuser_module_361728533238569985_231 scanchain_231/module_data_in[0] scanchain_231/module_data_in[1]
+ scanchain_231/module_data_in[2] scanchain_231/module_data_in[3] scanchain_231/module_data_in[4]
+ scanchain_231/module_data_in[5] scanchain_231/module_data_in[6] scanchain_231/module_data_in[7]
+ scanchain_231/module_data_out[0] scanchain_231/module_data_out[1] scanchain_231/module_data_out[2]
+ scanchain_231/module_data_out[3] scanchain_231/module_data_out[4] scanchain_231/module_data_out[5]
+ scanchain_231/module_data_out[6] scanchain_231/module_data_out[7] vccd1 vssd1 user_module_361728533238569985
Xuser_module_361728533238569985_242 scanchain_242/module_data_in[0] scanchain_242/module_data_in[1]
+ scanchain_242/module_data_in[2] scanchain_242/module_data_in[3] scanchain_242/module_data_in[4]
+ scanchain_242/module_data_in[5] scanchain_242/module_data_in[6] scanchain_242/module_data_in[7]
+ scanchain_242/module_data_out[0] scanchain_242/module_data_out[1] scanchain_242/module_data_out[2]
+ scanchain_242/module_data_out[3] scanchain_242/module_data_out[4] scanchain_242/module_data_out[5]
+ scanchain_242/module_data_out[6] scanchain_242/module_data_out[7] vccd1 vssd1 user_module_361728533238569985
Xuser_module_361728533238569985_220 scanchain_220/module_data_in[0] scanchain_220/module_data_in[1]
+ scanchain_220/module_data_in[2] scanchain_220/module_data_in[3] scanchain_220/module_data_in[4]
+ scanchain_220/module_data_in[5] scanchain_220/module_data_in[6] scanchain_220/module_data_in[7]
+ scanchain_220/module_data_out[0] scanchain_220/module_data_out[1] scanchain_220/module_data_out[2]
+ scanchain_220/module_data_out[3] scanchain_220/module_data_out[4] scanchain_220/module_data_out[5]
+ scanchain_220/module_data_out[6] scanchain_220/module_data_out[7] vccd1 vssd1 user_module_361728533238569985
Xuser_module_361728533238569985_094 scanchain_094/module_data_in[0] scanchain_094/module_data_in[1]
+ scanchain_094/module_data_in[2] scanchain_094/module_data_in[3] scanchain_094/module_data_in[4]
+ scanchain_094/module_data_in[5] scanchain_094/module_data_in[6] scanchain_094/module_data_in[7]
+ scanchain_094/module_data_out[0] scanchain_094/module_data_out[1] scanchain_094/module_data_out[2]
+ scanchain_094/module_data_out[3] scanchain_094/module_data_out[4] scanchain_094/module_data_out[5]
+ scanchain_094/module_data_out[6] scanchain_094/module_data_out[7] vccd1 vssd1 user_module_361728533238569985
Xuser_module_359372419264319489_014 scanchain_014/module_data_in[0] scanchain_014/module_data_in[1]
+ scanchain_014/module_data_in[2] scanchain_014/module_data_in[3] scanchain_014/module_data_in[4]
+ scanchain_014/module_data_in[5] scanchain_014/module_data_in[6] scanchain_014/module_data_in[7]
+ scanchain_014/module_data_out[0] scanchain_014/module_data_out[1] scanchain_014/module_data_out[2]
+ scanchain_014/module_data_out[3] scanchain_014/module_data_out[4] scanchain_014/module_data_out[5]
+ scanchain_014/module_data_out[6] scanchain_014/module_data_out[7] vccd1 vssd1 user_module_359372419264319489
Xdwisehart_top_043 dwisehart_top_043/io_in[0] dwisehart_top_043/io_in[1] dwisehart_top_043/io_in[2]
+ dwisehart_top_043/io_in[3] dwisehart_top_043/io_in[4] dwisehart_top_043/io_in[5]
+ dwisehart_top_043/io_in[6] dwisehart_top_043/io_in[7] dwisehart_top_043/io_out[0]
+ dwisehart_top_043/io_out[1] dwisehart_top_043/io_out[2] dwisehart_top_043/io_out[3]
+ dwisehart_top_043/io_out[4] dwisehart_top_043/io_out[5] dwisehart_top_043/io_out[6]
+ dwisehart_top_043/io_out[7] vccd1 vssd1 dwisehart_top
Xscanchain_127 scanchain_127/clk_in scanchain_128/clk_in scanchain_127/data_in scanchain_128/data_in
+ scanchain_127/latch_enable_in scanchain_128/latch_enable_in scanchain_127/module_data_in[0]
+ scanchain_127/module_data_in[1] scanchain_127/module_data_in[2] scanchain_127/module_data_in[3]
+ scanchain_127/module_data_in[4] scanchain_127/module_data_in[5] scanchain_127/module_data_in[6]
+ scanchain_127/module_data_in[7] scanchain_127/module_data_out[0] scanchain_127/module_data_out[1]
+ scanchain_127/module_data_out[2] scanchain_127/module_data_out[3] scanchain_127/module_data_out[4]
+ scanchain_127/module_data_out[5] scanchain_127/module_data_out[6] scanchain_127/module_data_out[7]
+ scanchain_127/scan_select_in scanchain_128/scan_select_in vccd1 vssd1 scanchain
Xscanchain_116 scanchain_116/clk_in scanchain_117/clk_in scanchain_116/data_in scanchain_117/data_in
+ scanchain_116/latch_enable_in scanchain_117/latch_enable_in scanchain_116/module_data_in[0]
+ scanchain_116/module_data_in[1] scanchain_116/module_data_in[2] scanchain_116/module_data_in[3]
+ scanchain_116/module_data_in[4] scanchain_116/module_data_in[5] scanchain_116/module_data_in[6]
+ scanchain_116/module_data_in[7] scanchain_116/module_data_out[0] scanchain_116/module_data_out[1]
+ scanchain_116/module_data_out[2] scanchain_116/module_data_out[3] scanchain_116/module_data_out[4]
+ scanchain_116/module_data_out[5] scanchain_116/module_data_out[6] scanchain_116/module_data_out[7]
+ scanchain_116/scan_select_in scanchain_117/scan_select_in vccd1 vssd1 scanchain
Xscanchain_138 scanchain_138/clk_in scanchain_139/clk_in scanchain_138/data_in scanchain_139/data_in
+ scanchain_138/latch_enable_in scanchain_139/latch_enable_in scanchain_138/module_data_in[0]
+ scanchain_138/module_data_in[1] scanchain_138/module_data_in[2] scanchain_138/module_data_in[3]
+ scanchain_138/module_data_in[4] scanchain_138/module_data_in[5] scanchain_138/module_data_in[6]
+ scanchain_138/module_data_in[7] scanchain_138/module_data_out[0] scanchain_138/module_data_out[1]
+ scanchain_138/module_data_out[2] scanchain_138/module_data_out[3] scanchain_138/module_data_out[4]
+ scanchain_138/module_data_out[5] scanchain_138/module_data_out[6] scanchain_138/module_data_out[7]
+ scanchain_138/scan_select_in scanchain_139/scan_select_in vccd1 vssd1 scanchain
Xscanchain_105 scanchain_105/clk_in scanchain_106/clk_in scanchain_105/data_in scanchain_106/data_in
+ scanchain_105/latch_enable_in scanchain_106/latch_enable_in scanchain_105/module_data_in[0]
+ scanchain_105/module_data_in[1] scanchain_105/module_data_in[2] scanchain_105/module_data_in[3]
+ scanchain_105/module_data_in[4] scanchain_105/module_data_in[5] scanchain_105/module_data_in[6]
+ scanchain_105/module_data_in[7] scanchain_105/module_data_out[0] scanchain_105/module_data_out[1]
+ scanchain_105/module_data_out[2] scanchain_105/module_data_out[3] scanchain_105/module_data_out[4]
+ scanchain_105/module_data_out[5] scanchain_105/module_data_out[6] scanchain_105/module_data_out[7]
+ scanchain_105/scan_select_in scanchain_106/scan_select_in vccd1 vssd1 scanchain
Xscanchain_149 scanchain_149/clk_in scanchain_150/clk_in scanchain_149/data_in scanchain_150/data_in
+ scanchain_149/latch_enable_in scanchain_150/latch_enable_in scanchain_149/module_data_in[0]
+ scanchain_149/module_data_in[1] scanchain_149/module_data_in[2] scanchain_149/module_data_in[3]
+ scanchain_149/module_data_in[4] scanchain_149/module_data_in[5] scanchain_149/module_data_in[6]
+ scanchain_149/module_data_in[7] scanchain_149/module_data_out[0] scanchain_149/module_data_out[1]
+ scanchain_149/module_data_out[2] scanchain_149/module_data_out[3] scanchain_149/module_data_out[4]
+ scanchain_149/module_data_out[5] scanchain_149/module_data_out[6] scanchain_149/module_data_out[7]
+ scanchain_149/scan_select_in scanchain_150/scan_select_in vccd1 vssd1 scanchain
Xuser_module_361728533238569985_232 scanchain_232/module_data_in[0] scanchain_232/module_data_in[1]
+ scanchain_232/module_data_in[2] scanchain_232/module_data_in[3] scanchain_232/module_data_in[4]
+ scanchain_232/module_data_in[5] scanchain_232/module_data_in[6] scanchain_232/module_data_in[7]
+ scanchain_232/module_data_out[0] scanchain_232/module_data_out[1] scanchain_232/module_data_out[2]
+ scanchain_232/module_data_out[3] scanchain_232/module_data_out[4] scanchain_232/module_data_out[5]
+ scanchain_232/module_data_out[6] scanchain_232/module_data_out[7] vccd1 vssd1 user_module_361728533238569985
Xuser_module_361728533238569985_243 scanchain_243/module_data_in[0] scanchain_243/module_data_in[1]
+ scanchain_243/module_data_in[2] scanchain_243/module_data_in[3] scanchain_243/module_data_in[4]
+ scanchain_243/module_data_in[5] scanchain_243/module_data_in[6] scanchain_243/module_data_in[7]
+ scanchain_243/module_data_out[0] scanchain_243/module_data_out[1] scanchain_243/module_data_out[2]
+ scanchain_243/module_data_out[3] scanchain_243/module_data_out[4] scanchain_243/module_data_out[5]
+ scanchain_243/module_data_out[6] scanchain_243/module_data_out[7] vccd1 vssd1 user_module_361728533238569985
Xuser_module_361728533238569985_221 scanchain_221/module_data_in[0] scanchain_221/module_data_in[1]
+ scanchain_221/module_data_in[2] scanchain_221/module_data_in[3] scanchain_221/module_data_in[4]
+ scanchain_221/module_data_in[5] scanchain_221/module_data_in[6] scanchain_221/module_data_in[7]
+ scanchain_221/module_data_out[0] scanchain_221/module_data_out[1] scanchain_221/module_data_out[2]
+ scanchain_221/module_data_out[3] scanchain_221/module_data_out[4] scanchain_221/module_data_out[5]
+ scanchain_221/module_data_out[6] scanchain_221/module_data_out[7] vccd1 vssd1 user_module_361728533238569985
Xuser_module_361728533238569985_210 scanchain_210/module_data_in[0] scanchain_210/module_data_in[1]
+ scanchain_210/module_data_in[2] scanchain_210/module_data_in[3] scanchain_210/module_data_in[4]
+ scanchain_210/module_data_in[5] scanchain_210/module_data_in[6] scanchain_210/module_data_in[7]
+ scanchain_210/module_data_out[0] scanchain_210/module_data_out[1] scanchain_210/module_data_out[2]
+ scanchain_210/module_data_out[3] scanchain_210/module_data_out[4] scanchain_210/module_data_out[5]
+ scanchain_210/module_data_out[6] scanchain_210/module_data_out[7] vccd1 vssd1 user_module_361728533238569985
Xuser_module_361728533238569985_040 scanchain_040/module_data_in[0] scanchain_040/module_data_in[1]
+ scanchain_040/module_data_in[2] scanchain_040/module_data_in[3] scanchain_040/module_data_in[4]
+ scanchain_040/module_data_in[5] scanchain_040/module_data_in[6] scanchain_040/module_data_in[7]
+ scanchain_040/module_data_out[0] scanchain_040/module_data_out[1] scanchain_040/module_data_out[2]
+ scanchain_040/module_data_out[3] scanchain_040/module_data_out[4] scanchain_040/module_data_out[5]
+ scanchain_040/module_data_out[6] scanchain_040/module_data_out[7] vccd1 vssd1 user_module_361728533238569985
Xuser_module_361728533238569985_095 scanchain_095/module_data_in[0] scanchain_095/module_data_in[1]
+ scanchain_095/module_data_in[2] scanchain_095/module_data_in[3] scanchain_095/module_data_in[4]
+ scanchain_095/module_data_in[5] scanchain_095/module_data_in[6] scanchain_095/module_data_in[7]
+ scanchain_095/module_data_out[0] scanchain_095/module_data_out[1] scanchain_095/module_data_out[2]
+ scanchain_095/module_data_out[3] scanchain_095/module_data_out[4] scanchain_095/module_data_out[5]
+ scanchain_095/module_data_out[6] scanchain_095/module_data_out[7] vccd1 vssd1 user_module_361728533238569985
Xuser_module_362336485347742721_080 scanchain_080/module_data_in[0] scanchain_080/module_data_in[1]
+ scanchain_080/module_data_in[2] scanchain_080/module_data_in[3] scanchain_080/module_data_in[4]
+ scanchain_080/module_data_in[5] scanchain_080/module_data_in[6] scanchain_080/module_data_in[7]
+ scanchain_080/module_data_out[0] scanchain_080/module_data_out[1] scanchain_080/module_data_out[2]
+ scanchain_080/module_data_out[3] scanchain_080/module_data_out[4] scanchain_080/module_data_out[5]
+ scanchain_080/module_data_out[6] scanchain_080/module_data_out[7] vccd1 vssd1 user_module_362336485347742721
Xkevinwguan_tiny_tapeout_061 scanchain_061/module_data_in[0] scanchain_061/module_data_in[1]
+ scanchain_061/module_data_in[2] scanchain_061/module_data_in[3] scanchain_061/module_data_in[4]
+ scanchain_061/module_data_in[5] scanchain_061/module_data_in[6] scanchain_061/module_data_in[7]
+ scanchain_061/module_data_out[0] scanchain_061/module_data_out[1] scanchain_061/module_data_out[2]
+ scanchain_061/module_data_out[3] scanchain_061/module_data_out[4] scanchain_061/module_data_out[5]
+ scanchain_061/module_data_out[6] scanchain_061/module_data_out[7] vccd1 vssd1 kevinwguan_tiny_tapeout
Xuser_module_361728533238569985_233 scanchain_233/module_data_in[0] scanchain_233/module_data_in[1]
+ scanchain_233/module_data_in[2] scanchain_233/module_data_in[3] scanchain_233/module_data_in[4]
+ scanchain_233/module_data_in[5] scanchain_233/module_data_in[6] scanchain_233/module_data_in[7]
+ scanchain_233/module_data_out[0] scanchain_233/module_data_out[1] scanchain_233/module_data_out[2]
+ scanchain_233/module_data_out[3] scanchain_233/module_data_out[4] scanchain_233/module_data_out[5]
+ scanchain_233/module_data_out[6] scanchain_233/module_data_out[7] vccd1 vssd1 user_module_361728533238569985
Xuser_module_361728533238569985_244 scanchain_244/module_data_in[0] scanchain_244/module_data_in[1]
+ scanchain_244/module_data_in[2] scanchain_244/module_data_in[3] scanchain_244/module_data_in[4]
+ scanchain_244/module_data_in[5] scanchain_244/module_data_in[6] scanchain_244/module_data_in[7]
+ scanchain_244/module_data_out[0] scanchain_244/module_data_out[1] scanchain_244/module_data_out[2]
+ scanchain_244/module_data_out[3] scanchain_244/module_data_out[4] scanchain_244/module_data_out[5]
+ scanchain_244/module_data_out[6] scanchain_244/module_data_out[7] vccd1 vssd1 user_module_361728533238569985
Xuser_module_361728533238569985_222 scanchain_222/module_data_in[0] scanchain_222/module_data_in[1]
+ scanchain_222/module_data_in[2] scanchain_222/module_data_in[3] scanchain_222/module_data_in[4]
+ scanchain_222/module_data_in[5] scanchain_222/module_data_in[6] scanchain_222/module_data_in[7]
+ scanchain_222/module_data_out[0] scanchain_222/module_data_out[1] scanchain_222/module_data_out[2]
+ scanchain_222/module_data_out[3] scanchain_222/module_data_out[4] scanchain_222/module_data_out[5]
+ scanchain_222/module_data_out[6] scanchain_222/module_data_out[7] vccd1 vssd1 user_module_361728533238569985
Xuser_module_361728533238569985_211 scanchain_211/module_data_in[0] scanchain_211/module_data_in[1]
+ scanchain_211/module_data_in[2] scanchain_211/module_data_in[3] scanchain_211/module_data_in[4]
+ scanchain_211/module_data_in[5] scanchain_211/module_data_in[6] scanchain_211/module_data_in[7]
+ scanchain_211/module_data_out[0] scanchain_211/module_data_out[1] scanchain_211/module_data_out[2]
+ scanchain_211/module_data_out[3] scanchain_211/module_data_out[4] scanchain_211/module_data_out[5]
+ scanchain_211/module_data_out[6] scanchain_211/module_data_out[7] vccd1 vssd1 user_module_361728533238569985
Xuser_module_361728533238569985_200 scanchain_200/module_data_in[0] scanchain_200/module_data_in[1]
+ scanchain_200/module_data_in[2] scanchain_200/module_data_in[3] scanchain_200/module_data_in[4]
+ scanchain_200/module_data_in[5] scanchain_200/module_data_in[6] scanchain_200/module_data_in[7]
+ scanchain_200/module_data_out[0] scanchain_200/module_data_out[1] scanchain_200/module_data_out[2]
+ scanchain_200/module_data_out[3] scanchain_200/module_data_out[4] scanchain_200/module_data_out[5]
+ scanchain_200/module_data_out[6] scanchain_200/module_data_out[7] vccd1 vssd1 user_module_361728533238569985
Xscanchain_128 scanchain_128/clk_in scanchain_129/clk_in scanchain_128/data_in scanchain_129/data_in
+ scanchain_128/latch_enable_in scanchain_129/latch_enable_in scanchain_128/module_data_in[0]
+ scanchain_128/module_data_in[1] scanchain_128/module_data_in[2] scanchain_128/module_data_in[3]
+ scanchain_128/module_data_in[4] scanchain_128/module_data_in[5] scanchain_128/module_data_in[6]
+ scanchain_128/module_data_in[7] scanchain_128/module_data_out[0] scanchain_128/module_data_out[1]
+ scanchain_128/module_data_out[2] scanchain_128/module_data_out[3] scanchain_128/module_data_out[4]
+ scanchain_128/module_data_out[5] scanchain_128/module_data_out[6] scanchain_128/module_data_out[7]
+ scanchain_128/scan_select_in scanchain_129/scan_select_in vccd1 vssd1 scanchain
Xscanchain_117 scanchain_117/clk_in scanchain_118/clk_in scanchain_117/data_in scanchain_118/data_in
+ scanchain_117/latch_enable_in scanchain_118/latch_enable_in scanchain_117/module_data_in[0]
+ scanchain_117/module_data_in[1] scanchain_117/module_data_in[2] scanchain_117/module_data_in[3]
+ scanchain_117/module_data_in[4] scanchain_117/module_data_in[5] scanchain_117/module_data_in[6]
+ scanchain_117/module_data_in[7] scanchain_117/module_data_out[0] scanchain_117/module_data_out[1]
+ scanchain_117/module_data_out[2] scanchain_117/module_data_out[3] scanchain_117/module_data_out[4]
+ scanchain_117/module_data_out[5] scanchain_117/module_data_out[6] scanchain_117/module_data_out[7]
+ scanchain_117/scan_select_in scanchain_118/scan_select_in vccd1 vssd1 scanchain
Xscanchain_106 scanchain_106/clk_in scanchain_107/clk_in scanchain_106/data_in scanchain_107/data_in
+ scanchain_106/latch_enable_in scanchain_107/latch_enable_in scanchain_106/module_data_in[0]
+ scanchain_106/module_data_in[1] scanchain_106/module_data_in[2] scanchain_106/module_data_in[3]
+ scanchain_106/module_data_in[4] scanchain_106/module_data_in[5] scanchain_106/module_data_in[6]
+ scanchain_106/module_data_in[7] scanchain_106/module_data_out[0] scanchain_106/module_data_out[1]
+ scanchain_106/module_data_out[2] scanchain_106/module_data_out[3] scanchain_106/module_data_out[4]
+ scanchain_106/module_data_out[5] scanchain_106/module_data_out[6] scanchain_106/module_data_out[7]
+ scanchain_106/scan_select_in scanchain_107/scan_select_in vccd1 vssd1 scanchain
Xscanchain_139 scanchain_139/clk_in scanchain_140/clk_in scanchain_139/data_in scanchain_140/data_in
+ scanchain_139/latch_enable_in scanchain_140/latch_enable_in scanchain_139/module_data_in[0]
+ scanchain_139/module_data_in[1] scanchain_139/module_data_in[2] scanchain_139/module_data_in[3]
+ scanchain_139/module_data_in[4] scanchain_139/module_data_in[5] scanchain_139/module_data_in[6]
+ scanchain_139/module_data_in[7] scanchain_139/module_data_out[0] scanchain_139/module_data_out[1]
+ scanchain_139/module_data_out[2] scanchain_139/module_data_out[3] scanchain_139/module_data_out[4]
+ scanchain_139/module_data_out[5] scanchain_139/module_data_out[6] scanchain_139/module_data_out[7]
+ scanchain_139/scan_select_in scanchain_140/scan_select_in vccd1 vssd1 scanchain
Xuser_module_361728533238569985_096 scanchain_096/module_data_in[0] scanchain_096/module_data_in[1]
+ scanchain_096/module_data_in[2] scanchain_096/module_data_in[3] scanchain_096/module_data_in[4]
+ scanchain_096/module_data_in[5] scanchain_096/module_data_in[6] scanchain_096/module_data_in[7]
+ scanchain_096/module_data_out[0] scanchain_096/module_data_out[1] scanchain_096/module_data_out[2]
+ scanchain_096/module_data_out[3] scanchain_096/module_data_out[4] scanchain_096/module_data_out[5]
+ scanchain_096/module_data_out[6] scanchain_096/module_data_out[7] vccd1 vssd1 user_module_361728533238569985
XMichaelBell_6bit_fifo_029 scanchain_029/module_data_in[0] scanchain_029/module_data_in[1]
+ scanchain_029/module_data_in[2] scanchain_029/module_data_in[3] scanchain_029/module_data_in[4]
+ scanchain_029/module_data_in[5] scanchain_029/module_data_in[6] scanchain_029/module_data_in[7]
+ scanchain_029/module_data_out[0] scanchain_029/module_data_out[1] scanchain_029/module_data_out[2]
+ scanchain_029/module_data_out[3] scanchain_029/module_data_out[4] scanchain_029/module_data_out[5]
+ scanchain_029/module_data_out[6] scanchain_029/module_data_out[7] vccd1 vssd1 MichaelBell_6bit_fifo
Xjblocklove_cgpt_benchmark_wrapper_064 scanchain_064/module_data_in[0] scanchain_064/module_data_in[1]
+ scanchain_064/module_data_in[2] scanchain_064/module_data_in[3] scanchain_064/module_data_in[4]
+ scanchain_064/module_data_in[5] scanchain_064/module_data_in[6] scanchain_064/module_data_in[7]
+ scanchain_064/module_data_out[0] scanchain_064/module_data_out[1] scanchain_064/module_data_out[2]
+ scanchain_064/module_data_out[3] scanchain_064/module_data_out[4] scanchain_064/module_data_out[5]
+ scanchain_064/module_data_out[6] scanchain_064/module_data_out[7] vccd1 vssd1 jblocklove_cgpt_benchmark_wrapper
Xuser_module_347497504164545108_088 scanchain_088/module_data_in[0] scanchain_088/module_data_in[1]
+ scanchain_088/module_data_in[2] scanchain_088/module_data_in[3] scanchain_088/module_data_in[4]
+ scanchain_088/module_data_in[5] scanchain_088/module_data_in[6] scanchain_088/module_data_in[7]
+ scanchain_088/module_data_out[0] scanchain_088/module_data_out[1] scanchain_088/module_data_out[2]
+ scanchain_088/module_data_out[3] scanchain_088/module_data_out[4] scanchain_088/module_data_out[5]
+ scanchain_088/module_data_out[6] scanchain_088/module_data_out[7] vccd1 vssd1 user_module_347497504164545108
Xscanchain_118 scanchain_118/clk_in scanchain_119/clk_in scanchain_118/data_in scanchain_119/data_in
+ scanchain_118/latch_enable_in scanchain_119/latch_enable_in scanchain_118/module_data_in[0]
+ scanchain_118/module_data_in[1] scanchain_118/module_data_in[2] scanchain_118/module_data_in[3]
+ scanchain_118/module_data_in[4] scanchain_118/module_data_in[5] scanchain_118/module_data_in[6]
+ scanchain_118/module_data_in[7] scanchain_118/module_data_out[0] scanchain_118/module_data_out[1]
+ scanchain_118/module_data_out[2] scanchain_118/module_data_out[3] scanchain_118/module_data_out[4]
+ scanchain_118/module_data_out[5] scanchain_118/module_data_out[6] scanchain_118/module_data_out[7]
+ scanchain_118/scan_select_in scanchain_119/scan_select_in vccd1 vssd1 scanchain
Xscanchain_129 scanchain_129/clk_in scanchain_130/clk_in scanchain_129/data_in scanchain_130/data_in
+ scanchain_129/latch_enable_in scanchain_130/latch_enable_in scanchain_129/module_data_in[0]
+ scanchain_129/module_data_in[1] scanchain_129/module_data_in[2] scanchain_129/module_data_in[3]
+ scanchain_129/module_data_in[4] scanchain_129/module_data_in[5] scanchain_129/module_data_in[6]
+ scanchain_129/module_data_in[7] scanchain_129/module_data_out[0] scanchain_129/module_data_out[1]
+ scanchain_129/module_data_out[2] scanchain_129/module_data_out[3] scanchain_129/module_data_out[4]
+ scanchain_129/module_data_out[5] scanchain_129/module_data_out[6] scanchain_129/module_data_out[7]
+ scanchain_129/scan_select_in scanchain_130/scan_select_in vccd1 vssd1 scanchain
Xscanchain_107 scanchain_107/clk_in scanchain_108/clk_in scanchain_107/data_in scanchain_108/data_in
+ scanchain_107/latch_enable_in scanchain_108/latch_enable_in scanchain_107/module_data_in[0]
+ scanchain_107/module_data_in[1] scanchain_107/module_data_in[2] scanchain_107/module_data_in[3]
+ scanchain_107/module_data_in[4] scanchain_107/module_data_in[5] scanchain_107/module_data_in[6]
+ scanchain_107/module_data_in[7] scanchain_107/module_data_out[0] scanchain_107/module_data_out[1]
+ scanchain_107/module_data_out[2] scanchain_107/module_data_out[3] scanchain_107/module_data_out[4]
+ scanchain_107/module_data_out[5] scanchain_107/module_data_out[6] scanchain_107/module_data_out[7]
+ scanchain_107/scan_select_in scanchain_108/scan_select_in vccd1 vssd1 scanchain
Xuser_module_361728533238569985_223 scanchain_223/module_data_in[0] scanchain_223/module_data_in[1]
+ scanchain_223/module_data_in[2] scanchain_223/module_data_in[3] scanchain_223/module_data_in[4]
+ scanchain_223/module_data_in[5] scanchain_223/module_data_in[6] scanchain_223/module_data_in[7]
+ scanchain_223/module_data_out[0] scanchain_223/module_data_out[1] scanchain_223/module_data_out[2]
+ scanchain_223/module_data_out[3] scanchain_223/module_data_out[4] scanchain_223/module_data_out[5]
+ scanchain_223/module_data_out[6] scanchain_223/module_data_out[7] vccd1 vssd1 user_module_361728533238569985
Xuser_module_361728533238569985_234 scanchain_234/module_data_in[0] scanchain_234/module_data_in[1]
+ scanchain_234/module_data_in[2] scanchain_234/module_data_in[3] scanchain_234/module_data_in[4]
+ scanchain_234/module_data_in[5] scanchain_234/module_data_in[6] scanchain_234/module_data_in[7]
+ scanchain_234/module_data_out[0] scanchain_234/module_data_out[1] scanchain_234/module_data_out[2]
+ scanchain_234/module_data_out[3] scanchain_234/module_data_out[4] scanchain_234/module_data_out[5]
+ scanchain_234/module_data_out[6] scanchain_234/module_data_out[7] vccd1 vssd1 user_module_361728533238569985
Xuser_module_361728533238569985_245 scanchain_245/module_data_in[0] scanchain_245/module_data_in[1]
+ scanchain_245/module_data_in[2] scanchain_245/module_data_in[3] scanchain_245/module_data_in[4]
+ scanchain_245/module_data_in[5] scanchain_245/module_data_in[6] scanchain_245/module_data_in[7]
+ scanchain_245/module_data_out[0] scanchain_245/module_data_out[1] scanchain_245/module_data_out[2]
+ scanchain_245/module_data_out[3] scanchain_245/module_data_out[4] scanchain_245/module_data_out[5]
+ scanchain_245/module_data_out[6] scanchain_245/module_data_out[7] vccd1 vssd1 user_module_361728533238569985
Xuser_module_361728533238569985_212 scanchain_212/module_data_in[0] scanchain_212/module_data_in[1]
+ scanchain_212/module_data_in[2] scanchain_212/module_data_in[3] scanchain_212/module_data_in[4]
+ scanchain_212/module_data_in[5] scanchain_212/module_data_in[6] scanchain_212/module_data_in[7]
+ scanchain_212/module_data_out[0] scanchain_212/module_data_out[1] scanchain_212/module_data_out[2]
+ scanchain_212/module_data_out[3] scanchain_212/module_data_out[4] scanchain_212/module_data_out[5]
+ scanchain_212/module_data_out[6] scanchain_212/module_data_out[7] vccd1 vssd1 user_module_361728533238569985
Xuser_module_361728533238569985_201 scanchain_201/module_data_in[0] scanchain_201/module_data_in[1]
+ scanchain_201/module_data_in[2] scanchain_201/module_data_in[3] scanchain_201/module_data_in[4]
+ scanchain_201/module_data_in[5] scanchain_201/module_data_in[6] scanchain_201/module_data_in[7]
+ scanchain_201/module_data_out[0] scanchain_201/module_data_out[1] scanchain_201/module_data_out[2]
+ scanchain_201/module_data_out[3] scanchain_201/module_data_out[4] scanchain_201/module_data_out[5]
+ scanchain_201/module_data_out[6] scanchain_201/module_data_out[7] vccd1 vssd1 user_module_361728533238569985
Xuser_module_361728533238569985_097 scanchain_097/module_data_in[0] scanchain_097/module_data_in[1]
+ scanchain_097/module_data_in[2] scanchain_097/module_data_in[3] scanchain_097/module_data_in[4]
+ scanchain_097/module_data_in[5] scanchain_097/module_data_in[6] scanchain_097/module_data_in[7]
+ scanchain_097/module_data_out[0] scanchain_097/module_data_out[1] scanchain_097/module_data_out[2]
+ scanchain_097/module_data_out[3] scanchain_097/module_data_out[4] scanchain_097/module_data_out[5]
+ scanchain_097/module_data_out[6] scanchain_097/module_data_out[7] vccd1 vssd1 user_module_361728533238569985
XMichaelBell_hovalaag_009 scanchain_009/module_data_in[0] scanchain_009/module_data_in[1]
+ scanchain_009/module_data_in[2] scanchain_009/module_data_in[3] scanchain_009/module_data_in[4]
+ scanchain_009/module_data_in[5] scanchain_009/module_data_in[6] scanchain_009/module_data_in[7]
+ scanchain_009/module_data_out[0] scanchain_009/module_data_out[1] scanchain_009/module_data_out[2]
+ scanchain_009/module_data_out[3] scanchain_009/module_data_out[4] scanchain_009/module_data_out[5]
+ scanchain_009/module_data_out[6] scanchain_009/module_data_out[7] vccd1 vssd1 MichaelBell_hovalaag
Xrobbertvanginkel_hamming74_068 scanchain_068/module_data_in[0] scanchain_068/module_data_in[1]
+ scanchain_068/module_data_in[2] scanchain_068/module_data_in[3] scanchain_068/module_data_in[4]
+ scanchain_068/module_data_in[5] scanchain_068/module_data_in[6] scanchain_068/module_data_in[7]
+ scanchain_068/module_data_out[0] scanchain_068/module_data_out[1] scanchain_068/module_data_out[2]
+ scanchain_068/module_data_out[3] scanchain_068/module_data_out[4] scanchain_068/module_data_out[5]
+ scanchain_068/module_data_out[6] scanchain_068/module_data_out[7] vccd1 vssd1 robbertvanginkel_hamming74
Xdratini0_fsk_modem_top_063 scanchain_063/module_data_in[0] scanchain_063/module_data_in[1]
+ scanchain_063/module_data_in[2] scanchain_063/module_data_in[3] scanchain_063/module_data_in[4]
+ scanchain_063/module_data_in[5] scanchain_063/module_data_in[6] scanchain_063/module_data_in[7]
+ scanchain_063/module_data_out[0] scanchain_063/module_data_out[1] scanchain_063/module_data_out[2]
+ scanchain_063/module_data_out[3] scanchain_063/module_data_out[4] scanchain_063/module_data_out[5]
+ scanchain_063/module_data_out[6] scanchain_063/module_data_out[7] vccd1 vssd1 dratini0_fsk_modem_top
Xshadow1229_player_016 shadow1229_player_016/io_in[0] shadow1229_player_016/io_in[1]
+ shadow1229_player_016/io_in[2] shadow1229_player_016/io_in[3] shadow1229_player_016/io_in[4]
+ shadow1229_player_016/io_in[5] shadow1229_player_016/io_in[6] shadow1229_player_016/io_in[7]
+ shadow1229_player_016/io_out[0] shadow1229_player_016/io_out[1] shadow1229_player_016/io_out[2]
+ shadow1229_player_016/io_out[3] shadow1229_player_016/io_out[4] shadow1229_player_016/io_out[5]
+ shadow1229_player_016/io_out[6] shadow1229_player_016/io_out[7] vccd1 vssd1 shadow1229_player
Xscanchain_119 scanchain_119/clk_in scanchain_120/clk_in scanchain_119/data_in scanchain_120/data_in
+ scanchain_119/latch_enable_in scanchain_120/latch_enable_in scanchain_119/module_data_in[0]
+ scanchain_119/module_data_in[1] scanchain_119/module_data_in[2] scanchain_119/module_data_in[3]
+ scanchain_119/module_data_in[4] scanchain_119/module_data_in[5] scanchain_119/module_data_in[6]
+ scanchain_119/module_data_in[7] scanchain_119/module_data_out[0] scanchain_119/module_data_out[1]
+ scanchain_119/module_data_out[2] scanchain_119/module_data_out[3] scanchain_119/module_data_out[4]
+ scanchain_119/module_data_out[5] scanchain_119/module_data_out[6] scanchain_119/module_data_out[7]
+ scanchain_119/scan_select_in scanchain_120/scan_select_in vccd1 vssd1 scanchain
Xscanchain_108 scanchain_108/clk_in scanchain_109/clk_in scanchain_108/data_in scanchain_109/data_in
+ scanchain_108/latch_enable_in scanchain_109/latch_enable_in scanchain_108/module_data_in[0]
+ scanchain_108/module_data_in[1] scanchain_108/module_data_in[2] scanchain_108/module_data_in[3]
+ scanchain_108/module_data_in[4] scanchain_108/module_data_in[5] scanchain_108/module_data_in[6]
+ scanchain_108/module_data_in[7] scanchain_108/module_data_out[0] scanchain_108/module_data_out[1]
+ scanchain_108/module_data_out[2] scanchain_108/module_data_out[3] scanchain_108/module_data_out[4]
+ scanchain_108/module_data_out[5] scanchain_108/module_data_out[6] scanchain_108/module_data_out[7]
+ scanchain_108/scan_select_in scanchain_109/scan_select_in vccd1 vssd1 scanchain
Xuser_module_361728533238569985_224 scanchain_224/module_data_in[0] scanchain_224/module_data_in[1]
+ scanchain_224/module_data_in[2] scanchain_224/module_data_in[3] scanchain_224/module_data_in[4]
+ scanchain_224/module_data_in[5] scanchain_224/module_data_in[6] scanchain_224/module_data_in[7]
+ scanchain_224/module_data_out[0] scanchain_224/module_data_out[1] scanchain_224/module_data_out[2]
+ scanchain_224/module_data_out[3] scanchain_224/module_data_out[4] scanchain_224/module_data_out[5]
+ scanchain_224/module_data_out[6] scanchain_224/module_data_out[7] vccd1 vssd1 user_module_361728533238569985
Xuser_module_361728533238569985_235 scanchain_235/module_data_in[0] scanchain_235/module_data_in[1]
+ scanchain_235/module_data_in[2] scanchain_235/module_data_in[3] scanchain_235/module_data_in[4]
+ scanchain_235/module_data_in[5] scanchain_235/module_data_in[6] scanchain_235/module_data_in[7]
+ scanchain_235/module_data_out[0] scanchain_235/module_data_out[1] scanchain_235/module_data_out[2]
+ scanchain_235/module_data_out[3] scanchain_235/module_data_out[4] scanchain_235/module_data_out[5]
+ scanchain_235/module_data_out[6] scanchain_235/module_data_out[7] vccd1 vssd1 user_module_361728533238569985
Xuser_module_361728533238569985_246 scanchain_246/module_data_in[0] scanchain_246/module_data_in[1]
+ scanchain_246/module_data_in[2] scanchain_246/module_data_in[3] scanchain_246/module_data_in[4]
+ scanchain_246/module_data_in[5] scanchain_246/module_data_in[6] scanchain_246/module_data_in[7]
+ scanchain_246/module_data_out[0] scanchain_246/module_data_out[1] scanchain_246/module_data_out[2]
+ scanchain_246/module_data_out[3] scanchain_246/module_data_out[4] scanchain_246/module_data_out[5]
+ scanchain_246/module_data_out[6] scanchain_246/module_data_out[7] vccd1 vssd1 user_module_361728533238569985
Xuser_module_361728533238569985_213 scanchain_213/module_data_in[0] scanchain_213/module_data_in[1]
+ scanchain_213/module_data_in[2] scanchain_213/module_data_in[3] scanchain_213/module_data_in[4]
+ scanchain_213/module_data_in[5] scanchain_213/module_data_in[6] scanchain_213/module_data_in[7]
+ scanchain_213/module_data_out[0] scanchain_213/module_data_out[1] scanchain_213/module_data_out[2]
+ scanchain_213/module_data_out[3] scanchain_213/module_data_out[4] scanchain_213/module_data_out[5]
+ scanchain_213/module_data_out[6] scanchain_213/module_data_out[7] vccd1 vssd1 user_module_361728533238569985
Xgbsha_ttfir_top_044 gbsha_ttfir_top_044/io_in[0] gbsha_ttfir_top_044/io_in[1] gbsha_ttfir_top_044/io_in[2]
+ gbsha_ttfir_top_044/io_in[3] gbsha_ttfir_top_044/io_in[4] gbsha_ttfir_top_044/io_in[5]
+ gbsha_ttfir_top_044/io_in[6] gbsha_ttfir_top_044/io_in[7] gbsha_ttfir_top_044/io_out[0]
+ gbsha_ttfir_top_044/io_out[1] gbsha_ttfir_top_044/io_out[2] gbsha_ttfir_top_044/io_out[3]
+ gbsha_ttfir_top_044/io_out[4] gbsha_ttfir_top_044/io_out[5] gbsha_ttfir_top_044/io_out[6]
+ gbsha_ttfir_top_044/io_out[7] vccd1 vssd1 gbsha_ttfir_top
Xuser_module_361728533238569985_202 scanchain_202/module_data_in[0] scanchain_202/module_data_in[1]
+ scanchain_202/module_data_in[2] scanchain_202/module_data_in[3] scanchain_202/module_data_in[4]
+ scanchain_202/module_data_in[5] scanchain_202/module_data_in[6] scanchain_202/module_data_in[7]
+ scanchain_202/module_data_out[0] scanchain_202/module_data_out[1] scanchain_202/module_data_out[2]
+ scanchain_202/module_data_out[3] scanchain_202/module_data_out[4] scanchain_202/module_data_out[5]
+ scanchain_202/module_data_out[6] scanchain_202/module_data_out[7] vccd1 vssd1 user_module_361728533238569985
Xuser_module_361728533238569985_098 scanchain_098/module_data_in[0] scanchain_098/module_data_in[1]
+ scanchain_098/module_data_in[2] scanchain_098/module_data_in[3] scanchain_098/module_data_in[4]
+ scanchain_098/module_data_in[5] scanchain_098/module_data_in[6] scanchain_098/module_data_in[7]
+ scanchain_098/module_data_out[0] scanchain_098/module_data_out[1] scanchain_098/module_data_out[2]
+ scanchain_098/module_data_out[3] scanchain_098/module_data_out[4] scanchain_098/module_data_out[5]
+ scanchain_098/module_data_out[6] scanchain_098/module_data_out[7] vccd1 vssd1 user_module_361728533238569985
Xdiferential_rvb2_023 diferential_rvb2_023/io_in[0] diferential_rvb2_023/io_in[1]
+ diferential_rvb2_023/io_in[2] diferential_rvb2_023/io_in[3] diferential_rvb2_023/io_in[4]
+ diferential_rvb2_023/io_in[5] diferential_rvb2_023/io_in[6] diferential_rvb2_023/io_in[7]
+ diferential_rvb2_023/io_out[0] diferential_rvb2_023/io_out[1] diferential_rvb2_023/io_out[2]
+ diferential_rvb2_023/io_out[3] diferential_rvb2_023/io_out[4] diferential_rvb2_023/io_out[5]
+ diferential_rvb2_023/io_out[6] diferential_rvb2_023/io_out[7] vccd1 vssd1 diferential_rvb2
Xgreenstyle_lfsr_013 greenstyle_lfsr_013/io_in[0] greenstyle_lfsr_013/io_in[1] greenstyle_lfsr_013/io_in[2]
+ greenstyle_lfsr_013/io_in[3] greenstyle_lfsr_013/io_in[4] greenstyle_lfsr_013/io_in[5]
+ greenstyle_lfsr_013/io_in[6] greenstyle_lfsr_013/io_in[7] greenstyle_lfsr_013/io_out[0]
+ greenstyle_lfsr_013/io_out[1] greenstyle_lfsr_013/io_out[2] greenstyle_lfsr_013/io_out[3]
+ greenstyle_lfsr_013/io_out[4] greenstyle_lfsr_013/io_out[5] greenstyle_lfsr_013/io_out[6]
+ greenstyle_lfsr_013/io_out[7] vccd1 vssd1 greenstyle_lfsr
XHiddenRoom_HiddenCPU_065 scanchain_065/module_data_in[0] scanchain_065/module_data_in[1]
+ scanchain_065/module_data_in[2] scanchain_065/module_data_in[3] scanchain_065/module_data_in[4]
+ scanchain_065/module_data_in[5] scanchain_065/module_data_in[6] scanchain_065/module_data_in[7]
+ scanchain_065/module_data_out[0] scanchain_065/module_data_out[1] scanchain_065/module_data_out[2]
+ scanchain_065/module_data_out[3] scanchain_065/module_data_out[4] scanchain_065/module_data_out[5]
+ scanchain_065/module_data_out[6] scanchain_065/module_data_out[7] vccd1 vssd1 HiddenRoom_HiddenCPU
Xscanchain_109 scanchain_109/clk_in scanchain_110/clk_in scanchain_109/data_in scanchain_110/data_in
+ scanchain_109/latch_enable_in scanchain_110/latch_enable_in scanchain_109/module_data_in[0]
+ scanchain_109/module_data_in[1] scanchain_109/module_data_in[2] scanchain_109/module_data_in[3]
+ scanchain_109/module_data_in[4] scanchain_109/module_data_in[5] scanchain_109/module_data_in[6]
+ scanchain_109/module_data_in[7] scanchain_109/module_data_out[0] scanchain_109/module_data_out[1]
+ scanchain_109/module_data_out[2] scanchain_109/module_data_out[3] scanchain_109/module_data_out[4]
+ scanchain_109/module_data_out[5] scanchain_109/module_data_out[6] scanchain_109/module_data_out[7]
+ scanchain_109/scan_select_in scanchain_110/scan_select_in vccd1 vssd1 scanchain
Xuser_module_361728533238569985_225 scanchain_225/module_data_in[0] scanchain_225/module_data_in[1]
+ scanchain_225/module_data_in[2] scanchain_225/module_data_in[3] scanchain_225/module_data_in[4]
+ scanchain_225/module_data_in[5] scanchain_225/module_data_in[6] scanchain_225/module_data_in[7]
+ scanchain_225/module_data_out[0] scanchain_225/module_data_out[1] scanchain_225/module_data_out[2]
+ scanchain_225/module_data_out[3] scanchain_225/module_data_out[4] scanchain_225/module_data_out[5]
+ scanchain_225/module_data_out[6] scanchain_225/module_data_out[7] vccd1 vssd1 user_module_361728533238569985
Xuser_module_361728533238569985_236 scanchain_236/module_data_in[0] scanchain_236/module_data_in[1]
+ scanchain_236/module_data_in[2] scanchain_236/module_data_in[3] scanchain_236/module_data_in[4]
+ scanchain_236/module_data_in[5] scanchain_236/module_data_in[6] scanchain_236/module_data_in[7]
+ scanchain_236/module_data_out[0] scanchain_236/module_data_out[1] scanchain_236/module_data_out[2]
+ scanchain_236/module_data_out[3] scanchain_236/module_data_out[4] scanchain_236/module_data_out[5]
+ scanchain_236/module_data_out[6] scanchain_236/module_data_out[7] vccd1 vssd1 user_module_361728533238569985
Xuser_module_361728533238569985_247 scanchain_247/module_data_in[0] scanchain_247/module_data_in[1]
+ scanchain_247/module_data_in[2] scanchain_247/module_data_in[3] scanchain_247/module_data_in[4]
+ scanchain_247/module_data_in[5] scanchain_247/module_data_in[6] scanchain_247/module_data_in[7]
+ scanchain_247/module_data_out[0] scanchain_247/module_data_out[1] scanchain_247/module_data_out[2]
+ scanchain_247/module_data_out[3] scanchain_247/module_data_out[4] scanchain_247/module_data_out[5]
+ scanchain_247/module_data_out[6] scanchain_247/module_data_out[7] vccd1 vssd1 user_module_361728533238569985
Xuser_module_361728533238569985_214 scanchain_214/module_data_in[0] scanchain_214/module_data_in[1]
+ scanchain_214/module_data_in[2] scanchain_214/module_data_in[3] scanchain_214/module_data_in[4]
+ scanchain_214/module_data_in[5] scanchain_214/module_data_in[6] scanchain_214/module_data_in[7]
+ scanchain_214/module_data_out[0] scanchain_214/module_data_out[1] scanchain_214/module_data_out[2]
+ scanchain_214/module_data_out[3] scanchain_214/module_data_out[4] scanchain_214/module_data_out[5]
+ scanchain_214/module_data_out[6] scanchain_214/module_data_out[7] vccd1 vssd1 user_module_361728533238569985
Xuser_module_361728533238569985_203 scanchain_203/module_data_in[0] scanchain_203/module_data_in[1]
+ scanchain_203/module_data_in[2] scanchain_203/module_data_in[3] scanchain_203/module_data_in[4]
+ scanchain_203/module_data_in[5] scanchain_203/module_data_in[6] scanchain_203/module_data_in[7]
+ scanchain_203/module_data_out[0] scanchain_203/module_data_out[1] scanchain_203/module_data_out[2]
+ scanchain_203/module_data_out[3] scanchain_203/module_data_out[4] scanchain_203/module_data_out[5]
+ scanchain_203/module_data_out[6] scanchain_203/module_data_out[7] vccd1 vssd1 user_module_361728533238569985
Xuser_module_361728533238569985_099 scanchain_099/module_data_in[0] scanchain_099/module_data_in[1]
+ scanchain_099/module_data_in[2] scanchain_099/module_data_in[3] scanchain_099/module_data_in[4]
+ scanchain_099/module_data_in[5] scanchain_099/module_data_in[6] scanchain_099/module_data_in[7]
+ scanchain_099/module_data_out[0] scanchain_099/module_data_out[1] scanchain_099/module_data_out[2]
+ scanchain_099/module_data_out[3] scanchain_099/module_data_out[4] scanchain_099/module_data_out[5]
+ scanchain_099/module_data_out[6] scanchain_099/module_data_out[7] vccd1 vssd1 user_module_361728533238569985
Xuser_module_361728533238569985_000 scanchain_000/module_data_in[0] scanchain_000/module_data_in[1]
+ scanchain_000/module_data_in[2] scanchain_000/module_data_in[3] scanchain_000/module_data_in[4]
+ scanchain_000/module_data_in[5] scanchain_000/module_data_in[6] scanchain_000/module_data_in[7]
+ scanchain_000/module_data_out[0] scanchain_000/module_data_out[1] scanchain_000/module_data_out[2]
+ scanchain_000/module_data_out[3] scanchain_000/module_data_out[4] scanchain_000/module_data_out[5]
+ scanchain_000/module_data_out[6] scanchain_000/module_data_out[7] vccd1 vssd1 user_module_361728533238569985
Xdratini0_pov_display_top_041 scanchain_041/module_data_in[0] scanchain_041/module_data_in[1]
+ scanchain_041/module_data_in[2] scanchain_041/module_data_in[3] scanchain_041/module_data_in[4]
+ scanchain_041/module_data_in[5] scanchain_041/module_data_in[6] scanchain_041/module_data_in[7]
+ scanchain_041/module_data_out[0] scanchain_041/module_data_out[1] scanchain_041/module_data_out[2]
+ scanchain_041/module_data_out[3] scanchain_041/module_data_out[4] scanchain_041/module_data_out[5]
+ scanchain_041/module_data_out[6] scanchain_041/module_data_out[7] vccd1 vssd1 dratini0_pov_display_top
Xwormy_top_004 wormy_top_004/io_in[0] wormy_top_004/io_in[1] wormy_top_004/io_in[2]
+ wormy_top_004/io_in[3] wormy_top_004/io_in[4] wormy_top_004/io_in[5] wormy_top_004/io_in[6]
+ wormy_top_004/io_in[7] wormy_top_004/io_out[0] wormy_top_004/io_out[1] wormy_top_004/io_out[2]
+ wormy_top_004/io_out[3] wormy_top_004/io_out[4] wormy_top_004/io_out[5] wormy_top_004/io_out[6]
+ wormy_top_004/io_out[7] vccd1 vssd1 wormy_top
Xbat52_pwm_ddpm_top_033 scanchain_033/module_data_in[0] scanchain_033/module_data_in[1]
+ scanchain_033/module_data_in[2] scanchain_033/module_data_in[3] scanchain_033/module_data_in[4]
+ scanchain_033/module_data_in[5] scanchain_033/module_data_in[6] scanchain_033/module_data_in[7]
+ scanchain_033/module_data_out[0] scanchain_033/module_data_out[1] scanchain_033/module_data_out[2]
+ scanchain_033/module_data_out[3] scanchain_033/module_data_out[4] scanchain_033/module_data_out[5]
+ scanchain_033/module_data_out[6] scanchain_033/module_data_out[7] vccd1 vssd1 bat52_pwm_ddpm_top
Xuser_module_361728533238569985_226 scanchain_226/module_data_in[0] scanchain_226/module_data_in[1]
+ scanchain_226/module_data_in[2] scanchain_226/module_data_in[3] scanchain_226/module_data_in[4]
+ scanchain_226/module_data_in[5] scanchain_226/module_data_in[6] scanchain_226/module_data_in[7]
+ scanchain_226/module_data_out[0] scanchain_226/module_data_out[1] scanchain_226/module_data_out[2]
+ scanchain_226/module_data_out[3] scanchain_226/module_data_out[4] scanchain_226/module_data_out[5]
+ scanchain_226/module_data_out[6] scanchain_226/module_data_out[7] vccd1 vssd1 user_module_361728533238569985
Xuser_module_361728533238569985_237 scanchain_237/module_data_in[0] scanchain_237/module_data_in[1]
+ scanchain_237/module_data_in[2] scanchain_237/module_data_in[3] scanchain_237/module_data_in[4]
+ scanchain_237/module_data_in[5] scanchain_237/module_data_in[6] scanchain_237/module_data_in[7]
+ scanchain_237/module_data_out[0] scanchain_237/module_data_out[1] scanchain_237/module_data_out[2]
+ scanchain_237/module_data_out[3] scanchain_237/module_data_out[4] scanchain_237/module_data_out[5]
+ scanchain_237/module_data_out[6] scanchain_237/module_data_out[7] vccd1 vssd1 user_module_361728533238569985
Xuser_module_361728533238569985_248 scanchain_248/module_data_in[0] scanchain_248/module_data_in[1]
+ scanchain_248/module_data_in[2] scanchain_248/module_data_in[3] scanchain_248/module_data_in[4]
+ scanchain_248/module_data_in[5] scanchain_248/module_data_in[6] scanchain_248/module_data_in[7]
+ scanchain_248/module_data_out[0] scanchain_248/module_data_out[1] scanchain_248/module_data_out[2]
+ scanchain_248/module_data_out[3] scanchain_248/module_data_out[4] scanchain_248/module_data_out[5]
+ scanchain_248/module_data_out[6] scanchain_248/module_data_out[7] vccd1 vssd1 user_module_361728533238569985
Xuser_module_361728533238569985_215 scanchain_215/module_data_in[0] scanchain_215/module_data_in[1]
+ scanchain_215/module_data_in[2] scanchain_215/module_data_in[3] scanchain_215/module_data_in[4]
+ scanchain_215/module_data_in[5] scanchain_215/module_data_in[6] scanchain_215/module_data_in[7]
+ scanchain_215/module_data_out[0] scanchain_215/module_data_out[1] scanchain_215/module_data_out[2]
+ scanchain_215/module_data_out[3] scanchain_215/module_data_out[4] scanchain_215/module_data_out[5]
+ scanchain_215/module_data_out[6] scanchain_215/module_data_out[7] vccd1 vssd1 user_module_361728533238569985
Xuser_module_361728533238569985_204 scanchain_204/module_data_in[0] scanchain_204/module_data_in[1]
+ scanchain_204/module_data_in[2] scanchain_204/module_data_in[3] scanchain_204/module_data_in[4]
+ scanchain_204/module_data_in[5] scanchain_204/module_data_in[6] scanchain_204/module_data_in[7]
+ scanchain_204/module_data_out[0] scanchain_204/module_data_out[1] scanchain_204/module_data_out[2]
+ scanchain_204/module_data_out[3] scanchain_204/module_data_out[4] scanchain_204/module_data_out[5]
+ scanchain_204/module_data_out[6] scanchain_204/module_data_out[7] vccd1 vssd1 user_module_361728533238569985
Xuser_module_361728533238569985_089 scanchain_089/module_data_in[0] scanchain_089/module_data_in[1]
+ scanchain_089/module_data_in[2] scanchain_089/module_data_in[3] scanchain_089/module_data_in[4]
+ scanchain_089/module_data_in[5] scanchain_089/module_data_in[6] scanchain_089/module_data_in[7]
+ scanchain_089/module_data_out[0] scanchain_089/module_data_out[1] scanchain_089/module_data_out[2]
+ scanchain_089/module_data_out[3] scanchain_089/module_data_out[4] scanchain_089/module_data_out[5]
+ scanchain_089/module_data_out[6] scanchain_089/module_data_out[7] vccd1 vssd1 user_module_361728533238569985
Xscanchain_090 scanchain_090/clk_in scanchain_091/clk_in scanchain_090/data_in scanchain_091/data_in
+ scanchain_090/latch_enable_in scanchain_091/latch_enable_in scanchain_090/module_data_in[0]
+ scanchain_090/module_data_in[1] scanchain_090/module_data_in[2] scanchain_090/module_data_in[3]
+ scanchain_090/module_data_in[4] scanchain_090/module_data_in[5] scanchain_090/module_data_in[6]
+ scanchain_090/module_data_in[7] scanchain_090/module_data_out[0] scanchain_090/module_data_out[1]
+ scanchain_090/module_data_out[2] scanchain_090/module_data_out[3] scanchain_090/module_data_out[4]
+ scanchain_090/module_data_out[5] scanchain_090/module_data_out[6] scanchain_090/module_data_out[7]
+ scanchain_090/scan_select_in scanchain_091/scan_select_in vccd1 vssd1 scanchain
Xuser_module_361728533238569985_238 scanchain_238/module_data_in[0] scanchain_238/module_data_in[1]
+ scanchain_238/module_data_in[2] scanchain_238/module_data_in[3] scanchain_238/module_data_in[4]
+ scanchain_238/module_data_in[5] scanchain_238/module_data_in[6] scanchain_238/module_data_in[7]
+ scanchain_238/module_data_out[0] scanchain_238/module_data_out[1] scanchain_238/module_data_out[2]
+ scanchain_238/module_data_out[3] scanchain_238/module_data_out[4] scanchain_238/module_data_out[5]
+ scanchain_238/module_data_out[6] scanchain_238/module_data_out[7] vccd1 vssd1 user_module_361728533238569985
Xuser_module_361728533238569985_249 scanchain_249/module_data_in[0] scanchain_249/module_data_in[1]
+ scanchain_249/module_data_in[2] scanchain_249/module_data_in[3] scanchain_249/module_data_in[4]
+ scanchain_249/module_data_in[5] scanchain_249/module_data_in[6] scanchain_249/module_data_in[7]
+ scanchain_249/module_data_out[0] scanchain_249/module_data_out[1] scanchain_249/module_data_out[2]
+ scanchain_249/module_data_out[3] scanchain_249/module_data_out[4] scanchain_249/module_data_out[5]
+ scanchain_249/module_data_out[6] scanchain_249/module_data_out[7] vccd1 vssd1 user_module_361728533238569985
Xuser_module_361728533238569985_227 scanchain_227/module_data_in[0] scanchain_227/module_data_in[1]
+ scanchain_227/module_data_in[2] scanchain_227/module_data_in[3] scanchain_227/module_data_in[4]
+ scanchain_227/module_data_in[5] scanchain_227/module_data_in[6] scanchain_227/module_data_in[7]
+ scanchain_227/module_data_out[0] scanchain_227/module_data_out[1] scanchain_227/module_data_out[2]
+ scanchain_227/module_data_out[3] scanchain_227/module_data_out[4] scanchain_227/module_data_out[5]
+ scanchain_227/module_data_out[6] scanchain_227/module_data_out[7] vccd1 vssd1 user_module_361728533238569985
Xuser_module_361728533238569985_216 scanchain_216/module_data_in[0] scanchain_216/module_data_in[1]
+ scanchain_216/module_data_in[2] scanchain_216/module_data_in[3] scanchain_216/module_data_in[4]
+ scanchain_216/module_data_in[5] scanchain_216/module_data_in[6] scanchain_216/module_data_in[7]
+ scanchain_216/module_data_out[0] scanchain_216/module_data_out[1] scanchain_216/module_data_out[2]
+ scanchain_216/module_data_out[3] scanchain_216/module_data_out[4] scanchain_216/module_data_out[5]
+ scanchain_216/module_data_out[6] scanchain_216/module_data_out[7] vccd1 vssd1 user_module_361728533238569985
Xuser_module_361728533238569985_205 scanchain_205/module_data_in[0] scanchain_205/module_data_in[1]
+ scanchain_205/module_data_in[2] scanchain_205/module_data_in[3] scanchain_205/module_data_in[4]
+ scanchain_205/module_data_in[5] scanchain_205/module_data_in[6] scanchain_205/module_data_in[7]
+ scanchain_205/module_data_out[0] scanchain_205/module_data_out[1] scanchain_205/module_data_out[2]
+ scanchain_205/module_data_out[3] scanchain_205/module_data_out[4] scanchain_205/module_data_out[5]
+ scanchain_205/module_data_out[6] scanchain_205/module_data_out[7] vccd1 vssd1 user_module_361728533238569985
Xuser_module_340805072482992722_056 scanchain_056/module_data_in[0] scanchain_056/module_data_in[1]
+ scanchain_056/module_data_in[2] scanchain_056/module_data_in[3] scanchain_056/module_data_in[4]
+ scanchain_056/module_data_in[5] scanchain_056/module_data_in[6] scanchain_056/module_data_in[7]
+ scanchain_056/module_data_out[0] scanchain_056/module_data_out[1] scanchain_056/module_data_out[2]
+ scanchain_056/module_data_out[3] scanchain_056/module_data_out[4] scanchain_056/module_data_out[5]
+ scanchain_056/module_data_out[6] scanchain_056/module_data_out[7] vccd1 vssd1 user_module_340805072482992722
Xclemensnasenberg_top_069 scanchain_069/module_data_in[0] scanchain_069/module_data_in[1]
+ scanchain_069/module_data_in[2] scanchain_069/module_data_in[3] scanchain_069/module_data_in[4]
+ scanchain_069/module_data_in[5] scanchain_069/module_data_in[6] scanchain_069/module_data_in[7]
+ scanchain_069/module_data_out[0] scanchain_069/module_data_out[1] scanchain_069/module_data_out[2]
+ scanchain_069/module_data_out[3] scanchain_069/module_data_out[4] scanchain_069/module_data_out[5]
+ scanchain_069/module_data_out[6] scanchain_069/module_data_out[7] vccd1 vssd1 clemensnasenberg_top
Xblueintegral_mat_mult_078 scanchain_078/module_data_in[0] scanchain_078/module_data_in[1]
+ scanchain_078/module_data_in[2] scanchain_078/module_data_in[3] scanchain_078/module_data_in[4]
+ scanchain_078/module_data_in[5] scanchain_078/module_data_in[6] scanchain_078/module_data_in[7]
+ scanchain_078/module_data_out[0] scanchain_078/module_data_out[1] scanchain_078/module_data_out[2]
+ scanchain_078/module_data_out[3] scanchain_078/module_data_out[4] scanchain_078/module_data_out[5]
+ scanchain_078/module_data_out[6] scanchain_078/module_data_out[7] vccd1 vssd1 blueintegral_mat_mult
Xscanchain_091 scanchain_091/clk_in scanchain_092/clk_in scanchain_091/data_in scanchain_092/data_in
+ scanchain_091/latch_enable_in scanchain_092/latch_enable_in scanchain_091/module_data_in[0]
+ scanchain_091/module_data_in[1] scanchain_091/module_data_in[2] scanchain_091/module_data_in[3]
+ scanchain_091/module_data_in[4] scanchain_091/module_data_in[5] scanchain_091/module_data_in[6]
+ scanchain_091/module_data_in[7] scanchain_091/module_data_out[0] scanchain_091/module_data_out[1]
+ scanchain_091/module_data_out[2] scanchain_091/module_data_out[3] scanchain_091/module_data_out[4]
+ scanchain_091/module_data_out[5] scanchain_091/module_data_out[6] scanchain_091/module_data_out[7]
+ scanchain_091/scan_select_in scanchain_092/scan_select_in vccd1 vssd1 scanchain
Xwokwi_tt03_simon_top_037 scanchain_037/module_data_in[0] scanchain_037/module_data_in[1]
+ scanchain_037/module_data_in[2] scanchain_037/module_data_in[3] scanchain_037/module_data_in[4]
+ scanchain_037/module_data_in[5] scanchain_037/module_data_in[6] scanchain_037/module_data_in[7]
+ scanchain_037/module_data_out[0] scanchain_037/module_data_out[1] scanchain_037/module_data_out[2]
+ scanchain_037/module_data_out[3] scanchain_037/module_data_out[4] scanchain_037/module_data_out[5]
+ scanchain_037/module_data_out[6] scanchain_037/module_data_out[7] vccd1 vssd1 wokwi_tt03_simon_top
Xscanchain_080 scanchain_080/clk_in scanchain_081/clk_in scanchain_080/data_in scanchain_081/data_in
+ scanchain_080/latch_enable_in scanchain_081/latch_enable_in scanchain_080/module_data_in[0]
+ scanchain_080/module_data_in[1] scanchain_080/module_data_in[2] scanchain_080/module_data_in[3]
+ scanchain_080/module_data_in[4] scanchain_080/module_data_in[5] scanchain_080/module_data_in[6]
+ scanchain_080/module_data_in[7] scanchain_080/module_data_out[0] scanchain_080/module_data_out[1]
+ scanchain_080/module_data_out[2] scanchain_080/module_data_out[3] scanchain_080/module_data_out[4]
+ scanchain_080/module_data_out[5] scanchain_080/module_data_out[6] scanchain_080/module_data_out[7]
+ scanchain_080/scan_select_in scanchain_081/scan_select_in vccd1 vssd1 scanchain
Xuser_module_361728533238569985_239 scanchain_239/module_data_in[0] scanchain_239/module_data_in[1]
+ scanchain_239/module_data_in[2] scanchain_239/module_data_in[3] scanchain_239/module_data_in[4]
+ scanchain_239/module_data_in[5] scanchain_239/module_data_in[6] scanchain_239/module_data_in[7]
+ scanchain_239/module_data_out[0] scanchain_239/module_data_out[1] scanchain_239/module_data_out[2]
+ scanchain_239/module_data_out[3] scanchain_239/module_data_out[4] scanchain_239/module_data_out[5]
+ scanchain_239/module_data_out[6] scanchain_239/module_data_out[7] vccd1 vssd1 user_module_361728533238569985
Xuser_module_361728533238569985_228 scanchain_228/module_data_in[0] scanchain_228/module_data_in[1]
+ scanchain_228/module_data_in[2] scanchain_228/module_data_in[3] scanchain_228/module_data_in[4]
+ scanchain_228/module_data_in[5] scanchain_228/module_data_in[6] scanchain_228/module_data_in[7]
+ scanchain_228/module_data_out[0] scanchain_228/module_data_out[1] scanchain_228/module_data_out[2]
+ scanchain_228/module_data_out[3] scanchain_228/module_data_out[4] scanchain_228/module_data_out[5]
+ scanchain_228/module_data_out[6] scanchain_228/module_data_out[7] vccd1 vssd1 user_module_361728533238569985
Xuser_module_361728533238569985_217 scanchain_217/module_data_in[0] scanchain_217/module_data_in[1]
+ scanchain_217/module_data_in[2] scanchain_217/module_data_in[3] scanchain_217/module_data_in[4]
+ scanchain_217/module_data_in[5] scanchain_217/module_data_in[6] scanchain_217/module_data_in[7]
+ scanchain_217/module_data_out[0] scanchain_217/module_data_out[1] scanchain_217/module_data_out[2]
+ scanchain_217/module_data_out[3] scanchain_217/module_data_out[4] scanchain_217/module_data_out[5]
+ scanchain_217/module_data_out[6] scanchain_217/module_data_out[7] vccd1 vssd1 user_module_361728533238569985
Xuser_module_361728533238569985_206 scanchain_206/module_data_in[0] scanchain_206/module_data_in[1]
+ scanchain_206/module_data_in[2] scanchain_206/module_data_in[3] scanchain_206/module_data_in[4]
+ scanchain_206/module_data_in[5] scanchain_206/module_data_in[6] scanchain_206/module_data_in[7]
+ scanchain_206/module_data_out[0] scanchain_206/module_data_out[1] scanchain_206/module_data_out[2]
+ scanchain_206/module_data_out[3] scanchain_206/module_data_out[4] scanchain_206/module_data_out[5]
+ scanchain_206/module_data_out[6] scanchain_206/module_data_out[7] vccd1 vssd1 user_module_361728533238569985
Xscanchain_240 scanchain_240/clk_in scanchain_241/clk_in scanchain_240/data_in scanchain_241/data_in
+ scanchain_240/latch_enable_in scanchain_241/latch_enable_in scanchain_240/module_data_in[0]
+ scanchain_240/module_data_in[1] scanchain_240/module_data_in[2] scanchain_240/module_data_in[3]
+ scanchain_240/module_data_in[4] scanchain_240/module_data_in[5] scanchain_240/module_data_in[6]
+ scanchain_240/module_data_in[7] scanchain_240/module_data_out[0] scanchain_240/module_data_out[1]
+ scanchain_240/module_data_out[2] scanchain_240/module_data_out[3] scanchain_240/module_data_out[4]
+ scanchain_240/module_data_out[5] scanchain_240/module_data_out[6] scanchain_240/module_data_out[7]
+ scanchain_240/scan_select_in scanchain_241/scan_select_in vccd1 vssd1 scanchain
Xscanchain_070 scanchain_070/clk_in scanchain_071/clk_in scanchain_070/data_in scanchain_071/data_in
+ scanchain_070/latch_enable_in scanchain_071/latch_enable_in s4ga_070/io_in[0] s4ga_070/io_in[1]
+ s4ga_070/io_in[2] s4ga_070/io_in[3] s4ga_070/io_in[4] s4ga_070/io_in[5] s4ga_070/io_in[6]
+ s4ga_070/io_in[7] s4ga_070/io_out[0] s4ga_070/io_out[1] s4ga_070/io_out[2] s4ga_070/io_out[3]
+ s4ga_070/io_out[4] s4ga_070/io_out[5] s4ga_070/io_out[6] s4ga_070/io_out[7] scanchain_070/scan_select_in
+ scanchain_071/scan_select_in vccd1 vssd1 scanchain
Xscanchain_081 scanchain_081/clk_in scanchain_082/clk_in scanchain_081/data_in scanchain_082/data_in
+ scanchain_081/latch_enable_in scanchain_082/latch_enable_in scanchain_081/module_data_in[0]
+ scanchain_081/module_data_in[1] scanchain_081/module_data_in[2] scanchain_081/module_data_in[3]
+ scanchain_081/module_data_in[4] scanchain_081/module_data_in[5] scanchain_081/module_data_in[6]
+ scanchain_081/module_data_in[7] scanchain_081/module_data_out[0] scanchain_081/module_data_out[1]
+ scanchain_081/module_data_out[2] scanchain_081/module_data_out[3] scanchain_081/module_data_out[4]
+ scanchain_081/module_data_out[5] scanchain_081/module_data_out[6] scanchain_081/module_data_out[7]
+ scanchain_081/scan_select_in scanchain_082/scan_select_in vccd1 vssd1 scanchain
Xuser_module_362867354023533569_083 scanchain_083/module_data_in[0] scanchain_083/module_data_in[1]
+ scanchain_083/module_data_in[2] scanchain_083/module_data_in[3] scanchain_083/module_data_in[4]
+ scanchain_083/module_data_in[5] scanchain_083/module_data_in[6] scanchain_083/module_data_in[7]
+ scanchain_083/module_data_out[0] scanchain_083/module_data_out[1] scanchain_083/module_data_out[2]
+ scanchain_083/module_data_out[3] scanchain_083/module_data_out[4] scanchain_083/module_data_out[5]
+ scanchain_083/module_data_out[6] scanchain_083/module_data_out[7] vccd1 vssd1 user_module_362867354023533569
Xscanchain_092 scanchain_092/clk_in scanchain_093/clk_in scanchain_092/data_in scanchain_093/data_in
+ scanchain_092/latch_enable_in scanchain_093/latch_enable_in scanchain_092/module_data_in[0]
+ scanchain_092/module_data_in[1] scanchain_092/module_data_in[2] scanchain_092/module_data_in[3]
+ scanchain_092/module_data_in[4] scanchain_092/module_data_in[5] scanchain_092/module_data_in[6]
+ scanchain_092/module_data_in[7] scanchain_092/module_data_out[0] scanchain_092/module_data_out[1]
+ scanchain_092/module_data_out[2] scanchain_092/module_data_out[3] scanchain_092/module_data_out[4]
+ scanchain_092/module_data_out[5] scanchain_092/module_data_out[6] scanchain_092/module_data_out[7]
+ scanchain_092/scan_select_in scanchain_093/scan_select_in vccd1 vssd1 scanchain
Xuser_module_362249236392794113_079 scanchain_079/module_data_in[0] scanchain_079/module_data_in[1]
+ scanchain_079/module_data_in[2] scanchain_079/module_data_in[3] scanchain_079/module_data_in[4]
+ scanchain_079/module_data_in[5] scanchain_079/module_data_in[6] scanchain_079/module_data_in[7]
+ scanchain_079/module_data_out[0] scanchain_079/module_data_out[1] scanchain_079/module_data_out[2]
+ scanchain_079/module_data_out[3] scanchain_079/module_data_out[4] scanchain_079/module_data_out[5]
+ scanchain_079/module_data_out[6] scanchain_079/module_data_out[7] vccd1 vssd1 user_module_362249236392794113
Xuser_module_362441918332875777_084 scanchain_084/module_data_in[0] scanchain_084/module_data_in[1]
+ scanchain_084/module_data_in[2] scanchain_084/module_data_in[3] scanchain_084/module_data_in[4]
+ scanchain_084/module_data_in[5] scanchain_084/module_data_in[6] scanchain_084/module_data_in[7]
+ scanchain_084/module_data_out[0] scanchain_084/module_data_out[1] scanchain_084/module_data_out[2]
+ scanchain_084/module_data_out[3] scanchain_084/module_data_out[4] scanchain_084/module_data_out[5]
+ scanchain_084/module_data_out[6] scanchain_084/module_data_out[7] vccd1 vssd1 user_module_362441918332875777
Xuser_module_361728533238569985_229 scanchain_229/module_data_in[0] scanchain_229/module_data_in[1]
+ scanchain_229/module_data_in[2] scanchain_229/module_data_in[3] scanchain_229/module_data_in[4]
+ scanchain_229/module_data_in[5] scanchain_229/module_data_in[6] scanchain_229/module_data_in[7]
+ scanchain_229/module_data_out[0] scanchain_229/module_data_out[1] scanchain_229/module_data_out[2]
+ scanchain_229/module_data_out[3] scanchain_229/module_data_out[4] scanchain_229/module_data_out[5]
+ scanchain_229/module_data_out[6] scanchain_229/module_data_out[7] vccd1 vssd1 user_module_361728533238569985
Xuser_module_361728533238569985_218 scanchain_218/module_data_in[0] scanchain_218/module_data_in[1]
+ scanchain_218/module_data_in[2] scanchain_218/module_data_in[3] scanchain_218/module_data_in[4]
+ scanchain_218/module_data_in[5] scanchain_218/module_data_in[6] scanchain_218/module_data_in[7]
+ scanchain_218/module_data_out[0] scanchain_218/module_data_out[1] scanchain_218/module_data_out[2]
+ scanchain_218/module_data_out[3] scanchain_218/module_data_out[4] scanchain_218/module_data_out[5]
+ scanchain_218/module_data_out[6] scanchain_218/module_data_out[7] vccd1 vssd1 user_module_361728533238569985
Xuser_module_361728533238569985_207 scanchain_207/module_data_in[0] scanchain_207/module_data_in[1]
+ scanchain_207/module_data_in[2] scanchain_207/module_data_in[3] scanchain_207/module_data_in[4]
+ scanchain_207/module_data_in[5] scanchain_207/module_data_in[6] scanchain_207/module_data_in[7]
+ scanchain_207/module_data_out[0] scanchain_207/module_data_out[1] scanchain_207/module_data_out[2]
+ scanchain_207/module_data_out[3] scanchain_207/module_data_out[4] scanchain_207/module_data_out[5]
+ scanchain_207/module_data_out[6] scanchain_207/module_data_out[7] vccd1 vssd1 user_module_361728533238569985
Xhtfab_microtapeout_046 scanchain_046/module_data_in[0] scanchain_046/module_data_in[1]
+ scanchain_046/module_data_in[2] scanchain_046/module_data_in[3] scanchain_046/module_data_in[4]
+ scanchain_046/module_data_in[5] scanchain_046/module_data_in[6] scanchain_046/module_data_in[7]
+ scanchain_046/module_data_out[0] scanchain_046/module_data_out[1] scanchain_046/module_data_out[2]
+ scanchain_046/module_data_out[3] scanchain_046/module_data_out[4] scanchain_046/module_data_out[5]
+ scanchain_046/module_data_out[6] scanchain_046/module_data_out[7] vccd1 vssd1 htfab_microtapeout
Xhpretl_tt03_temperature_sensor_048 scanchain_048/module_data_in[0] scanchain_048/module_data_in[1]
+ scanchain_048/module_data_in[2] scanchain_048/module_data_in[3] scanchain_048/module_data_in[4]
+ scanchain_048/module_data_in[5] scanchain_048/module_data_in[6] scanchain_048/module_data_in[7]
+ scanchain_048/module_data_out[0] scanchain_048/module_data_out[1] scanchain_048/module_data_out[2]
+ scanchain_048/module_data_out[3] scanchain_048/module_data_out[4] scanchain_048/module_data_out[5]
+ scanchain_048/module_data_out[6] scanchain_048/module_data_out[7] vccd1 vssd1 hpretl_tt03_temperature_sensor
Xscanchain_230 scanchain_230/clk_in scanchain_231/clk_in scanchain_230/data_in scanchain_231/data_in
+ scanchain_230/latch_enable_in scanchain_231/latch_enable_in scanchain_230/module_data_in[0]
+ scanchain_230/module_data_in[1] scanchain_230/module_data_in[2] scanchain_230/module_data_in[3]
+ scanchain_230/module_data_in[4] scanchain_230/module_data_in[5] scanchain_230/module_data_in[6]
+ scanchain_230/module_data_in[7] scanchain_230/module_data_out[0] scanchain_230/module_data_out[1]
+ scanchain_230/module_data_out[2] scanchain_230/module_data_out[3] scanchain_230/module_data_out[4]
+ scanchain_230/module_data_out[5] scanchain_230/module_data_out[6] scanchain_230/module_data_out[7]
+ scanchain_230/scan_select_in scanchain_231/scan_select_in vccd1 vssd1 scanchain
Xscanchain_241 scanchain_241/clk_in scanchain_242/clk_in scanchain_241/data_in scanchain_242/data_in
+ scanchain_241/latch_enable_in scanchain_242/latch_enable_in scanchain_241/module_data_in[0]
+ scanchain_241/module_data_in[1] scanchain_241/module_data_in[2] scanchain_241/module_data_in[3]
+ scanchain_241/module_data_in[4] scanchain_241/module_data_in[5] scanchain_241/module_data_in[6]
+ scanchain_241/module_data_in[7] scanchain_241/module_data_out[0] scanchain_241/module_data_out[1]
+ scanchain_241/module_data_out[2] scanchain_241/module_data_out[3] scanchain_241/module_data_out[4]
+ scanchain_241/module_data_out[5] scanchain_241/module_data_out[6] scanchain_241/module_data_out[7]
+ scanchain_241/scan_select_in scanchain_242/scan_select_in vccd1 vssd1 scanchain
Xzl_uart_066 zl_uart_066/io_in[0] zl_uart_066/io_in[1] zl_uart_066/io_in[2] zl_uart_066/io_in[3]
+ zl_uart_066/io_in[4] zl_uart_066/io_in[5] zl_uart_066/io_in[6] zl_uart_066/io_in[7]
+ zl_uart_066/io_out[0] zl_uart_066/io_out[1] zl_uart_066/io_out[2] zl_uart_066/io_out[3]
+ zl_uart_066/io_out[4] zl_uart_066/io_out[5] zl_uart_066/io_out[6] zl_uart_066/io_out[7]
+ vccd1 vssd1 zl_uart
Xtinysat_039 tinysat_039/io_in[0] tinysat_039/io_in[1] tinysat_039/io_in[2] tinysat_039/io_in[3]
+ tinysat_039/io_in[4] tinysat_039/io_in[5] tinysat_039/io_in[6] tinysat_039/io_in[7]
+ tinysat_039/io_out[0] tinysat_039/io_out[1] tinysat_039/io_out[2] tinysat_039/io_out[3]
+ tinysat_039/io_out[4] tinysat_039/io_out[5] tinysat_039/io_out[6] tinysat_039/io_out[7]
+ vccd1 vssd1 tinysat
Xscanchain_060 scanchain_060/clk_in scanchain_061/clk_in scanchain_060/data_in scanchain_061/data_in
+ scanchain_060/latch_enable_in scanchain_061/latch_enable_in FSM_LAT_060/io_in[0]
+ FSM_LAT_060/io_in[1] FSM_LAT_060/io_in[2] FSM_LAT_060/io_in[3] FSM_LAT_060/io_in[4]
+ FSM_LAT_060/io_in[5] FSM_LAT_060/io_in[6] FSM_LAT_060/io_in[7] FSM_LAT_060/io_out[0]
+ FSM_LAT_060/io_out[1] FSM_LAT_060/io_out[2] FSM_LAT_060/io_out[3] FSM_LAT_060/io_out[4]
+ FSM_LAT_060/io_out[5] FSM_LAT_060/io_out[6] FSM_LAT_060/io_out[7] scanchain_060/scan_select_in
+ scanchain_061/scan_select_in vccd1 vssd1 scanchain
Xscanchain_071 scanchain_071/clk_in scanchain_072/clk_in scanchain_071/data_in scanchain_072/data_in
+ scanchain_071/latch_enable_in scanchain_072/latch_enable_in scanchain_071/module_data_in[0]
+ scanchain_071/module_data_in[1] scanchain_071/module_data_in[2] scanchain_071/module_data_in[3]
+ scanchain_071/module_data_in[4] scanchain_071/module_data_in[5] scanchain_071/module_data_in[6]
+ scanchain_071/module_data_in[7] scanchain_071/module_data_out[0] scanchain_071/module_data_out[1]
+ scanchain_071/module_data_out[2] scanchain_071/module_data_out[3] scanchain_071/module_data_out[4]
+ scanchain_071/module_data_out[5] scanchain_071/module_data_out[6] scanchain_071/module_data_out[7]
+ scanchain_071/scan_select_in scanchain_072/scan_select_in vccd1 vssd1 scanchain
Xscanchain_082 scanchain_082/clk_in scanchain_083/clk_in scanchain_082/data_in scanchain_083/data_in
+ scanchain_082/latch_enable_in scanchain_083/latch_enable_in scanchain_082/module_data_in[0]
+ scanchain_082/module_data_in[1] scanchain_082/module_data_in[2] scanchain_082/module_data_in[3]
+ scanchain_082/module_data_in[4] scanchain_082/module_data_in[5] scanchain_082/module_data_in[6]
+ scanchain_082/module_data_in[7] scanchain_082/module_data_out[0] scanchain_082/module_data_out[1]
+ scanchain_082/module_data_out[2] scanchain_082/module_data_out[3] scanchain_082/module_data_out[4]
+ scanchain_082/module_data_out[5] scanchain_082/module_data_out[6] scanchain_082/module_data_out[7]
+ scanchain_082/scan_select_in scanchain_083/scan_select_in vccd1 vssd1 scanchain
Xscanchain_093 scanchain_093/clk_in scanchain_094/clk_in scanchain_093/data_in scanchain_094/data_in
+ scanchain_093/latch_enable_in scanchain_094/latch_enable_in scanchain_093/module_data_in[0]
+ scanchain_093/module_data_in[1] scanchain_093/module_data_in[2] scanchain_093/module_data_in[3]
+ scanchain_093/module_data_in[4] scanchain_093/module_data_in[5] scanchain_093/module_data_in[6]
+ scanchain_093/module_data_in[7] scanchain_093/module_data_out[0] scanchain_093/module_data_out[1]
+ scanchain_093/module_data_out[2] scanchain_093/module_data_out[3] scanchain_093/module_data_out[4]
+ scanchain_093/module_data_out[5] scanchain_093/module_data_out[6] scanchain_093/module_data_out[7]
+ scanchain_093/scan_select_in scanchain_094/scan_select_in vccd1 vssd1 scanchain
Xuser_module_361728533238569985_219 scanchain_219/module_data_in[0] scanchain_219/module_data_in[1]
+ scanchain_219/module_data_in[2] scanchain_219/module_data_in[3] scanchain_219/module_data_in[4]
+ scanchain_219/module_data_in[5] scanchain_219/module_data_in[6] scanchain_219/module_data_in[7]
+ scanchain_219/module_data_out[0] scanchain_219/module_data_out[1] scanchain_219/module_data_out[2]
+ scanchain_219/module_data_out[3] scanchain_219/module_data_out[4] scanchain_219/module_data_out[5]
+ scanchain_219/module_data_out[6] scanchain_219/module_data_out[7] vccd1 vssd1 user_module_361728533238569985
Xuser_module_361728533238569985_208 scanchain_208/module_data_in[0] scanchain_208/module_data_in[1]
+ scanchain_208/module_data_in[2] scanchain_208/module_data_in[3] scanchain_208/module_data_in[4]
+ scanchain_208/module_data_in[5] scanchain_208/module_data_in[6] scanchain_208/module_data_in[7]
+ scanchain_208/module_data_out[0] scanchain_208/module_data_out[1] scanchain_208/module_data_out[2]
+ scanchain_208/module_data_out[3] scanchain_208/module_data_out[4] scanchain_208/module_data_out[5]
+ scanchain_208/module_data_out[6] scanchain_208/module_data_out[7] vccd1 vssd1 user_module_361728533238569985
Xdwisehart_ring_top_081 scanchain_081/module_data_in[0] scanchain_081/module_data_in[1]
+ scanchain_081/module_data_in[2] scanchain_081/module_data_in[3] scanchain_081/module_data_in[4]
+ scanchain_081/module_data_in[5] scanchain_081/module_data_in[6] scanchain_081/module_data_in[7]
+ scanchain_081/module_data_out[0] scanchain_081/module_data_out[1] scanchain_081/module_data_out[2]
+ scanchain_081/module_data_out[3] scanchain_081/module_data_out[4] scanchain_081/module_data_out[5]
+ scanchain_081/module_data_out[6] scanchain_081/module_data_out[7] vccd1 vssd1 dwisehart_ring_top
Xjmw95_top_067 jmw95_top_067/io_in[0] jmw95_top_067/io_in[1] jmw95_top_067/io_in[2]
+ jmw95_top_067/io_in[3] jmw95_top_067/io_in[4] jmw95_top_067/io_in[5] jmw95_top_067/io_in[6]
+ jmw95_top_067/io_in[7] jmw95_top_067/io_out[0] jmw95_top_067/io_out[1] jmw95_top_067/io_out[2]
+ jmw95_top_067/io_out[3] jmw95_top_067/io_out[4] jmw95_top_067/io_out[5] jmw95_top_067/io_out[6]
+ jmw95_top_067/io_out[7] vccd1 vssd1 jmw95_top
Xscanchain_231 scanchain_231/clk_in scanchain_232/clk_in scanchain_231/data_in scanchain_232/data_in
+ scanchain_231/latch_enable_in scanchain_232/latch_enable_in scanchain_231/module_data_in[0]
+ scanchain_231/module_data_in[1] scanchain_231/module_data_in[2] scanchain_231/module_data_in[3]
+ scanchain_231/module_data_in[4] scanchain_231/module_data_in[5] scanchain_231/module_data_in[6]
+ scanchain_231/module_data_in[7] scanchain_231/module_data_out[0] scanchain_231/module_data_out[1]
+ scanchain_231/module_data_out[2] scanchain_231/module_data_out[3] scanchain_231/module_data_out[4]
+ scanchain_231/module_data_out[5] scanchain_231/module_data_out[6] scanchain_231/module_data_out[7]
+ scanchain_231/scan_select_in scanchain_232/scan_select_in vccd1 vssd1 scanchain
Xscanchain_242 scanchain_242/clk_in scanchain_243/clk_in scanchain_242/data_in scanchain_243/data_in
+ scanchain_242/latch_enable_in scanchain_243/latch_enable_in scanchain_242/module_data_in[0]
+ scanchain_242/module_data_in[1] scanchain_242/module_data_in[2] scanchain_242/module_data_in[3]
+ scanchain_242/module_data_in[4] scanchain_242/module_data_in[5] scanchain_242/module_data_in[6]
+ scanchain_242/module_data_in[7] scanchain_242/module_data_out[0] scanchain_242/module_data_out[1]
+ scanchain_242/module_data_out[2] scanchain_242/module_data_out[3] scanchain_242/module_data_out[4]
+ scanchain_242/module_data_out[5] scanchain_242/module_data_out[6] scanchain_242/module_data_out[7]
+ scanchain_242/scan_select_in scanchain_243/scan_select_in vccd1 vssd1 scanchain
Xscanchain_220 scanchain_220/clk_in scanchain_221/clk_in scanchain_220/data_in scanchain_221/data_in
+ scanchain_220/latch_enable_in scanchain_221/latch_enable_in scanchain_220/module_data_in[0]
+ scanchain_220/module_data_in[1] scanchain_220/module_data_in[2] scanchain_220/module_data_in[3]
+ scanchain_220/module_data_in[4] scanchain_220/module_data_in[5] scanchain_220/module_data_in[6]
+ scanchain_220/module_data_in[7] scanchain_220/module_data_out[0] scanchain_220/module_data_out[1]
+ scanchain_220/module_data_out[2] scanchain_220/module_data_out[3] scanchain_220/module_data_out[4]
+ scanchain_220/module_data_out[5] scanchain_220/module_data_out[6] scanchain_220/module_data_out[7]
+ scanchain_220/scan_select_in scanchain_221/scan_select_in vccd1 vssd1 scanchain
Xscanchain_050 scanchain_050/clk_in scanchain_051/clk_in scanchain_050/data_in scanchain_051/data_in
+ scanchain_050/latch_enable_in scanchain_051/latch_enable_in pwm_050/io_in[0] pwm_050/io_in[1]
+ pwm_050/io_in[2] pwm_050/io_in[3] pwm_050/io_in[4] pwm_050/io_in[5] pwm_050/io_in[6]
+ pwm_050/io_in[7] pwm_050/io_out[0] pwm_050/io_out[1] pwm_050/io_out[2] pwm_050/io_out[3]
+ pwm_050/io_out[4] pwm_050/io_out[5] pwm_050/io_out[6] pwm_050/io_out[7] scanchain_050/scan_select_in
+ scanchain_051/scan_select_in vccd1 vssd1 scanchain
Xscanchain_061 scanchain_061/clk_in scanchain_062/clk_in scanchain_061/data_in scanchain_062/data_in
+ scanchain_061/latch_enable_in scanchain_062/latch_enable_in scanchain_061/module_data_in[0]
+ scanchain_061/module_data_in[1] scanchain_061/module_data_in[2] scanchain_061/module_data_in[3]
+ scanchain_061/module_data_in[4] scanchain_061/module_data_in[5] scanchain_061/module_data_in[6]
+ scanchain_061/module_data_in[7] scanchain_061/module_data_out[0] scanchain_061/module_data_out[1]
+ scanchain_061/module_data_out[2] scanchain_061/module_data_out[3] scanchain_061/module_data_out[4]
+ scanchain_061/module_data_out[5] scanchain_061/module_data_out[6] scanchain_061/module_data_out[7]
+ scanchain_061/scan_select_in scanchain_062/scan_select_in vccd1 vssd1 scanchain
Xscanchain_072 scanchain_072/clk_in scanchain_073/clk_in scanchain_072/data_in scanchain_073/data_in
+ scanchain_072/latch_enable_in scanchain_073/latch_enable_in tiny_bnn_072/io_in[0]
+ tiny_bnn_072/io_in[1] tiny_bnn_072/io_in[2] tiny_bnn_072/io_in[3] tiny_bnn_072/io_in[4]
+ tiny_bnn_072/io_in[5] tiny_bnn_072/io_in[6] tiny_bnn_072/io_in[7] tiny_bnn_072/io_out[0]
+ tiny_bnn_072/io_out[1] tiny_bnn_072/io_out[2] tiny_bnn_072/io_out[3] tiny_bnn_072/io_out[4]
+ tiny_bnn_072/io_out[5] tiny_bnn_072/io_out[6] tiny_bnn_072/io_out[7] scanchain_072/scan_select_in
+ scanchain_073/scan_select_in vccd1 vssd1 scanchain
Xscanchain_083 scanchain_083/clk_in scanchain_084/clk_in scanchain_083/data_in scanchain_084/data_in
+ scanchain_083/latch_enable_in scanchain_084/latch_enable_in scanchain_083/module_data_in[0]
+ scanchain_083/module_data_in[1] scanchain_083/module_data_in[2] scanchain_083/module_data_in[3]
+ scanchain_083/module_data_in[4] scanchain_083/module_data_in[5] scanchain_083/module_data_in[6]
+ scanchain_083/module_data_in[7] scanchain_083/module_data_out[0] scanchain_083/module_data_out[1]
+ scanchain_083/module_data_out[2] scanchain_083/module_data_out[3] scanchain_083/module_data_out[4]
+ scanchain_083/module_data_out[5] scanchain_083/module_data_out[6] scanchain_083/module_data_out[7]
+ scanchain_083/scan_select_in scanchain_084/scan_select_in vccd1 vssd1 scanchain
Xscanchain_094 scanchain_094/clk_in scanchain_095/clk_in scanchain_094/data_in scanchain_095/data_in
+ scanchain_094/latch_enable_in scanchain_095/latch_enable_in scanchain_094/module_data_in[0]
+ scanchain_094/module_data_in[1] scanchain_094/module_data_in[2] scanchain_094/module_data_in[3]
+ scanchain_094/module_data_in[4] scanchain_094/module_data_in[5] scanchain_094/module_data_in[6]
+ scanchain_094/module_data_in[7] scanchain_094/module_data_out[0] scanchain_094/module_data_out[1]
+ scanchain_094/module_data_out[2] scanchain_094/module_data_out[3] scanchain_094/module_data_out[4]
+ scanchain_094/module_data_out[5] scanchain_094/module_data_out[6] scanchain_094/module_data_out[7]
+ scanchain_094/scan_select_in scanchain_095/scan_select_in vccd1 vssd1 scanchain
Xuser_module_361728533238569985_209 scanchain_209/module_data_in[0] scanchain_209/module_data_in[1]
+ scanchain_209/module_data_in[2] scanchain_209/module_data_in[3] scanchain_209/module_data_in[4]
+ scanchain_209/module_data_in[5] scanchain_209/module_data_in[6] scanchain_209/module_data_in[7]
+ scanchain_209/module_data_out[0] scanchain_209/module_data_out[1] scanchain_209/module_data_out[2]
+ scanchain_209/module_data_out[3] scanchain_209/module_data_out[4] scanchain_209/module_data_out[5]
+ scanchain_209/module_data_out[6] scanchain_209/module_data_out[7] vccd1 vssd1 user_module_361728533238569985
Xuser_module_361684719151591425_036 scanchain_036/module_data_in[0] scanchain_036/module_data_in[1]
+ scanchain_036/module_data_in[2] scanchain_036/module_data_in[3] scanchain_036/module_data_in[4]
+ scanchain_036/module_data_in[5] scanchain_036/module_data_in[6] scanchain_036/module_data_in[7]
+ scanchain_036/module_data_out[0] scanchain_036/module_data_out[1] scanchain_036/module_data_out[2]
+ scanchain_036/module_data_out[3] scanchain_036/module_data_out[4] scanchain_036/module_data_out[5]
+ scanchain_036/module_data_out[6] scanchain_036/module_data_out[7] vccd1 vssd1 user_module_361684719151591425
Xdsp_4bits_seq_alu_049 dsp_4bits_seq_alu_049/io_in[0] dsp_4bits_seq_alu_049/io_in[1]
+ dsp_4bits_seq_alu_049/io_in[2] dsp_4bits_seq_alu_049/io_in[3] dsp_4bits_seq_alu_049/io_in[4]
+ dsp_4bits_seq_alu_049/io_in[5] dsp_4bits_seq_alu_049/io_in[6] dsp_4bits_seq_alu_049/io_in[7]
+ dsp_4bits_seq_alu_049/io_out[0] dsp_4bits_seq_alu_049/io_out[1] dsp_4bits_seq_alu_049/io_out[2]
+ dsp_4bits_seq_alu_049/io_out[3] dsp_4bits_seq_alu_049/io_out[4] dsp_4bits_seq_alu_049/io_out[5]
+ dsp_4bits_seq_alu_049/io_out[6] dsp_4bits_seq_alu_049/io_out[7] vccd1 vssd1 dsp_4bits_seq_alu
Xscanchain_232 scanchain_232/clk_in scanchain_233/clk_in scanchain_232/data_in scanchain_233/data_in
+ scanchain_232/latch_enable_in scanchain_233/latch_enable_in scanchain_232/module_data_in[0]
+ scanchain_232/module_data_in[1] scanchain_232/module_data_in[2] scanchain_232/module_data_in[3]
+ scanchain_232/module_data_in[4] scanchain_232/module_data_in[5] scanchain_232/module_data_in[6]
+ scanchain_232/module_data_in[7] scanchain_232/module_data_out[0] scanchain_232/module_data_out[1]
+ scanchain_232/module_data_out[2] scanchain_232/module_data_out[3] scanchain_232/module_data_out[4]
+ scanchain_232/module_data_out[5] scanchain_232/module_data_out[6] scanchain_232/module_data_out[7]
+ scanchain_232/scan_select_in scanchain_233/scan_select_in vccd1 vssd1 scanchain
Xscanchain_243 scanchain_243/clk_in scanchain_244/clk_in scanchain_243/data_in scanchain_244/data_in
+ scanchain_243/latch_enable_in scanchain_244/latch_enable_in scanchain_243/module_data_in[0]
+ scanchain_243/module_data_in[1] scanchain_243/module_data_in[2] scanchain_243/module_data_in[3]
+ scanchain_243/module_data_in[4] scanchain_243/module_data_in[5] scanchain_243/module_data_in[6]
+ scanchain_243/module_data_in[7] scanchain_243/module_data_out[0] scanchain_243/module_data_out[1]
+ scanchain_243/module_data_out[2] scanchain_243/module_data_out[3] scanchain_243/module_data_out[4]
+ scanchain_243/module_data_out[5] scanchain_243/module_data_out[6] scanchain_243/module_data_out[7]
+ scanchain_243/scan_select_in scanchain_244/scan_select_in vccd1 vssd1 scanchain
Xscanchain_221 scanchain_221/clk_in scanchain_222/clk_in scanchain_221/data_in scanchain_222/data_in
+ scanchain_221/latch_enable_in scanchain_222/latch_enable_in scanchain_221/module_data_in[0]
+ scanchain_221/module_data_in[1] scanchain_221/module_data_in[2] scanchain_221/module_data_in[3]
+ scanchain_221/module_data_in[4] scanchain_221/module_data_in[5] scanchain_221/module_data_in[6]
+ scanchain_221/module_data_in[7] scanchain_221/module_data_out[0] scanchain_221/module_data_out[1]
+ scanchain_221/module_data_out[2] scanchain_221/module_data_out[3] scanchain_221/module_data_out[4]
+ scanchain_221/module_data_out[5] scanchain_221/module_data_out[6] scanchain_221/module_data_out[7]
+ scanchain_221/scan_select_in scanchain_222/scan_select_in vccd1 vssd1 scanchain
Xscanchain_210 scanchain_210/clk_in scanchain_211/clk_in scanchain_210/data_in scanchain_211/data_in
+ scanchain_210/latch_enable_in scanchain_211/latch_enable_in scanchain_210/module_data_in[0]
+ scanchain_210/module_data_in[1] scanchain_210/module_data_in[2] scanchain_210/module_data_in[3]
+ scanchain_210/module_data_in[4] scanchain_210/module_data_in[5] scanchain_210/module_data_in[6]
+ scanchain_210/module_data_in[7] scanchain_210/module_data_out[0] scanchain_210/module_data_out[1]
+ scanchain_210/module_data_out[2] scanchain_210/module_data_out[3] scanchain_210/module_data_out[4]
+ scanchain_210/module_data_out[5] scanchain_210/module_data_out[6] scanchain_210/module_data_out[7]
+ scanchain_210/scan_select_in scanchain_211/scan_select_in vccd1 vssd1 scanchain
Xscanchain_040 scanchain_040/clk_in scanchain_041/clk_in scanchain_040/data_in scanchain_041/data_in
+ scanchain_040/latch_enable_in scanchain_041/latch_enable_in scanchain_040/module_data_in[0]
+ scanchain_040/module_data_in[1] scanchain_040/module_data_in[2] scanchain_040/module_data_in[3]
+ scanchain_040/module_data_in[4] scanchain_040/module_data_in[5] scanchain_040/module_data_in[6]
+ scanchain_040/module_data_in[7] scanchain_040/module_data_out[0] scanchain_040/module_data_out[1]
+ scanchain_040/module_data_out[2] scanchain_040/module_data_out[3] scanchain_040/module_data_out[4]
+ scanchain_040/module_data_out[5] scanchain_040/module_data_out[6] scanchain_040/module_data_out[7]
+ scanchain_040/scan_select_in scanchain_041/scan_select_in vccd1 vssd1 scanchain
Xscanchain_051 scanchain_051/clk_in scanchain_052/clk_in scanchain_051/data_in scanchain_052/data_in
+ scanchain_051/latch_enable_in scanchain_052/latch_enable_in scanchain_051/module_data_in[0]
+ scanchain_051/module_data_in[1] scanchain_051/module_data_in[2] scanchain_051/module_data_in[3]
+ scanchain_051/module_data_in[4] scanchain_051/module_data_in[5] scanchain_051/module_data_in[6]
+ scanchain_051/module_data_in[7] scanchain_051/module_data_out[0] scanchain_051/module_data_out[1]
+ scanchain_051/module_data_out[2] scanchain_051/module_data_out[3] scanchain_051/module_data_out[4]
+ scanchain_051/module_data_out[5] scanchain_051/module_data_out[6] scanchain_051/module_data_out[7]
+ scanchain_051/scan_select_in scanchain_052/scan_select_in vccd1 vssd1 scanchain
Xscanchain_073 scanchain_073/clk_in scanchain_074/clk_in scanchain_073/data_in scanchain_074/data_in
+ scanchain_073/latch_enable_in scanchain_074/latch_enable_in lucaz97_tt_top_073/io_in[0]
+ lucaz97_tt_top_073/io_in[1] lucaz97_tt_top_073/io_in[2] lucaz97_tt_top_073/io_in[3]
+ lucaz97_tt_top_073/io_in[4] lucaz97_tt_top_073/io_in[5] lucaz97_tt_top_073/io_in[6]
+ lucaz97_tt_top_073/io_in[7] lucaz97_tt_top_073/io_out[0] lucaz97_tt_top_073/io_out[1]
+ lucaz97_tt_top_073/io_out[2] lucaz97_tt_top_073/io_out[3] lucaz97_tt_top_073/io_out[4]
+ lucaz97_tt_top_073/io_out[5] lucaz97_tt_top_073/io_out[6] lucaz97_tt_top_073/io_out[7]
+ scanchain_073/scan_select_in scanchain_074/scan_select_in vccd1 vssd1 scanchain
Xscanchain_062 scanchain_062/clk_in scanchain_063/clk_in scanchain_062/data_in scanchain_063/data_in
+ scanchain_062/latch_enable_in scanchain_063/latch_enable_in scanchain_062/module_data_in[0]
+ scanchain_062/module_data_in[1] scanchain_062/module_data_in[2] scanchain_062/module_data_in[3]
+ scanchain_062/module_data_in[4] scanchain_062/module_data_in[5] scanchain_062/module_data_in[6]
+ scanchain_062/module_data_in[7] scanchain_062/module_data_out[0] scanchain_062/module_data_out[1]
+ scanchain_062/module_data_out[2] scanchain_062/module_data_out[3] scanchain_062/module_data_out[4]
+ scanchain_062/module_data_out[5] scanchain_062/module_data_out[6] scanchain_062/module_data_out[7]
+ scanchain_062/scan_select_in scanchain_063/scan_select_in vccd1 vssd1 scanchain
Xscanchain_084 scanchain_084/clk_in scanchain_085/clk_in scanchain_084/data_in scanchain_085/data_in
+ scanchain_084/latch_enable_in scanchain_085/latch_enable_in scanchain_084/module_data_in[0]
+ scanchain_084/module_data_in[1] scanchain_084/module_data_in[2] scanchain_084/module_data_in[3]
+ scanchain_084/module_data_in[4] scanchain_084/module_data_in[5] scanchain_084/module_data_in[6]
+ scanchain_084/module_data_in[7] scanchain_084/module_data_out[0] scanchain_084/module_data_out[1]
+ scanchain_084/module_data_out[2] scanchain_084/module_data_out[3] scanchain_084/module_data_out[4]
+ scanchain_084/module_data_out[5] scanchain_084/module_data_out[6] scanchain_084/module_data_out[7]
+ scanchain_084/scan_select_in scanchain_085/scan_select_in vccd1 vssd1 scanchain
Xscanchain_095 scanchain_095/clk_in scanchain_096/clk_in scanchain_095/data_in scanchain_096/data_in
+ scanchain_095/latch_enable_in scanchain_096/latch_enable_in scanchain_095/module_data_in[0]
+ scanchain_095/module_data_in[1] scanchain_095/module_data_in[2] scanchain_095/module_data_in[3]
+ scanchain_095/module_data_in[4] scanchain_095/module_data_in[5] scanchain_095/module_data_in[6]
+ scanchain_095/module_data_in[7] scanchain_095/module_data_out[0] scanchain_095/module_data_out[1]
+ scanchain_095/module_data_out[2] scanchain_095/module_data_out[3] scanchain_095/module_data_out[4]
+ scanchain_095/module_data_out[5] scanchain_095/module_data_out[6] scanchain_095/module_data_out[7]
+ scanchain_095/scan_select_in scanchain_096/scan_select_in vccd1 vssd1 scanchain
Xguianmonezm_ezmcpu_030 scanchain_030/module_data_in[0] scanchain_030/module_data_in[1]
+ scanchain_030/module_data_in[2] scanchain_030/module_data_in[3] scanchain_030/module_data_in[4]
+ scanchain_030/module_data_in[5] scanchain_030/module_data_in[6] scanchain_030/module_data_in[7]
+ scanchain_030/module_data_out[0] scanchain_030/module_data_out[1] scanchain_030/module_data_out[2]
+ scanchain_030/module_data_out[3] scanchain_030/module_data_out[4] scanchain_030/module_data_out[5]
+ scanchain_030/module_data_out[6] scanchain_030/module_data_out[7] vccd1 vssd1 guianmonezm_ezmcpu
Xlukevassallo_xor_cipher_027 scanchain_027/module_data_in[0] scanchain_027/module_data_in[1]
+ scanchain_027/module_data_in[2] scanchain_027/module_data_in[3] scanchain_027/module_data_in[4]
+ scanchain_027/module_data_in[5] scanchain_027/module_data_in[6] scanchain_027/module_data_in[7]
+ scanchain_027/module_data_out[0] scanchain_027/module_data_out[1] scanchain_027/module_data_out[2]
+ scanchain_027/module_data_out[3] scanchain_027/module_data_out[4] scanchain_027/module_data_out[5]
+ scanchain_027/module_data_out[6] scanchain_027/module_data_out[7] vccd1 vssd1 lukevassallo_xor_cipher
Xscanchain_233 scanchain_233/clk_in scanchain_234/clk_in scanchain_233/data_in scanchain_234/data_in
+ scanchain_233/latch_enable_in scanchain_234/latch_enable_in scanchain_233/module_data_in[0]
+ scanchain_233/module_data_in[1] scanchain_233/module_data_in[2] scanchain_233/module_data_in[3]
+ scanchain_233/module_data_in[4] scanchain_233/module_data_in[5] scanchain_233/module_data_in[6]
+ scanchain_233/module_data_in[7] scanchain_233/module_data_out[0] scanchain_233/module_data_out[1]
+ scanchain_233/module_data_out[2] scanchain_233/module_data_out[3] scanchain_233/module_data_out[4]
+ scanchain_233/module_data_out[5] scanchain_233/module_data_out[6] scanchain_233/module_data_out[7]
+ scanchain_233/scan_select_in scanchain_234/scan_select_in vccd1 vssd1 scanchain
Xscanchain_244 scanchain_244/clk_in scanchain_245/clk_in scanchain_244/data_in scanchain_245/data_in
+ scanchain_244/latch_enable_in scanchain_245/latch_enable_in scanchain_244/module_data_in[0]
+ scanchain_244/module_data_in[1] scanchain_244/module_data_in[2] scanchain_244/module_data_in[3]
+ scanchain_244/module_data_in[4] scanchain_244/module_data_in[5] scanchain_244/module_data_in[6]
+ scanchain_244/module_data_in[7] scanchain_244/module_data_out[0] scanchain_244/module_data_out[1]
+ scanchain_244/module_data_out[2] scanchain_244/module_data_out[3] scanchain_244/module_data_out[4]
+ scanchain_244/module_data_out[5] scanchain_244/module_data_out[6] scanchain_244/module_data_out[7]
+ scanchain_244/scan_select_in scanchain_245/scan_select_in vccd1 vssd1 scanchain
Xscanchain_222 scanchain_222/clk_in scanchain_223/clk_in scanchain_222/data_in scanchain_223/data_in
+ scanchain_222/latch_enable_in scanchain_223/latch_enable_in scanchain_222/module_data_in[0]
+ scanchain_222/module_data_in[1] scanchain_222/module_data_in[2] scanchain_222/module_data_in[3]
+ scanchain_222/module_data_in[4] scanchain_222/module_data_in[5] scanchain_222/module_data_in[6]
+ scanchain_222/module_data_in[7] scanchain_222/module_data_out[0] scanchain_222/module_data_out[1]
+ scanchain_222/module_data_out[2] scanchain_222/module_data_out[3] scanchain_222/module_data_out[4]
+ scanchain_222/module_data_out[5] scanchain_222/module_data_out[6] scanchain_222/module_data_out[7]
+ scanchain_222/scan_select_in scanchain_223/scan_select_in vccd1 vssd1 scanchain
Xscanchain_211 scanchain_211/clk_in scanchain_212/clk_in scanchain_211/data_in scanchain_212/data_in
+ scanchain_211/latch_enable_in scanchain_212/latch_enable_in scanchain_211/module_data_in[0]
+ scanchain_211/module_data_in[1] scanchain_211/module_data_in[2] scanchain_211/module_data_in[3]
+ scanchain_211/module_data_in[4] scanchain_211/module_data_in[5] scanchain_211/module_data_in[6]
+ scanchain_211/module_data_in[7] scanchain_211/module_data_out[0] scanchain_211/module_data_out[1]
+ scanchain_211/module_data_out[2] scanchain_211/module_data_out[3] scanchain_211/module_data_out[4]
+ scanchain_211/module_data_out[5] scanchain_211/module_data_out[6] scanchain_211/module_data_out[7]
+ scanchain_211/scan_select_in scanchain_212/scan_select_in vccd1 vssd1 scanchain
Xscanchain_200 scanchain_200/clk_in scanchain_201/clk_in scanchain_200/data_in scanchain_201/data_in
+ scanchain_200/latch_enable_in scanchain_201/latch_enable_in scanchain_200/module_data_in[0]
+ scanchain_200/module_data_in[1] scanchain_200/module_data_in[2] scanchain_200/module_data_in[3]
+ scanchain_200/module_data_in[4] scanchain_200/module_data_in[5] scanchain_200/module_data_in[6]
+ scanchain_200/module_data_in[7] scanchain_200/module_data_out[0] scanchain_200/module_data_out[1]
+ scanchain_200/module_data_out[2] scanchain_200/module_data_out[3] scanchain_200/module_data_out[4]
+ scanchain_200/module_data_out[5] scanchain_200/module_data_out[6] scanchain_200/module_data_out[7]
+ scanchain_200/scan_select_in scanchain_201/scan_select_in vccd1 vssd1 scanchain
Xscanchain_030 scanchain_030/clk_in scanchain_031/clk_in scanchain_030/data_in scanchain_031/data_in
+ scanchain_030/latch_enable_in scanchain_031/latch_enable_in scanchain_030/module_data_in[0]
+ scanchain_030/module_data_in[1] scanchain_030/module_data_in[2] scanchain_030/module_data_in[3]
+ scanchain_030/module_data_in[4] scanchain_030/module_data_in[5] scanchain_030/module_data_in[6]
+ scanchain_030/module_data_in[7] scanchain_030/module_data_out[0] scanchain_030/module_data_out[1]
+ scanchain_030/module_data_out[2] scanchain_030/module_data_out[3] scanchain_030/module_data_out[4]
+ scanchain_030/module_data_out[5] scanchain_030/module_data_out[6] scanchain_030/module_data_out[7]
+ scanchain_030/scan_select_in scanchain_031/scan_select_in vccd1 vssd1 scanchain
Xscanchain_041 scanchain_041/clk_in scanchain_042/clk_in scanchain_041/data_in scanchain_042/data_in
+ scanchain_041/latch_enable_in scanchain_042/latch_enable_in scanchain_041/module_data_in[0]
+ scanchain_041/module_data_in[1] scanchain_041/module_data_in[2] scanchain_041/module_data_in[3]
+ scanchain_041/module_data_in[4] scanchain_041/module_data_in[5] scanchain_041/module_data_in[6]
+ scanchain_041/module_data_in[7] scanchain_041/module_data_out[0] scanchain_041/module_data_out[1]
+ scanchain_041/module_data_out[2] scanchain_041/module_data_out[3] scanchain_041/module_data_out[4]
+ scanchain_041/module_data_out[5] scanchain_041/module_data_out[6] scanchain_041/module_data_out[7]
+ scanchain_041/scan_select_in scanchain_042/scan_select_in vccd1 vssd1 scanchain
Xuser_module_361728533238569985_190 scanchain_190/module_data_in[0] scanchain_190/module_data_in[1]
+ scanchain_190/module_data_in[2] scanchain_190/module_data_in[3] scanchain_190/module_data_in[4]
+ scanchain_190/module_data_in[5] scanchain_190/module_data_in[6] scanchain_190/module_data_in[7]
+ scanchain_190/module_data_out[0] scanchain_190/module_data_out[1] scanchain_190/module_data_out[2]
+ scanchain_190/module_data_out[3] scanchain_190/module_data_out[4] scanchain_190/module_data_out[5]
+ scanchain_190/module_data_out[6] scanchain_190/module_data_out[7] vccd1 vssd1 user_module_361728533238569985
Xscanchain_052 scanchain_052/clk_in scanchain_053/clk_in scanchain_052/data_in scanchain_053/data_in
+ scanchain_052/latch_enable_in scanchain_053/latch_enable_in scanchain_052/module_data_in[0]
+ scanchain_052/module_data_in[1] scanchain_052/module_data_in[2] scanchain_052/module_data_in[3]
+ scanchain_052/module_data_in[4] scanchain_052/module_data_in[5] scanchain_052/module_data_in[6]
+ scanchain_052/module_data_in[7] scanchain_052/module_data_out[0] scanchain_052/module_data_out[1]
+ scanchain_052/module_data_out[2] scanchain_052/module_data_out[3] scanchain_052/module_data_out[4]
+ scanchain_052/module_data_out[5] scanchain_052/module_data_out[6] scanchain_052/module_data_out[7]
+ scanchain_052/scan_select_in scanchain_053/scan_select_in vccd1 vssd1 scanchain
Xscanchain_074 scanchain_074/clk_in scanchain_075/clk_in scanchain_074/data_in scanchain_075/data_in
+ scanchain_074/latch_enable_in scanchain_075/latch_enable_in scanchain_074/module_data_in[0]
+ scanchain_074/module_data_in[1] scanchain_074/module_data_in[2] scanchain_074/module_data_in[3]
+ scanchain_074/module_data_in[4] scanchain_074/module_data_in[5] scanchain_074/module_data_in[6]
+ scanchain_074/module_data_in[7] scanchain_074/module_data_out[0] scanchain_074/module_data_out[1]
+ scanchain_074/module_data_out[2] scanchain_074/module_data_out[3] scanchain_074/module_data_out[4]
+ scanchain_074/module_data_out[5] scanchain_074/module_data_out[6] scanchain_074/module_data_out[7]
+ scanchain_074/scan_select_in scanchain_075/scan_select_in vccd1 vssd1 scanchain
Xscanchain_063 scanchain_063/clk_in scanchain_064/clk_in scanchain_063/data_in scanchain_064/data_in
+ scanchain_063/latch_enable_in scanchain_064/latch_enable_in scanchain_063/module_data_in[0]
+ scanchain_063/module_data_in[1] scanchain_063/module_data_in[2] scanchain_063/module_data_in[3]
+ scanchain_063/module_data_in[4] scanchain_063/module_data_in[5] scanchain_063/module_data_in[6]
+ scanchain_063/module_data_in[7] scanchain_063/module_data_out[0] scanchain_063/module_data_out[1]
+ scanchain_063/module_data_out[2] scanchain_063/module_data_out[3] scanchain_063/module_data_out[4]
+ scanchain_063/module_data_out[5] scanchain_063/module_data_out[6] scanchain_063/module_data_out[7]
+ scanchain_063/scan_select_in scanchain_064/scan_select_in vccd1 vssd1 scanchain
Xscanchain_085 scanchain_085/clk_in scanchain_086/clk_in scanchain_085/data_in scanchain_086/data_in
+ scanchain_085/latch_enable_in scanchain_086/latch_enable_in scanchain_085/module_data_in[0]
+ scanchain_085/module_data_in[1] scanchain_085/module_data_in[2] scanchain_085/module_data_in[3]
+ scanchain_085/module_data_in[4] scanchain_085/module_data_in[5] scanchain_085/module_data_in[6]
+ scanchain_085/module_data_in[7] scanchain_085/module_data_out[0] scanchain_085/module_data_out[1]
+ scanchain_085/module_data_out[2] scanchain_085/module_data_out[3] scanchain_085/module_data_out[4]
+ scanchain_085/module_data_out[5] scanchain_085/module_data_out[6] scanchain_085/module_data_out[7]
+ scanchain_085/scan_select_in scanchain_086/scan_select_in vccd1 vssd1 scanchain
Xscanchain_096 scanchain_096/clk_in scanchain_097/clk_in scanchain_096/data_in scanchain_097/data_in
+ scanchain_096/latch_enable_in scanchain_097/latch_enable_in scanchain_096/module_data_in[0]
+ scanchain_096/module_data_in[1] scanchain_096/module_data_in[2] scanchain_096/module_data_in[3]
+ scanchain_096/module_data_in[4] scanchain_096/module_data_in[5] scanchain_096/module_data_in[6]
+ scanchain_096/module_data_in[7] scanchain_096/module_data_out[0] scanchain_096/module_data_out[1]
+ scanchain_096/module_data_out[2] scanchain_096/module_data_out[3] scanchain_096/module_data_out[4]
+ scanchain_096/module_data_out[5] scanchain_096/module_data_out[6] scanchain_096/module_data_out[7]
+ scanchain_096/scan_select_in scanchain_097/scan_select_in vccd1 vssd1 scanchain
Xuser_module_360745091952588801_032 scanchain_032/module_data_in[0] scanchain_032/module_data_in[1]
+ scanchain_032/module_data_in[2] scanchain_032/module_data_in[3] scanchain_032/module_data_in[4]
+ scanchain_032/module_data_in[5] scanchain_032/module_data_in[6] scanchain_032/module_data_in[7]
+ scanchain_032/module_data_out[0] scanchain_032/module_data_out[1] scanchain_032/module_data_out[2]
+ scanchain_032/module_data_out[3] scanchain_032/module_data_out[4] scanchain_032/module_data_out[5]
+ scanchain_032/module_data_out[6] scanchain_032/module_data_out[7] vccd1 vssd1 user_module_360745091952588801
Xuser_module_358370685977079809_051 scanchain_051/module_data_in[0] scanchain_051/module_data_in[1]
+ scanchain_051/module_data_in[2] scanchain_051/module_data_in[3] scanchain_051/module_data_in[4]
+ scanchain_051/module_data_in[5] scanchain_051/module_data_in[6] scanchain_051/module_data_in[7]
+ scanchain_051/module_data_out[0] scanchain_051/module_data_out[1] scanchain_051/module_data_out[2]
+ scanchain_051/module_data_out[3] scanchain_051/module_data_out[4] scanchain_051/module_data_out[5]
+ scanchain_051/module_data_out[6] scanchain_051/module_data_out[7] vccd1 vssd1 user_module_358370685977079809
Xuser_module_362675777226104833_062 scanchain_062/module_data_in[0] scanchain_062/module_data_in[1]
+ scanchain_062/module_data_in[2] scanchain_062/module_data_in[3] scanchain_062/module_data_in[4]
+ scanchain_062/module_data_in[5] scanchain_062/module_data_in[6] scanchain_062/module_data_in[7]
+ scanchain_062/module_data_out[0] scanchain_062/module_data_out[1] scanchain_062/module_data_out[2]
+ scanchain_062/module_data_out[3] scanchain_062/module_data_out[4] scanchain_062/module_data_out[5]
+ scanchain_062/module_data_out[6] scanchain_062/module_data_out[7] vccd1 vssd1 user_module_362675777226104833
Xscanchain_223 scanchain_223/clk_in scanchain_224/clk_in scanchain_223/data_in scanchain_224/data_in
+ scanchain_223/latch_enable_in scanchain_224/latch_enable_in scanchain_223/module_data_in[0]
+ scanchain_223/module_data_in[1] scanchain_223/module_data_in[2] scanchain_223/module_data_in[3]
+ scanchain_223/module_data_in[4] scanchain_223/module_data_in[5] scanchain_223/module_data_in[6]
+ scanchain_223/module_data_in[7] scanchain_223/module_data_out[0] scanchain_223/module_data_out[1]
+ scanchain_223/module_data_out[2] scanchain_223/module_data_out[3] scanchain_223/module_data_out[4]
+ scanchain_223/module_data_out[5] scanchain_223/module_data_out[6] scanchain_223/module_data_out[7]
+ scanchain_223/scan_select_in scanchain_224/scan_select_in vccd1 vssd1 scanchain
Xscanchain_234 scanchain_234/clk_in scanchain_235/clk_in scanchain_234/data_in scanchain_235/data_in
+ scanchain_234/latch_enable_in scanchain_235/latch_enable_in scanchain_234/module_data_in[0]
+ scanchain_234/module_data_in[1] scanchain_234/module_data_in[2] scanchain_234/module_data_in[3]
+ scanchain_234/module_data_in[4] scanchain_234/module_data_in[5] scanchain_234/module_data_in[6]
+ scanchain_234/module_data_in[7] scanchain_234/module_data_out[0] scanchain_234/module_data_out[1]
+ scanchain_234/module_data_out[2] scanchain_234/module_data_out[3] scanchain_234/module_data_out[4]
+ scanchain_234/module_data_out[5] scanchain_234/module_data_out[6] scanchain_234/module_data_out[7]
+ scanchain_234/scan_select_in scanchain_235/scan_select_in vccd1 vssd1 scanchain
Xscanchain_245 scanchain_245/clk_in scanchain_246/clk_in scanchain_245/data_in scanchain_246/data_in
+ scanchain_245/latch_enable_in scanchain_246/latch_enable_in scanchain_245/module_data_in[0]
+ scanchain_245/module_data_in[1] scanchain_245/module_data_in[2] scanchain_245/module_data_in[3]
+ scanchain_245/module_data_in[4] scanchain_245/module_data_in[5] scanchain_245/module_data_in[6]
+ scanchain_245/module_data_in[7] scanchain_245/module_data_out[0] scanchain_245/module_data_out[1]
+ scanchain_245/module_data_out[2] scanchain_245/module_data_out[3] scanchain_245/module_data_out[4]
+ scanchain_245/module_data_out[5] scanchain_245/module_data_out[6] scanchain_245/module_data_out[7]
+ scanchain_245/scan_select_in scanchain_246/scan_select_in vccd1 vssd1 scanchain
Xscanchain_212 scanchain_212/clk_in scanchain_213/clk_in scanchain_212/data_in scanchain_213/data_in
+ scanchain_212/latch_enable_in scanchain_213/latch_enable_in scanchain_212/module_data_in[0]
+ scanchain_212/module_data_in[1] scanchain_212/module_data_in[2] scanchain_212/module_data_in[3]
+ scanchain_212/module_data_in[4] scanchain_212/module_data_in[5] scanchain_212/module_data_in[6]
+ scanchain_212/module_data_in[7] scanchain_212/module_data_out[0] scanchain_212/module_data_out[1]
+ scanchain_212/module_data_out[2] scanchain_212/module_data_out[3] scanchain_212/module_data_out[4]
+ scanchain_212/module_data_out[5] scanchain_212/module_data_out[6] scanchain_212/module_data_out[7]
+ scanchain_212/scan_select_in scanchain_213/scan_select_in vccd1 vssd1 scanchain
Xscanchain_201 scanchain_201/clk_in scanchain_202/clk_in scanchain_201/data_in scanchain_202/data_in
+ scanchain_201/latch_enable_in scanchain_202/latch_enable_in scanchain_201/module_data_in[0]
+ scanchain_201/module_data_in[1] scanchain_201/module_data_in[2] scanchain_201/module_data_in[3]
+ scanchain_201/module_data_in[4] scanchain_201/module_data_in[5] scanchain_201/module_data_in[6]
+ scanchain_201/module_data_in[7] scanchain_201/module_data_out[0] scanchain_201/module_data_out[1]
+ scanchain_201/module_data_out[2] scanchain_201/module_data_out[3] scanchain_201/module_data_out[4]
+ scanchain_201/module_data_out[5] scanchain_201/module_data_out[6] scanchain_201/module_data_out[7]
+ scanchain_201/scan_select_in scanchain_202/scan_select_in vccd1 vssd1 scanchain
Xscanchain_097 scanchain_097/clk_in scanchain_098/clk_in scanchain_097/data_in scanchain_098/data_in
+ scanchain_097/latch_enable_in scanchain_098/latch_enable_in scanchain_097/module_data_in[0]
+ scanchain_097/module_data_in[1] scanchain_097/module_data_in[2] scanchain_097/module_data_in[3]
+ scanchain_097/module_data_in[4] scanchain_097/module_data_in[5] scanchain_097/module_data_in[6]
+ scanchain_097/module_data_in[7] scanchain_097/module_data_out[0] scanchain_097/module_data_out[1]
+ scanchain_097/module_data_out[2] scanchain_097/module_data_out[3] scanchain_097/module_data_out[4]
+ scanchain_097/module_data_out[5] scanchain_097/module_data_out[6] scanchain_097/module_data_out[7]
+ scanchain_097/scan_select_in scanchain_098/scan_select_in vccd1 vssd1 scanchain
Xscanchain_020 scanchain_020/clk_in scanchain_021/clk_in scanchain_020/data_in scanchain_021/data_in
+ scanchain_020/latch_enable_in scanchain_021/latch_enable_in scanchain_020/module_data_in[0]
+ scanchain_020/module_data_in[1] scanchain_020/module_data_in[2] scanchain_020/module_data_in[3]
+ scanchain_020/module_data_in[4] scanchain_020/module_data_in[5] scanchain_020/module_data_in[6]
+ scanchain_020/module_data_in[7] scanchain_020/module_data_out[0] scanchain_020/module_data_out[1]
+ scanchain_020/module_data_out[2] scanchain_020/module_data_out[3] scanchain_020/module_data_out[4]
+ scanchain_020/module_data_out[5] scanchain_020/module_data_out[6] scanchain_020/module_data_out[7]
+ scanchain_020/scan_select_in scanchain_021/scan_select_in vccd1 vssd1 scanchain
Xscanchain_031 scanchain_031/clk_in scanchain_032/clk_in scanchain_031/data_in scanchain_032/data_in
+ scanchain_031/latch_enable_in scanchain_032/latch_enable_in scanchain_031/module_data_in[0]
+ scanchain_031/module_data_in[1] scanchain_031/module_data_in[2] scanchain_031/module_data_in[3]
+ scanchain_031/module_data_in[4] scanchain_031/module_data_in[5] scanchain_031/module_data_in[6]
+ scanchain_031/module_data_in[7] scanchain_031/module_data_out[0] scanchain_031/module_data_out[1]
+ scanchain_031/module_data_out[2] scanchain_031/module_data_out[3] scanchain_031/module_data_out[4]
+ scanchain_031/module_data_out[5] scanchain_031/module_data_out[6] scanchain_031/module_data_out[7]
+ scanchain_031/scan_select_in scanchain_032/scan_select_in vccd1 vssd1 scanchain
Xscanchain_042 scanchain_042/clk_in scanchain_043/clk_in scanchain_042/data_in scanchain_043/data_in
+ scanchain_042/latch_enable_in scanchain_043/latch_enable_in jordan336_toy_cpu_042/io_in[0]
+ jordan336_toy_cpu_042/io_in[1] jordan336_toy_cpu_042/io_in[2] jordan336_toy_cpu_042/io_in[3]
+ jordan336_toy_cpu_042/io_in[4] jordan336_toy_cpu_042/io_in[5] jordan336_toy_cpu_042/io_in[6]
+ jordan336_toy_cpu_042/io_in[7] jordan336_toy_cpu_042/io_out[0] jordan336_toy_cpu_042/io_out[1]
+ jordan336_toy_cpu_042/io_out[2] jordan336_toy_cpu_042/io_out[3] jordan336_toy_cpu_042/io_out[4]
+ jordan336_toy_cpu_042/io_out[5] jordan336_toy_cpu_042/io_out[6] jordan336_toy_cpu_042/io_out[7]
+ scanchain_042/scan_select_in scanchain_043/scan_select_in vccd1 vssd1 scanchain
Xscanchain_053 scanchain_053/clk_in scanchain_054/clk_in scanchain_053/data_in scanchain_054/data_in
+ scanchain_053/latch_enable_in scanchain_054/latch_enable_in scanchain_053/module_data_in[0]
+ scanchain_053/module_data_in[1] scanchain_053/module_data_in[2] scanchain_053/module_data_in[3]
+ scanchain_053/module_data_in[4] scanchain_053/module_data_in[5] scanchain_053/module_data_in[6]
+ scanchain_053/module_data_in[7] scanchain_053/module_data_out[0] scanchain_053/module_data_out[1]
+ scanchain_053/module_data_out[2] scanchain_053/module_data_out[3] scanchain_053/module_data_out[4]
+ scanchain_053/module_data_out[5] scanchain_053/module_data_out[6] scanchain_053/module_data_out[7]
+ scanchain_053/scan_select_in scanchain_054/scan_select_in vccd1 vssd1 scanchain
Xuser_module_361728533238569985_191 scanchain_191/module_data_in[0] scanchain_191/module_data_in[1]
+ scanchain_191/module_data_in[2] scanchain_191/module_data_in[3] scanchain_191/module_data_in[4]
+ scanchain_191/module_data_in[5] scanchain_191/module_data_in[6] scanchain_191/module_data_in[7]
+ scanchain_191/module_data_out[0] scanchain_191/module_data_out[1] scanchain_191/module_data_out[2]
+ scanchain_191/module_data_out[3] scanchain_191/module_data_out[4] scanchain_191/module_data_out[5]
+ scanchain_191/module_data_out[6] scanchain_191/module_data_out[7] vccd1 vssd1 user_module_361728533238569985
Xuser_module_361728533238569985_180 scanchain_180/module_data_in[0] scanchain_180/module_data_in[1]
+ scanchain_180/module_data_in[2] scanchain_180/module_data_in[3] scanchain_180/module_data_in[4]
+ scanchain_180/module_data_in[5] scanchain_180/module_data_in[6] scanchain_180/module_data_in[7]
+ scanchain_180/module_data_out[0] scanchain_180/module_data_out[1] scanchain_180/module_data_out[2]
+ scanchain_180/module_data_out[3] scanchain_180/module_data_out[4] scanchain_180/module_data_out[5]
+ scanchain_180/module_data_out[6] scanchain_180/module_data_out[7] vccd1 vssd1 user_module_361728533238569985
Xscanchain_064 scanchain_064/clk_in scanchain_065/clk_in scanchain_064/data_in scanchain_065/data_in
+ scanchain_064/latch_enable_in scanchain_065/latch_enable_in scanchain_064/module_data_in[0]
+ scanchain_064/module_data_in[1] scanchain_064/module_data_in[2] scanchain_064/module_data_in[3]
+ scanchain_064/module_data_in[4] scanchain_064/module_data_in[5] scanchain_064/module_data_in[6]
+ scanchain_064/module_data_in[7] scanchain_064/module_data_out[0] scanchain_064/module_data_out[1]
+ scanchain_064/module_data_out[2] scanchain_064/module_data_out[3] scanchain_064/module_data_out[4]
+ scanchain_064/module_data_out[5] scanchain_064/module_data_out[6] scanchain_064/module_data_out[7]
+ scanchain_064/scan_select_in scanchain_065/scan_select_in vccd1 vssd1 scanchain
Xscanchain_075 scanchain_075/clk_in scanchain_076/clk_in scanchain_075/data_in scanchain_076/data_in
+ scanchain_075/latch_enable_in scanchain_076/latch_enable_in scanchain_075/module_data_in[0]
+ scanchain_075/module_data_in[1] scanchain_075/module_data_in[2] scanchain_075/module_data_in[3]
+ scanchain_075/module_data_in[4] scanchain_075/module_data_in[5] scanchain_075/module_data_in[6]
+ scanchain_075/module_data_in[7] scanchain_075/module_data_out[0] scanchain_075/module_data_out[1]
+ scanchain_075/module_data_out[2] scanchain_075/module_data_out[3] scanchain_075/module_data_out[4]
+ scanchain_075/module_data_out[5] scanchain_075/module_data_out[6] scanchain_075/module_data_out[7]
+ scanchain_075/scan_select_in scanchain_076/scan_select_in vccd1 vssd1 scanchain
Xscanchain_086 scanchain_086/clk_in scanchain_087/clk_in scanchain_086/data_in scanchain_087/data_in
+ scanchain_086/latch_enable_in scanchain_087/latch_enable_in scanchain_086/module_data_in[0]
+ scanchain_086/module_data_in[1] scanchain_086/module_data_in[2] scanchain_086/module_data_in[3]
+ scanchain_086/module_data_in[4] scanchain_086/module_data_in[5] scanchain_086/module_data_in[6]
+ scanchain_086/module_data_in[7] scanchain_086/module_data_out[0] scanchain_086/module_data_out[1]
+ scanchain_086/module_data_out[2] scanchain_086/module_data_out[3] scanchain_086/module_data_out[4]
+ scanchain_086/module_data_out[5] scanchain_086/module_data_out[6] scanchain_086/module_data_out[7]
+ scanchain_086/scan_select_in scanchain_087/scan_select_in vccd1 vssd1 scanchain
Xmeiniki_pi_003 meiniki_pi_003/io_in[0] meiniki_pi_003/io_in[1] meiniki_pi_003/io_in[2]
+ meiniki_pi_003/io_in[3] meiniki_pi_003/io_in[4] meiniki_pi_003/io_in[5] meiniki_pi_003/io_in[6]
+ meiniki_pi_003/io_in[7] meiniki_pi_003/io_out[0] meiniki_pi_003/io_out[1] meiniki_pi_003/io_out[2]
+ meiniki_pi_003/io_out[3] meiniki_pi_003/io_out[4] meiniki_pi_003/io_out[5] meiniki_pi_003/io_out[6]
+ meiniki_pi_003/io_out[7] vccd1 vssd1 meiniki_pi
Xuser_module_347417602591556180_085 scanchain_085/module_data_in[0] scanchain_085/module_data_in[1]
+ scanchain_085/module_data_in[2] scanchain_085/module_data_in[3] scanchain_085/module_data_in[4]
+ scanchain_085/module_data_in[5] scanchain_085/module_data_in[6] scanchain_085/module_data_in[7]
+ scanchain_085/module_data_out[0] scanchain_085/module_data_out[1] scanchain_085/module_data_out[2]
+ scanchain_085/module_data_out[3] scanchain_085/module_data_out[4] scanchain_085/module_data_out[5]
+ scanchain_085/module_data_out[6] scanchain_085/module_data_out[7] vccd1 vssd1 user_module_347417602591556180
Xseven_segment_seconds_055 scanchain_055/module_data_in[0] scanchain_055/module_data_in[1]
+ scanchain_055/module_data_in[2] scanchain_055/module_data_in[3] scanchain_055/module_data_in[4]
+ scanchain_055/module_data_in[5] scanchain_055/module_data_in[6] scanchain_055/module_data_in[7]
+ scanchain_055/module_data_out[0] scanchain_055/module_data_out[1] scanchain_055/module_data_out[2]
+ scanchain_055/module_data_out[3] scanchain_055/module_data_out[4] scanchain_055/module_data_out[5]
+ scanchain_055/module_data_out[6] scanchain_055/module_data_out[7] vccd1 vssd1 seven_segment_seconds
Xtomkeddie_top_tto_a_028 scanchain_028/module_data_in[0] scanchain_028/module_data_in[1]
+ scanchain_028/module_data_in[2] scanchain_028/module_data_in[3] scanchain_028/module_data_in[4]
+ scanchain_028/module_data_in[5] scanchain_028/module_data_in[6] scanchain_028/module_data_in[7]
+ scanchain_028/module_data_out[0] scanchain_028/module_data_out[1] scanchain_028/module_data_out[2]
+ scanchain_028/module_data_out[3] scanchain_028/module_data_out[4] scanchain_028/module_data_out[5]
+ scanchain_028/module_data_out[6] scanchain_028/module_data_out[7] vccd1 vssd1 tomkeddie_top_tto_a
Xdiferential_rvb1_022 diferential_rvb1_022/io_in[0] diferential_rvb1_022/io_in[1]
+ diferential_rvb1_022/io_in[2] diferential_rvb1_022/io_in[3] diferential_rvb1_022/io_in[4]
+ diferential_rvb1_022/io_in[5] diferential_rvb1_022/io_in[6] diferential_rvb1_022/io_in[7]
+ diferential_rvb1_022/io_out[0] diferential_rvb1_022/io_out[1] diferential_rvb1_022/io_out[2]
+ diferential_rvb1_022/io_out[3] diferential_rvb1_022/io_out[4] diferential_rvb1_022/io_out[5]
+ diferential_rvb1_022/io_out[6] diferential_rvb1_022/io_out[7] vccd1 vssd1 diferential_rvb1
Xscanchain_224 scanchain_224/clk_in scanchain_225/clk_in scanchain_224/data_in scanchain_225/data_in
+ scanchain_224/latch_enable_in scanchain_225/latch_enable_in scanchain_224/module_data_in[0]
+ scanchain_224/module_data_in[1] scanchain_224/module_data_in[2] scanchain_224/module_data_in[3]
+ scanchain_224/module_data_in[4] scanchain_224/module_data_in[5] scanchain_224/module_data_in[6]
+ scanchain_224/module_data_in[7] scanchain_224/module_data_out[0] scanchain_224/module_data_out[1]
+ scanchain_224/module_data_out[2] scanchain_224/module_data_out[3] scanchain_224/module_data_out[4]
+ scanchain_224/module_data_out[5] scanchain_224/module_data_out[6] scanchain_224/module_data_out[7]
+ scanchain_224/scan_select_in scanchain_225/scan_select_in vccd1 vssd1 scanchain
Xscanchain_235 scanchain_235/clk_in scanchain_236/clk_in scanchain_235/data_in scanchain_236/data_in
+ scanchain_235/latch_enable_in scanchain_236/latch_enable_in scanchain_235/module_data_in[0]
+ scanchain_235/module_data_in[1] scanchain_235/module_data_in[2] scanchain_235/module_data_in[3]
+ scanchain_235/module_data_in[4] scanchain_235/module_data_in[5] scanchain_235/module_data_in[6]
+ scanchain_235/module_data_in[7] scanchain_235/module_data_out[0] scanchain_235/module_data_out[1]
+ scanchain_235/module_data_out[2] scanchain_235/module_data_out[3] scanchain_235/module_data_out[4]
+ scanchain_235/module_data_out[5] scanchain_235/module_data_out[6] scanchain_235/module_data_out[7]
+ scanchain_235/scan_select_in scanchain_236/scan_select_in vccd1 vssd1 scanchain
Xscanchain_246 scanchain_246/clk_in scanchain_247/clk_in scanchain_246/data_in scanchain_247/data_in
+ scanchain_246/latch_enable_in scanchain_247/latch_enable_in scanchain_246/module_data_in[0]
+ scanchain_246/module_data_in[1] scanchain_246/module_data_in[2] scanchain_246/module_data_in[3]
+ scanchain_246/module_data_in[4] scanchain_246/module_data_in[5] scanchain_246/module_data_in[6]
+ scanchain_246/module_data_in[7] scanchain_246/module_data_out[0] scanchain_246/module_data_out[1]
+ scanchain_246/module_data_out[2] scanchain_246/module_data_out[3] scanchain_246/module_data_out[4]
+ scanchain_246/module_data_out[5] scanchain_246/module_data_out[6] scanchain_246/module_data_out[7]
+ scanchain_246/scan_select_in scanchain_247/scan_select_in vccd1 vssd1 scanchain
Xscanchain_213 scanchain_213/clk_in scanchain_214/clk_in scanchain_213/data_in scanchain_214/data_in
+ scanchain_213/latch_enable_in scanchain_214/latch_enable_in scanchain_213/module_data_in[0]
+ scanchain_213/module_data_in[1] scanchain_213/module_data_in[2] scanchain_213/module_data_in[3]
+ scanchain_213/module_data_in[4] scanchain_213/module_data_in[5] scanchain_213/module_data_in[6]
+ scanchain_213/module_data_in[7] scanchain_213/module_data_out[0] scanchain_213/module_data_out[1]
+ scanchain_213/module_data_out[2] scanchain_213/module_data_out[3] scanchain_213/module_data_out[4]
+ scanchain_213/module_data_out[5] scanchain_213/module_data_out[6] scanchain_213/module_data_out[7]
+ scanchain_213/scan_select_in scanchain_214/scan_select_in vccd1 vssd1 scanchain
Xscanchain_202 scanchain_202/clk_in scanchain_203/clk_in scanchain_202/data_in scanchain_203/data_in
+ scanchain_202/latch_enable_in scanchain_203/latch_enable_in scanchain_202/module_data_in[0]
+ scanchain_202/module_data_in[1] scanchain_202/module_data_in[2] scanchain_202/module_data_in[3]
+ scanchain_202/module_data_in[4] scanchain_202/module_data_in[5] scanchain_202/module_data_in[6]
+ scanchain_202/module_data_in[7] scanchain_202/module_data_out[0] scanchain_202/module_data_out[1]
+ scanchain_202/module_data_out[2] scanchain_202/module_data_out[3] scanchain_202/module_data_out[4]
+ scanchain_202/module_data_out[5] scanchain_202/module_data_out[6] scanchain_202/module_data_out[7]
+ scanchain_202/scan_select_in scanchain_203/scan_select_in vccd1 vssd1 scanchain
Xscanchain_098 scanchain_098/clk_in scanchain_099/clk_in scanchain_098/data_in scanchain_099/data_in
+ scanchain_098/latch_enable_in scanchain_099/latch_enable_in scanchain_098/module_data_in[0]
+ scanchain_098/module_data_in[1] scanchain_098/module_data_in[2] scanchain_098/module_data_in[3]
+ scanchain_098/module_data_in[4] scanchain_098/module_data_in[5] scanchain_098/module_data_in[6]
+ scanchain_098/module_data_in[7] scanchain_098/module_data_out[0] scanchain_098/module_data_out[1]
+ scanchain_098/module_data_out[2] scanchain_098/module_data_out[3] scanchain_098/module_data_out[4]
+ scanchain_098/module_data_out[5] scanchain_098/module_data_out[6] scanchain_098/module_data_out[7]
+ scanchain_098/scan_select_in scanchain_099/scan_select_in vccd1 vssd1 scanchain
Xscanchain_010 scanchain_010/clk_in scanchain_011/clk_in scanchain_010/data_in scanchain_011/data_in
+ scanchain_010/latch_enable_in scanchain_011/latch_enable_in scanchain_010/module_data_in[0]
+ scanchain_010/module_data_in[1] scanchain_010/module_data_in[2] scanchain_010/module_data_in[3]
+ scanchain_010/module_data_in[4] scanchain_010/module_data_in[5] scanchain_010/module_data_in[6]
+ scanchain_010/module_data_in[7] scanchain_010/module_data_out[0] scanchain_010/module_data_out[1]
+ scanchain_010/module_data_out[2] scanchain_010/module_data_out[3] scanchain_010/module_data_out[4]
+ scanchain_010/module_data_out[5] scanchain_010/module_data_out[6] scanchain_010/module_data_out[7]
+ scanchain_010/scan_select_in scanchain_011/scan_select_in vccd1 vssd1 scanchain
Xscanchain_021 scanchain_021/clk_in scanchain_022/clk_in scanchain_021/data_in scanchain_022/data_in
+ scanchain_021/latch_enable_in scanchain_022/latch_enable_in scanchain_021/module_data_in[0]
+ scanchain_021/module_data_in[1] scanchain_021/module_data_in[2] scanchain_021/module_data_in[3]
+ scanchain_021/module_data_in[4] scanchain_021/module_data_in[5] scanchain_021/module_data_in[6]
+ scanchain_021/module_data_in[7] scanchain_021/module_data_out[0] scanchain_021/module_data_out[1]
+ scanchain_021/module_data_out[2] scanchain_021/module_data_out[3] scanchain_021/module_data_out[4]
+ scanchain_021/module_data_out[5] scanchain_021/module_data_out[6] scanchain_021/module_data_out[7]
+ scanchain_021/scan_select_in scanchain_022/scan_select_in vccd1 vssd1 scanchain
Xscanchain_032 scanchain_032/clk_in scanchain_033/clk_in scanchain_032/data_in scanchain_033/data_in
+ scanchain_032/latch_enable_in scanchain_033/latch_enable_in scanchain_032/module_data_in[0]
+ scanchain_032/module_data_in[1] scanchain_032/module_data_in[2] scanchain_032/module_data_in[3]
+ scanchain_032/module_data_in[4] scanchain_032/module_data_in[5] scanchain_032/module_data_in[6]
+ scanchain_032/module_data_in[7] scanchain_032/module_data_out[0] scanchain_032/module_data_out[1]
+ scanchain_032/module_data_out[2] scanchain_032/module_data_out[3] scanchain_032/module_data_out[4]
+ scanchain_032/module_data_out[5] scanchain_032/module_data_out[6] scanchain_032/module_data_out[7]
+ scanchain_032/scan_select_in scanchain_033/scan_select_in vccd1 vssd1 scanchain
Xscanchain_043 scanchain_043/clk_in scanchain_044/clk_in scanchain_043/data_in scanchain_044/data_in
+ scanchain_043/latch_enable_in scanchain_044/latch_enable_in dwisehart_top_043/io_in[0]
+ dwisehart_top_043/io_in[1] dwisehart_top_043/io_in[2] dwisehart_top_043/io_in[3]
+ dwisehart_top_043/io_in[4] dwisehart_top_043/io_in[5] dwisehart_top_043/io_in[6]
+ dwisehart_top_043/io_in[7] dwisehart_top_043/io_out[0] dwisehart_top_043/io_out[1]
+ dwisehart_top_043/io_out[2] dwisehart_top_043/io_out[3] dwisehart_top_043/io_out[4]
+ dwisehart_top_043/io_out[5] dwisehart_top_043/io_out[6] dwisehart_top_043/io_out[7]
+ scanchain_043/scan_select_in scanchain_044/scan_select_in vccd1 vssd1 scanchain
Xscanchain_054 scanchain_054/clk_in scanchain_055/clk_in scanchain_054/data_in scanchain_055/data_in
+ scanchain_054/latch_enable_in scanchain_055/latch_enable_in scanchain_054/module_data_in[0]
+ scanchain_054/module_data_in[1] scanchain_054/module_data_in[2] scanchain_054/module_data_in[3]
+ scanchain_054/module_data_in[4] scanchain_054/module_data_in[5] scanchain_054/module_data_in[6]
+ scanchain_054/module_data_in[7] scanchain_054/module_data_out[0] scanchain_054/module_data_out[1]
+ scanchain_054/module_data_out[2] scanchain_054/module_data_out[3] scanchain_054/module_data_out[4]
+ scanchain_054/module_data_out[5] scanchain_054/module_data_out[6] scanchain_054/module_data_out[7]
+ scanchain_054/scan_select_in scanchain_055/scan_select_in vccd1 vssd1 scanchain
Xuser_module_361728533238569985_192 scanchain_192/module_data_in[0] scanchain_192/module_data_in[1]
+ scanchain_192/module_data_in[2] scanchain_192/module_data_in[3] scanchain_192/module_data_in[4]
+ scanchain_192/module_data_in[5] scanchain_192/module_data_in[6] scanchain_192/module_data_in[7]
+ scanchain_192/module_data_out[0] scanchain_192/module_data_out[1] scanchain_192/module_data_out[2]
+ scanchain_192/module_data_out[3] scanchain_192/module_data_out[4] scanchain_192/module_data_out[5]
+ scanchain_192/module_data_out[6] scanchain_192/module_data_out[7] vccd1 vssd1 user_module_361728533238569985
Xuser_module_361728533238569985_181 scanchain_181/module_data_in[0] scanchain_181/module_data_in[1]
+ scanchain_181/module_data_in[2] scanchain_181/module_data_in[3] scanchain_181/module_data_in[4]
+ scanchain_181/module_data_in[5] scanchain_181/module_data_in[6] scanchain_181/module_data_in[7]
+ scanchain_181/module_data_out[0] scanchain_181/module_data_out[1] scanchain_181/module_data_out[2]
+ scanchain_181/module_data_out[3] scanchain_181/module_data_out[4] scanchain_181/module_data_out[5]
+ scanchain_181/module_data_out[6] scanchain_181/module_data_out[7] vccd1 vssd1 user_module_361728533238569985
Xscanchain_065 scanchain_065/clk_in scanchain_066/clk_in scanchain_065/data_in scanchain_066/data_in
+ scanchain_065/latch_enable_in scanchain_066/latch_enable_in scanchain_065/module_data_in[0]
+ scanchain_065/module_data_in[1] scanchain_065/module_data_in[2] scanchain_065/module_data_in[3]
+ scanchain_065/module_data_in[4] scanchain_065/module_data_in[5] scanchain_065/module_data_in[6]
+ scanchain_065/module_data_in[7] scanchain_065/module_data_out[0] scanchain_065/module_data_out[1]
+ scanchain_065/module_data_out[2] scanchain_065/module_data_out[3] scanchain_065/module_data_out[4]
+ scanchain_065/module_data_out[5] scanchain_065/module_data_out[6] scanchain_065/module_data_out[7]
+ scanchain_065/scan_select_in scanchain_066/scan_select_in vccd1 vssd1 scanchain
Xuser_module_361728533238569985_170 scanchain_170/module_data_in[0] scanchain_170/module_data_in[1]
+ scanchain_170/module_data_in[2] scanchain_170/module_data_in[3] scanchain_170/module_data_in[4]
+ scanchain_170/module_data_in[5] scanchain_170/module_data_in[6] scanchain_170/module_data_in[7]
+ scanchain_170/module_data_out[0] scanchain_170/module_data_out[1] scanchain_170/module_data_out[2]
+ scanchain_170/module_data_out[3] scanchain_170/module_data_out[4] scanchain_170/module_data_out[5]
+ scanchain_170/module_data_out[6] scanchain_170/module_data_out[7] vccd1 vssd1 user_module_361728533238569985
Xscanchain_076 scanchain_076/clk_in scanchain_077/clk_in scanchain_076/data_in scanchain_077/data_in
+ scanchain_076/latch_enable_in scanchain_077/latch_enable_in scanchain_076/module_data_in[0]
+ scanchain_076/module_data_in[1] scanchain_076/module_data_in[2] scanchain_076/module_data_in[3]
+ scanchain_076/module_data_in[4] scanchain_076/module_data_in[5] scanchain_076/module_data_in[6]
+ scanchain_076/module_data_in[7] scanchain_076/module_data_out[0] scanchain_076/module_data_out[1]
+ scanchain_076/module_data_out[2] scanchain_076/module_data_out[3] scanchain_076/module_data_out[4]
+ scanchain_076/module_data_out[5] scanchain_076/module_data_out[6] scanchain_076/module_data_out[7]
+ scanchain_076/scan_select_in scanchain_077/scan_select_in vccd1 vssd1 scanchain
Xscanchain_087 scanchain_087/clk_in scanchain_088/clk_in scanchain_087/data_in scanchain_088/data_in
+ scanchain_087/latch_enable_in scanchain_088/latch_enable_in scanchain_087/module_data_in[0]
+ scanchain_087/module_data_in[1] scanchain_087/module_data_in[2] scanchain_087/module_data_in[3]
+ scanchain_087/module_data_in[4] scanchain_087/module_data_in[5] scanchain_087/module_data_in[6]
+ scanchain_087/module_data_in[7] scanchain_087/module_data_out[0] scanchain_087/module_data_out[1]
+ scanchain_087/module_data_out[2] scanchain_087/module_data_out[3] scanchain_087/module_data_out[4]
+ scanchain_087/module_data_out[5] scanchain_087/module_data_out[6] scanchain_087/module_data_out[7]
+ scanchain_087/scan_select_in scanchain_088/scan_select_in vccd1 vssd1 scanchain
Xjordan336_toy_cpu_042 jordan336_toy_cpu_042/io_in[0] jordan336_toy_cpu_042/io_in[1]
+ jordan336_toy_cpu_042/io_in[2] jordan336_toy_cpu_042/io_in[3] jordan336_toy_cpu_042/io_in[4]
+ jordan336_toy_cpu_042/io_in[5] jordan336_toy_cpu_042/io_in[6] jordan336_toy_cpu_042/io_in[7]
+ jordan336_toy_cpu_042/io_out[0] jordan336_toy_cpu_042/io_out[1] jordan336_toy_cpu_042/io_out[2]
+ jordan336_toy_cpu_042/io_out[3] jordan336_toy_cpu_042/io_out[4] jordan336_toy_cpu_042/io_out[5]
+ jordan336_toy_cpu_042/io_out[6] jordan336_toy_cpu_042/io_out[7] vccd1 vssd1 jordan336_toy_cpu
Xknight_rider_KolosKoblasz_005 scanchain_005/module_data_in[0] scanchain_005/module_data_in[1]
+ scanchain_005/module_data_in[2] scanchain_005/module_data_in[3] scanchain_005/module_data_in[4]
+ scanchain_005/module_data_in[5] scanchain_005/module_data_in[6] scanchain_005/module_data_in[7]
+ scanchain_005/module_data_out[0] scanchain_005/module_data_out[1] scanchain_005/module_data_out[2]
+ scanchain_005/module_data_out[3] scanchain_005/module_data_out[4] scanchain_005/module_data_out[5]
+ scanchain_005/module_data_out[6] scanchain_005/module_data_out[7] vccd1 vssd1 knight_rider_KolosKoblasz
Xscanchain_225 scanchain_225/clk_in scanchain_226/clk_in scanchain_225/data_in scanchain_226/data_in
+ scanchain_225/latch_enable_in scanchain_226/latch_enable_in scanchain_225/module_data_in[0]
+ scanchain_225/module_data_in[1] scanchain_225/module_data_in[2] scanchain_225/module_data_in[3]
+ scanchain_225/module_data_in[4] scanchain_225/module_data_in[5] scanchain_225/module_data_in[6]
+ scanchain_225/module_data_in[7] scanchain_225/module_data_out[0] scanchain_225/module_data_out[1]
+ scanchain_225/module_data_out[2] scanchain_225/module_data_out[3] scanchain_225/module_data_out[4]
+ scanchain_225/module_data_out[5] scanchain_225/module_data_out[6] scanchain_225/module_data_out[7]
+ scanchain_225/scan_select_in scanchain_226/scan_select_in vccd1 vssd1 scanchain
Xscanchain_236 scanchain_236/clk_in scanchain_237/clk_in scanchain_236/data_in scanchain_237/data_in
+ scanchain_236/latch_enable_in scanchain_237/latch_enable_in scanchain_236/module_data_in[0]
+ scanchain_236/module_data_in[1] scanchain_236/module_data_in[2] scanchain_236/module_data_in[3]
+ scanchain_236/module_data_in[4] scanchain_236/module_data_in[5] scanchain_236/module_data_in[6]
+ scanchain_236/module_data_in[7] scanchain_236/module_data_out[0] scanchain_236/module_data_out[1]
+ scanchain_236/module_data_out[2] scanchain_236/module_data_out[3] scanchain_236/module_data_out[4]
+ scanchain_236/module_data_out[5] scanchain_236/module_data_out[6] scanchain_236/module_data_out[7]
+ scanchain_236/scan_select_in scanchain_237/scan_select_in vccd1 vssd1 scanchain
Xscanchain_247 scanchain_247/clk_in scanchain_248/clk_in scanchain_247/data_in scanchain_248/data_in
+ scanchain_247/latch_enable_in scanchain_248/latch_enable_in scanchain_247/module_data_in[0]
+ scanchain_247/module_data_in[1] scanchain_247/module_data_in[2] scanchain_247/module_data_in[3]
+ scanchain_247/module_data_in[4] scanchain_247/module_data_in[5] scanchain_247/module_data_in[6]
+ scanchain_247/module_data_in[7] scanchain_247/module_data_out[0] scanchain_247/module_data_out[1]
+ scanchain_247/module_data_out[2] scanchain_247/module_data_out[3] scanchain_247/module_data_out[4]
+ scanchain_247/module_data_out[5] scanchain_247/module_data_out[6] scanchain_247/module_data_out[7]
+ scanchain_247/scan_select_in scanchain_248/scan_select_in vccd1 vssd1 scanchain
Xscanchain_214 scanchain_214/clk_in scanchain_215/clk_in scanchain_214/data_in scanchain_215/data_in
+ scanchain_214/latch_enable_in scanchain_215/latch_enable_in scanchain_214/module_data_in[0]
+ scanchain_214/module_data_in[1] scanchain_214/module_data_in[2] scanchain_214/module_data_in[3]
+ scanchain_214/module_data_in[4] scanchain_214/module_data_in[5] scanchain_214/module_data_in[6]
+ scanchain_214/module_data_in[7] scanchain_214/module_data_out[0] scanchain_214/module_data_out[1]
+ scanchain_214/module_data_out[2] scanchain_214/module_data_out[3] scanchain_214/module_data_out[4]
+ scanchain_214/module_data_out[5] scanchain_214/module_data_out[6] scanchain_214/module_data_out[7]
+ scanchain_214/scan_select_in scanchain_215/scan_select_in vccd1 vssd1 scanchain
Xscanchain_203 scanchain_203/clk_in scanchain_204/clk_in scanchain_203/data_in scanchain_204/data_in
+ scanchain_203/latch_enable_in scanchain_204/latch_enable_in scanchain_203/module_data_in[0]
+ scanchain_203/module_data_in[1] scanchain_203/module_data_in[2] scanchain_203/module_data_in[3]
+ scanchain_203/module_data_in[4] scanchain_203/module_data_in[5] scanchain_203/module_data_in[6]
+ scanchain_203/module_data_in[7] scanchain_203/module_data_out[0] scanchain_203/module_data_out[1]
+ scanchain_203/module_data_out[2] scanchain_203/module_data_out[3] scanchain_203/module_data_out[4]
+ scanchain_203/module_data_out[5] scanchain_203/module_data_out[6] scanchain_203/module_data_out[7]
+ scanchain_203/scan_select_in scanchain_204/scan_select_in vccd1 vssd1 scanchain
Xscanchain_099 scanchain_099/clk_in scanchain_100/clk_in scanchain_099/data_in scanchain_100/data_in
+ scanchain_099/latch_enable_in scanchain_100/latch_enable_in scanchain_099/module_data_in[0]
+ scanchain_099/module_data_in[1] scanchain_099/module_data_in[2] scanchain_099/module_data_in[3]
+ scanchain_099/module_data_in[4] scanchain_099/module_data_in[5] scanchain_099/module_data_in[6]
+ scanchain_099/module_data_in[7] scanchain_099/module_data_out[0] scanchain_099/module_data_out[1]
+ scanchain_099/module_data_out[2] scanchain_099/module_data_out[3] scanchain_099/module_data_out[4]
+ scanchain_099/module_data_out[5] scanchain_099/module_data_out[6] scanchain_099/module_data_out[7]
+ scanchain_099/scan_select_in scanchain_100/scan_select_in vccd1 vssd1 scanchain
Xscanchain_011 scanchain_011/clk_in scanchain_012/clk_in scanchain_011/data_in scanchain_012/data_in
+ scanchain_011/latch_enable_in scanchain_012/latch_enable_in scanchain_011/module_data_in[0]
+ scanchain_011/module_data_in[1] scanchain_011/module_data_in[2] scanchain_011/module_data_in[3]
+ scanchain_011/module_data_in[4] scanchain_011/module_data_in[5] scanchain_011/module_data_in[6]
+ scanchain_011/module_data_in[7] scanchain_011/module_data_out[0] scanchain_011/module_data_out[1]
+ scanchain_011/module_data_out[2] scanchain_011/module_data_out[3] scanchain_011/module_data_out[4]
+ scanchain_011/module_data_out[5] scanchain_011/module_data_out[6] scanchain_011/module_data_out[7]
+ scanchain_011/scan_select_in scanchain_012/scan_select_in vccd1 vssd1 scanchain
Xscanchain_000 scanchain_000/clk_in scanchain_001/clk_in scanchain_000/data_in scanchain_001/data_in
+ scanchain_000/latch_enable_in scanchain_001/latch_enable_in scanchain_000/module_data_in[0]
+ scanchain_000/module_data_in[1] scanchain_000/module_data_in[2] scanchain_000/module_data_in[3]
+ scanchain_000/module_data_in[4] scanchain_000/module_data_in[5] scanchain_000/module_data_in[6]
+ scanchain_000/module_data_in[7] scanchain_000/module_data_out[0] scanchain_000/module_data_out[1]
+ scanchain_000/module_data_out[2] scanchain_000/module_data_out[3] scanchain_000/module_data_out[4]
+ scanchain_000/module_data_out[5] scanchain_000/module_data_out[6] scanchain_000/module_data_out[7]
+ scan_controller/scan_select scanchain_001/scan_select_in vccd1 vssd1 scanchain
Xscanchain_022 scanchain_022/clk_in scanchain_023/clk_in scanchain_022/data_in scanchain_023/data_in
+ scanchain_022/latch_enable_in scanchain_023/latch_enable_in diferential_rvb1_022/io_in[0]
+ diferential_rvb1_022/io_in[1] diferential_rvb1_022/io_in[2] diferential_rvb1_022/io_in[3]
+ diferential_rvb1_022/io_in[4] diferential_rvb1_022/io_in[5] diferential_rvb1_022/io_in[6]
+ diferential_rvb1_022/io_in[7] diferential_rvb1_022/io_out[0] diferential_rvb1_022/io_out[1]
+ diferential_rvb1_022/io_out[2] diferential_rvb1_022/io_out[3] diferential_rvb1_022/io_out[4]
+ diferential_rvb1_022/io_out[5] diferential_rvb1_022/io_out[6] diferential_rvb1_022/io_out[7]
+ scanchain_022/scan_select_in scanchain_023/scan_select_in vccd1 vssd1 scanchain
Xscanchain_033 scanchain_033/clk_in scanchain_034/clk_in scanchain_033/data_in scanchain_034/data_in
+ scanchain_033/latch_enable_in scanchain_034/latch_enable_in scanchain_033/module_data_in[0]
+ scanchain_033/module_data_in[1] scanchain_033/module_data_in[2] scanchain_033/module_data_in[3]
+ scanchain_033/module_data_in[4] scanchain_033/module_data_in[5] scanchain_033/module_data_in[6]
+ scanchain_033/module_data_in[7] scanchain_033/module_data_out[0] scanchain_033/module_data_out[1]
+ scanchain_033/module_data_out[2] scanchain_033/module_data_out[3] scanchain_033/module_data_out[4]
+ scanchain_033/module_data_out[5] scanchain_033/module_data_out[6] scanchain_033/module_data_out[7]
+ scanchain_033/scan_select_in scanchain_034/scan_select_in vccd1 vssd1 scanchain
Xscanchain_044 scanchain_044/clk_in scanchain_045/clk_in scanchain_044/data_in scanchain_045/data_in
+ scanchain_044/latch_enable_in scanchain_045/latch_enable_in gbsha_ttfir_top_044/io_in[0]
+ gbsha_ttfir_top_044/io_in[1] gbsha_ttfir_top_044/io_in[2] gbsha_ttfir_top_044/io_in[3]
+ gbsha_ttfir_top_044/io_in[4] gbsha_ttfir_top_044/io_in[5] gbsha_ttfir_top_044/io_in[6]
+ gbsha_ttfir_top_044/io_in[7] gbsha_ttfir_top_044/io_out[0] gbsha_ttfir_top_044/io_out[1]
+ gbsha_ttfir_top_044/io_out[2] gbsha_ttfir_top_044/io_out[3] gbsha_ttfir_top_044/io_out[4]
+ gbsha_ttfir_top_044/io_out[5] gbsha_ttfir_top_044/io_out[6] gbsha_ttfir_top_044/io_out[7]
+ scanchain_044/scan_select_in scanchain_045/scan_select_in vccd1 vssd1 scanchain
Xscanchain_055 scanchain_055/clk_in scanchain_056/clk_in scanchain_055/data_in scanchain_056/data_in
+ scanchain_055/latch_enable_in scanchain_056/latch_enable_in scanchain_055/module_data_in[0]
+ scanchain_055/module_data_in[1] scanchain_055/module_data_in[2] scanchain_055/module_data_in[3]
+ scanchain_055/module_data_in[4] scanchain_055/module_data_in[5] scanchain_055/module_data_in[6]
+ scanchain_055/module_data_in[7] scanchain_055/module_data_out[0] scanchain_055/module_data_out[1]
+ scanchain_055/module_data_out[2] scanchain_055/module_data_out[3] scanchain_055/module_data_out[4]
+ scanchain_055/module_data_out[5] scanchain_055/module_data_out[6] scanchain_055/module_data_out[7]
+ scanchain_055/scan_select_in scanchain_056/scan_select_in vccd1 vssd1 scanchain
Xuser_module_361728533238569985_193 scanchain_193/module_data_in[0] scanchain_193/module_data_in[1]
+ scanchain_193/module_data_in[2] scanchain_193/module_data_in[3] scanchain_193/module_data_in[4]
+ scanchain_193/module_data_in[5] scanchain_193/module_data_in[6] scanchain_193/module_data_in[7]
+ scanchain_193/module_data_out[0] scanchain_193/module_data_out[1] scanchain_193/module_data_out[2]
+ scanchain_193/module_data_out[3] scanchain_193/module_data_out[4] scanchain_193/module_data_out[5]
+ scanchain_193/module_data_out[6] scanchain_193/module_data_out[7] vccd1 vssd1 user_module_361728533238569985
Xuser_module_361728533238569985_182 scanchain_182/module_data_in[0] scanchain_182/module_data_in[1]
+ scanchain_182/module_data_in[2] scanchain_182/module_data_in[3] scanchain_182/module_data_in[4]
+ scanchain_182/module_data_in[5] scanchain_182/module_data_in[6] scanchain_182/module_data_in[7]
+ scanchain_182/module_data_out[0] scanchain_182/module_data_out[1] scanchain_182/module_data_out[2]
+ scanchain_182/module_data_out[3] scanchain_182/module_data_out[4] scanchain_182/module_data_out[5]
+ scanchain_182/module_data_out[6] scanchain_182/module_data_out[7] vccd1 vssd1 user_module_361728533238569985
Xscanchain_066 scanchain_066/clk_in scanchain_067/clk_in scanchain_066/data_in scanchain_067/data_in
+ scanchain_066/latch_enable_in scanchain_067/latch_enable_in zl_uart_066/io_in[0]
+ zl_uart_066/io_in[1] zl_uart_066/io_in[2] zl_uart_066/io_in[3] zl_uart_066/io_in[4]
+ zl_uart_066/io_in[5] zl_uart_066/io_in[6] zl_uart_066/io_in[7] zl_uart_066/io_out[0]
+ zl_uart_066/io_out[1] zl_uart_066/io_out[2] zl_uart_066/io_out[3] zl_uart_066/io_out[4]
+ zl_uart_066/io_out[5] zl_uart_066/io_out[6] zl_uart_066/io_out[7] scanchain_066/scan_select_in
+ scanchain_067/scan_select_in vccd1 vssd1 scanchain
Xuser_module_361728533238569985_171 scanchain_171/module_data_in[0] scanchain_171/module_data_in[1]
+ scanchain_171/module_data_in[2] scanchain_171/module_data_in[3] scanchain_171/module_data_in[4]
+ scanchain_171/module_data_in[5] scanchain_171/module_data_in[6] scanchain_171/module_data_in[7]
+ scanchain_171/module_data_out[0] scanchain_171/module_data_out[1] scanchain_171/module_data_out[2]
+ scanchain_171/module_data_out[3] scanchain_171/module_data_out[4] scanchain_171/module_data_out[5]
+ scanchain_171/module_data_out[6] scanchain_171/module_data_out[7] vccd1 vssd1 user_module_361728533238569985
Xscanchain_077 scanchain_077/clk_in scanchain_078/clk_in scanchain_077/data_in scanchain_078/data_in
+ scanchain_077/latch_enable_in scanchain_078/latch_enable_in scanchain_077/module_data_in[0]
+ scanchain_077/module_data_in[1] scanchain_077/module_data_in[2] scanchain_077/module_data_in[3]
+ scanchain_077/module_data_in[4] scanchain_077/module_data_in[5] scanchain_077/module_data_in[6]
+ scanchain_077/module_data_in[7] scanchain_077/module_data_out[0] scanchain_077/module_data_out[1]
+ scanchain_077/module_data_out[2] scanchain_077/module_data_out[3] scanchain_077/module_data_out[4]
+ scanchain_077/module_data_out[5] scanchain_077/module_data_out[6] scanchain_077/module_data_out[7]
+ scanchain_077/scan_select_in scanchain_078/scan_select_in vccd1 vssd1 scanchain
Xscanchain_088 scanchain_088/clk_in scanchain_089/clk_in scanchain_088/data_in scanchain_089/data_in
+ scanchain_088/latch_enable_in scanchain_089/latch_enable_in scanchain_088/module_data_in[0]
+ scanchain_088/module_data_in[1] scanchain_088/module_data_in[2] scanchain_088/module_data_in[3]
+ scanchain_088/module_data_in[4] scanchain_088/module_data_in[5] scanchain_088/module_data_in[6]
+ scanchain_088/module_data_in[7] scanchain_088/module_data_out[0] scanchain_088/module_data_out[1]
+ scanchain_088/module_data_out[2] scanchain_088/module_data_out[3] scanchain_088/module_data_out[4]
+ scanchain_088/module_data_out[5] scanchain_088/module_data_out[6] scanchain_088/module_data_out[7]
+ scanchain_088/scan_select_in scanchain_089/scan_select_in vccd1 vssd1 scanchain
Xuser_module_361728533238569985_160 scanchain_160/module_data_in[0] scanchain_160/module_data_in[1]
+ scanchain_160/module_data_in[2] scanchain_160/module_data_in[3] scanchain_160/module_data_in[4]
+ scanchain_160/module_data_in[5] scanchain_160/module_data_in[6] scanchain_160/module_data_in[7]
+ scanchain_160/module_data_out[0] scanchain_160/module_data_out[1] scanchain_160/module_data_out[2]
+ scanchain_160/module_data_out[3] scanchain_160/module_data_out[4] scanchain_160/module_data_out[5]
+ scanchain_160/module_data_out[6] scanchain_160/module_data_out[7] vccd1 vssd1 user_module_361728533238569985
Xuser_module_357752736742764545_002 scanchain_002/module_data_in[0] scanchain_002/module_data_in[1]
+ scanchain_002/module_data_in[2] scanchain_002/module_data_in[3] scanchain_002/module_data_in[4]
+ scanchain_002/module_data_in[5] scanchain_002/module_data_in[6] scanchain_002/module_data_in[7]
+ scanchain_002/module_data_out[0] scanchain_002/module_data_out[1] scanchain_002/module_data_out[2]
+ scanchain_002/module_data_out[3] scanchain_002/module_data_out[4] scanchain_002/module_data_out[5]
+ scanchain_002/module_data_out[6] scanchain_002/module_data_out[7] vccd1 vssd1 user_module_357752736742764545
Xscanchain_226 scanchain_226/clk_in scanchain_227/clk_in scanchain_226/data_in scanchain_227/data_in
+ scanchain_226/latch_enable_in scanchain_227/latch_enable_in scanchain_226/module_data_in[0]
+ scanchain_226/module_data_in[1] scanchain_226/module_data_in[2] scanchain_226/module_data_in[3]
+ scanchain_226/module_data_in[4] scanchain_226/module_data_in[5] scanchain_226/module_data_in[6]
+ scanchain_226/module_data_in[7] scanchain_226/module_data_out[0] scanchain_226/module_data_out[1]
+ scanchain_226/module_data_out[2] scanchain_226/module_data_out[3] scanchain_226/module_data_out[4]
+ scanchain_226/module_data_out[5] scanchain_226/module_data_out[6] scanchain_226/module_data_out[7]
+ scanchain_226/scan_select_in scanchain_227/scan_select_in vccd1 vssd1 scanchain
Xscanchain_237 scanchain_237/clk_in scanchain_238/clk_in scanchain_237/data_in scanchain_238/data_in
+ scanchain_237/latch_enable_in scanchain_238/latch_enable_in scanchain_237/module_data_in[0]
+ scanchain_237/module_data_in[1] scanchain_237/module_data_in[2] scanchain_237/module_data_in[3]
+ scanchain_237/module_data_in[4] scanchain_237/module_data_in[5] scanchain_237/module_data_in[6]
+ scanchain_237/module_data_in[7] scanchain_237/module_data_out[0] scanchain_237/module_data_out[1]
+ scanchain_237/module_data_out[2] scanchain_237/module_data_out[3] scanchain_237/module_data_out[4]
+ scanchain_237/module_data_out[5] scanchain_237/module_data_out[6] scanchain_237/module_data_out[7]
+ scanchain_237/scan_select_in scanchain_238/scan_select_in vccd1 vssd1 scanchain
Xscanchain_248 scanchain_248/clk_in scanchain_249/clk_in scanchain_248/data_in scanchain_249/data_in
+ scanchain_248/latch_enable_in scanchain_249/latch_enable_in scanchain_248/module_data_in[0]
+ scanchain_248/module_data_in[1] scanchain_248/module_data_in[2] scanchain_248/module_data_in[3]
+ scanchain_248/module_data_in[4] scanchain_248/module_data_in[5] scanchain_248/module_data_in[6]
+ scanchain_248/module_data_in[7] scanchain_248/module_data_out[0] scanchain_248/module_data_out[1]
+ scanchain_248/module_data_out[2] scanchain_248/module_data_out[3] scanchain_248/module_data_out[4]
+ scanchain_248/module_data_out[5] scanchain_248/module_data_out[6] scanchain_248/module_data_out[7]
+ scanchain_248/scan_select_in scanchain_249/scan_select_in vccd1 vssd1 scanchain
Xscanchain_215 scanchain_215/clk_in scanchain_216/clk_in scanchain_215/data_in scanchain_216/data_in
+ scanchain_215/latch_enable_in scanchain_216/latch_enable_in scanchain_215/module_data_in[0]
+ scanchain_215/module_data_in[1] scanchain_215/module_data_in[2] scanchain_215/module_data_in[3]
+ scanchain_215/module_data_in[4] scanchain_215/module_data_in[5] scanchain_215/module_data_in[6]
+ scanchain_215/module_data_in[7] scanchain_215/module_data_out[0] scanchain_215/module_data_out[1]
+ scanchain_215/module_data_out[2] scanchain_215/module_data_out[3] scanchain_215/module_data_out[4]
+ scanchain_215/module_data_out[5] scanchain_215/module_data_out[6] scanchain_215/module_data_out[7]
+ scanchain_215/scan_select_in scanchain_216/scan_select_in vccd1 vssd1 scanchain
Xscanchain_204 scanchain_204/clk_in scanchain_205/clk_in scanchain_204/data_in scanchain_205/data_in
+ scanchain_204/latch_enable_in scanchain_205/latch_enable_in scanchain_204/module_data_in[0]
+ scanchain_204/module_data_in[1] scanchain_204/module_data_in[2] scanchain_204/module_data_in[3]
+ scanchain_204/module_data_in[4] scanchain_204/module_data_in[5] scanchain_204/module_data_in[6]
+ scanchain_204/module_data_in[7] scanchain_204/module_data_out[0] scanchain_204/module_data_out[1]
+ scanchain_204/module_data_out[2] scanchain_204/module_data_out[3] scanchain_204/module_data_out[4]
+ scanchain_204/module_data_out[5] scanchain_204/module_data_out[6] scanchain_204/module_data_out[7]
+ scanchain_204/scan_select_in scanchain_205/scan_select_in vccd1 vssd1 scanchain
Xuser_module_362208154278843393_075 scanchain_075/module_data_in[0] scanchain_075/module_data_in[1]
+ scanchain_075/module_data_in[2] scanchain_075/module_data_in[3] scanchain_075/module_data_in[4]
+ scanchain_075/module_data_in[5] scanchain_075/module_data_in[6] scanchain_075/module_data_in[7]
+ scanchain_075/module_data_out[0] scanchain_075/module_data_out[1] scanchain_075/module_data_out[2]
+ scanchain_075/module_data_out[3] scanchain_075/module_data_out[4] scanchain_075/module_data_out[5]
+ scanchain_075/module_data_out[6] scanchain_075/module_data_out[7] vccd1 vssd1 user_module_362208154278843393
Xuser_module_361728533238569985_150 scanchain_150/module_data_in[0] scanchain_150/module_data_in[1]
+ scanchain_150/module_data_in[2] scanchain_150/module_data_in[3] scanchain_150/module_data_in[4]
+ scanchain_150/module_data_in[5] scanchain_150/module_data_in[6] scanchain_150/module_data_in[7]
+ scanchain_150/module_data_out[0] scanchain_150/module_data_out[1] scanchain_150/module_data_out[2]
+ scanchain_150/module_data_out[3] scanchain_150/module_data_out[4] scanchain_150/module_data_out[5]
+ scanchain_150/module_data_out[6] scanchain_150/module_data_out[7] vccd1 vssd1 user_module_361728533238569985
Xscanchain_012 scanchain_012/clk_in scanchain_013/clk_in scanchain_012/data_in scanchain_013/data_in
+ scanchain_012/latch_enable_in scanchain_013/latch_enable_in scanchain_012/module_data_in[0]
+ scanchain_012/module_data_in[1] scanchain_012/module_data_in[2] scanchain_012/module_data_in[3]
+ scanchain_012/module_data_in[4] scanchain_012/module_data_in[5] scanchain_012/module_data_in[6]
+ scanchain_012/module_data_in[7] scanchain_012/module_data_out[0] scanchain_012/module_data_out[1]
+ scanchain_012/module_data_out[2] scanchain_012/module_data_out[3] scanchain_012/module_data_out[4]
+ scanchain_012/module_data_out[5] scanchain_012/module_data_out[6] scanchain_012/module_data_out[7]
+ scanchain_012/scan_select_in scanchain_013/scan_select_in vccd1 vssd1 scanchain
Xscanchain_001 scanchain_001/clk_in scanchain_002/clk_in scanchain_001/data_in scanchain_002/data_in
+ scanchain_001/latch_enable_in scanchain_002/latch_enable_in morningjava_top_001/io_in[0]
+ morningjava_top_001/io_in[1] morningjava_top_001/io_in[2] morningjava_top_001/io_in[3]
+ morningjava_top_001/io_in[4] morningjava_top_001/io_in[5] morningjava_top_001/io_in[6]
+ morningjava_top_001/io_in[7] morningjava_top_001/io_out[0] morningjava_top_001/io_out[1]
+ morningjava_top_001/io_out[2] morningjava_top_001/io_out[3] morningjava_top_001/io_out[4]
+ morningjava_top_001/io_out[5] morningjava_top_001/io_out[6] morningjava_top_001/io_out[7]
+ scanchain_001/scan_select_in scanchain_002/scan_select_in vccd1 vssd1 scanchain
Xscanchain_023 scanchain_023/clk_in scanchain_024/clk_in scanchain_023/data_in scanchain_024/data_in
+ scanchain_023/latch_enable_in scanchain_024/latch_enable_in diferential_rvb2_023/io_in[0]
+ diferential_rvb2_023/io_in[1] diferential_rvb2_023/io_in[2] diferential_rvb2_023/io_in[3]
+ diferential_rvb2_023/io_in[4] diferential_rvb2_023/io_in[5] diferential_rvb2_023/io_in[6]
+ diferential_rvb2_023/io_in[7] diferential_rvb2_023/io_out[0] diferential_rvb2_023/io_out[1]
+ diferential_rvb2_023/io_out[2] diferential_rvb2_023/io_out[3] diferential_rvb2_023/io_out[4]
+ diferential_rvb2_023/io_out[5] diferential_rvb2_023/io_out[6] diferential_rvb2_023/io_out[7]
+ scanchain_023/scan_select_in scanchain_024/scan_select_in vccd1 vssd1 scanchain
Xscanchain_034 scanchain_034/clk_in scanchain_035/clk_in scanchain_034/data_in scanchain_035/data_in
+ scanchain_034/latch_enable_in scanchain_035/latch_enable_in scanchain_034/module_data_in[0]
+ scanchain_034/module_data_in[1] scanchain_034/module_data_in[2] scanchain_034/module_data_in[3]
+ scanchain_034/module_data_in[4] scanchain_034/module_data_in[5] scanchain_034/module_data_in[6]
+ scanchain_034/module_data_in[7] scanchain_034/module_data_out[0] scanchain_034/module_data_out[1]
+ scanchain_034/module_data_out[2] scanchain_034/module_data_out[3] scanchain_034/module_data_out[4]
+ scanchain_034/module_data_out[5] scanchain_034/module_data_out[6] scanchain_034/module_data_out[7]
+ scanchain_034/scan_select_in scanchain_035/scan_select_in vccd1 vssd1 scanchain
Xscanchain_045 scanchain_045/clk_in scanchain_046/clk_in scanchain_045/data_in scanchain_046/data_in
+ scanchain_045/latch_enable_in scanchain_046/latch_enable_in kiwih_tt_top_045/io_in[0]
+ kiwih_tt_top_045/io_in[1] kiwih_tt_top_045/io_in[2] kiwih_tt_top_045/io_in[3] kiwih_tt_top_045/io_in[4]
+ kiwih_tt_top_045/io_in[5] kiwih_tt_top_045/io_in[6] kiwih_tt_top_045/io_in[7] kiwih_tt_top_045/io_out[0]
+ kiwih_tt_top_045/io_out[1] kiwih_tt_top_045/io_out[2] kiwih_tt_top_045/io_out[3]
+ kiwih_tt_top_045/io_out[4] kiwih_tt_top_045/io_out[5] kiwih_tt_top_045/io_out[6]
+ kiwih_tt_top_045/io_out[7] scanchain_045/scan_select_in scanchain_046/scan_select_in
+ vccd1 vssd1 scanchain
Xuser_module_361728533238569985_194 scanchain_194/module_data_in[0] scanchain_194/module_data_in[1]
+ scanchain_194/module_data_in[2] scanchain_194/module_data_in[3] scanchain_194/module_data_in[4]
+ scanchain_194/module_data_in[5] scanchain_194/module_data_in[6] scanchain_194/module_data_in[7]
+ scanchain_194/module_data_out[0] scanchain_194/module_data_out[1] scanchain_194/module_data_out[2]
+ scanchain_194/module_data_out[3] scanchain_194/module_data_out[4] scanchain_194/module_data_out[5]
+ scanchain_194/module_data_out[6] scanchain_194/module_data_out[7] vccd1 vssd1 user_module_361728533238569985
Xscanchain_056 scanchain_056/clk_in scanchain_057/clk_in scanchain_056/data_in scanchain_057/data_in
+ scanchain_056/latch_enable_in scanchain_057/latch_enable_in scanchain_056/module_data_in[0]
+ scanchain_056/module_data_in[1] scanchain_056/module_data_in[2] scanchain_056/module_data_in[3]
+ scanchain_056/module_data_in[4] scanchain_056/module_data_in[5] scanchain_056/module_data_in[6]
+ scanchain_056/module_data_in[7] scanchain_056/module_data_out[0] scanchain_056/module_data_out[1]
+ scanchain_056/module_data_out[2] scanchain_056/module_data_out[3] scanchain_056/module_data_out[4]
+ scanchain_056/module_data_out[5] scanchain_056/module_data_out[6] scanchain_056/module_data_out[7]
+ scanchain_056/scan_select_in scanchain_057/scan_select_in vccd1 vssd1 scanchain
Xuser_module_361728533238569985_183 scanchain_183/module_data_in[0] scanchain_183/module_data_in[1]
+ scanchain_183/module_data_in[2] scanchain_183/module_data_in[3] scanchain_183/module_data_in[4]
+ scanchain_183/module_data_in[5] scanchain_183/module_data_in[6] scanchain_183/module_data_in[7]
+ scanchain_183/module_data_out[0] scanchain_183/module_data_out[1] scanchain_183/module_data_out[2]
+ scanchain_183/module_data_out[3] scanchain_183/module_data_out[4] scanchain_183/module_data_out[5]
+ scanchain_183/module_data_out[6] scanchain_183/module_data_out[7] vccd1 vssd1 user_module_361728533238569985
Xscanchain_067 scanchain_067/clk_in scanchain_068/clk_in scanchain_067/data_in scanchain_068/data_in
+ scanchain_067/latch_enable_in scanchain_068/latch_enable_in jmw95_top_067/io_in[0]
+ jmw95_top_067/io_in[1] jmw95_top_067/io_in[2] jmw95_top_067/io_in[3] jmw95_top_067/io_in[4]
+ jmw95_top_067/io_in[5] jmw95_top_067/io_in[6] jmw95_top_067/io_in[7] jmw95_top_067/io_out[0]
+ jmw95_top_067/io_out[1] jmw95_top_067/io_out[2] jmw95_top_067/io_out[3] jmw95_top_067/io_out[4]
+ jmw95_top_067/io_out[5] jmw95_top_067/io_out[6] jmw95_top_067/io_out[7] scanchain_067/scan_select_in
+ scanchain_068/scan_select_in vccd1 vssd1 scanchain
Xscanchain_078 scanchain_078/clk_in scanchain_079/clk_in scanchain_078/data_in scanchain_079/data_in
+ scanchain_078/latch_enable_in scanchain_079/latch_enable_in scanchain_078/module_data_in[0]
+ scanchain_078/module_data_in[1] scanchain_078/module_data_in[2] scanchain_078/module_data_in[3]
+ scanchain_078/module_data_in[4] scanchain_078/module_data_in[5] scanchain_078/module_data_in[6]
+ scanchain_078/module_data_in[7] scanchain_078/module_data_out[0] scanchain_078/module_data_out[1]
+ scanchain_078/module_data_out[2] scanchain_078/module_data_out[3] scanchain_078/module_data_out[4]
+ scanchain_078/module_data_out[5] scanchain_078/module_data_out[6] scanchain_078/module_data_out[7]
+ scanchain_078/scan_select_in scanchain_079/scan_select_in vccd1 vssd1 scanchain
Xuser_module_361728533238569985_172 scanchain_172/module_data_in[0] scanchain_172/module_data_in[1]
+ scanchain_172/module_data_in[2] scanchain_172/module_data_in[3] scanchain_172/module_data_in[4]
+ scanchain_172/module_data_in[5] scanchain_172/module_data_in[6] scanchain_172/module_data_in[7]
+ scanchain_172/module_data_out[0] scanchain_172/module_data_out[1] scanchain_172/module_data_out[2]
+ scanchain_172/module_data_out[3] scanchain_172/module_data_out[4] scanchain_172/module_data_out[5]
+ scanchain_172/module_data_out[6] scanchain_172/module_data_out[7] vccd1 vssd1 user_module_361728533238569985
Xuser_module_361728533238569985_161 scanchain_161/module_data_in[0] scanchain_161/module_data_in[1]
+ scanchain_161/module_data_in[2] scanchain_161/module_data_in[3] scanchain_161/module_data_in[4]
+ scanchain_161/module_data_in[5] scanchain_161/module_data_in[6] scanchain_161/module_data_in[7]
+ scanchain_161/module_data_out[0] scanchain_161/module_data_out[1] scanchain_161/module_data_out[2]
+ scanchain_161/module_data_out[3] scanchain_161/module_data_out[4] scanchain_161/module_data_out[5]
+ scanchain_161/module_data_out[6] scanchain_161/module_data_out[7] vccd1 vssd1 user_module_361728533238569985
Xscanchain_089 scanchain_089/clk_in scanchain_090/clk_in scanchain_089/data_in scanchain_090/data_in
+ scanchain_089/latch_enable_in scanchain_090/latch_enable_in scanchain_089/module_data_in[0]
+ scanchain_089/module_data_in[1] scanchain_089/module_data_in[2] scanchain_089/module_data_in[3]
+ scanchain_089/module_data_in[4] scanchain_089/module_data_in[5] scanchain_089/module_data_in[6]
+ scanchain_089/module_data_in[7] scanchain_089/module_data_out[0] scanchain_089/module_data_out[1]
+ scanchain_089/module_data_out[2] scanchain_089/module_data_out[3] scanchain_089/module_data_out[4]
+ scanchain_089/module_data_out[5] scanchain_089/module_data_out[6] scanchain_089/module_data_out[7]
+ scanchain_089/scan_select_in scanchain_090/scan_select_in vccd1 vssd1 scanchain
Xscanchain_238 scanchain_238/clk_in scanchain_239/clk_in scanchain_238/data_in scanchain_239/data_in
+ scanchain_238/latch_enable_in scanchain_239/latch_enable_in scanchain_238/module_data_in[0]
+ scanchain_238/module_data_in[1] scanchain_238/module_data_in[2] scanchain_238/module_data_in[3]
+ scanchain_238/module_data_in[4] scanchain_238/module_data_in[5] scanchain_238/module_data_in[6]
+ scanchain_238/module_data_in[7] scanchain_238/module_data_out[0] scanchain_238/module_data_out[1]
+ scanchain_238/module_data_out[2] scanchain_238/module_data_out[3] scanchain_238/module_data_out[4]
+ scanchain_238/module_data_out[5] scanchain_238/module_data_out[6] scanchain_238/module_data_out[7]
+ scanchain_238/scan_select_in scanchain_239/scan_select_in vccd1 vssd1 scanchain
Xscanchain_249 scanchain_249/clk_in scanchain_249/clk_out scanchain_249/data_in scanchain_249/data_out
+ scanchain_249/latch_enable_in scanchain_249/latch_enable_out scanchain_249/module_data_in[0]
+ scanchain_249/module_data_in[1] scanchain_249/module_data_in[2] scanchain_249/module_data_in[3]
+ scanchain_249/module_data_in[4] scanchain_249/module_data_in[5] scanchain_249/module_data_in[6]
+ scanchain_249/module_data_in[7] scanchain_249/module_data_out[0] scanchain_249/module_data_out[1]
+ scanchain_249/module_data_out[2] scanchain_249/module_data_out[3] scanchain_249/module_data_out[4]
+ scanchain_249/module_data_out[5] scanchain_249/module_data_out[6] scanchain_249/module_data_out[7]
+ scanchain_249/scan_select_in scanchain_249/scan_select_out vccd1 vssd1 scanchain
Xscanchain_227 scanchain_227/clk_in scanchain_228/clk_in scanchain_227/data_in scanchain_228/data_in
+ scanchain_227/latch_enable_in scanchain_228/latch_enable_in scanchain_227/module_data_in[0]
+ scanchain_227/module_data_in[1] scanchain_227/module_data_in[2] scanchain_227/module_data_in[3]
+ scanchain_227/module_data_in[4] scanchain_227/module_data_in[5] scanchain_227/module_data_in[6]
+ scanchain_227/module_data_in[7] scanchain_227/module_data_out[0] scanchain_227/module_data_out[1]
+ scanchain_227/module_data_out[2] scanchain_227/module_data_out[3] scanchain_227/module_data_out[4]
+ scanchain_227/module_data_out[5] scanchain_227/module_data_out[6] scanchain_227/module_data_out[7]
+ scanchain_227/scan_select_in scanchain_228/scan_select_in vccd1 vssd1 scanchain
Xscanchain_216 scanchain_216/clk_in scanchain_217/clk_in scanchain_216/data_in scanchain_217/data_in
+ scanchain_216/latch_enable_in scanchain_217/latch_enable_in scanchain_216/module_data_in[0]
+ scanchain_216/module_data_in[1] scanchain_216/module_data_in[2] scanchain_216/module_data_in[3]
+ scanchain_216/module_data_in[4] scanchain_216/module_data_in[5] scanchain_216/module_data_in[6]
+ scanchain_216/module_data_in[7] scanchain_216/module_data_out[0] scanchain_216/module_data_out[1]
+ scanchain_216/module_data_out[2] scanchain_216/module_data_out[3] scanchain_216/module_data_out[4]
+ scanchain_216/module_data_out[5] scanchain_216/module_data_out[6] scanchain_216/module_data_out[7]
+ scanchain_216/scan_select_in scanchain_217/scan_select_in vccd1 vssd1 scanchain
Xscanchain_205 scanchain_205/clk_in scanchain_206/clk_in scanchain_205/data_in scanchain_206/data_in
+ scanchain_205/latch_enable_in scanchain_206/latch_enable_in scanchain_205/module_data_in[0]
+ scanchain_205/module_data_in[1] scanchain_205/module_data_in[2] scanchain_205/module_data_in[3]
+ scanchain_205/module_data_in[4] scanchain_205/module_data_in[5] scanchain_205/module_data_in[6]
+ scanchain_205/module_data_in[7] scanchain_205/module_data_out[0] scanchain_205/module_data_out[1]
+ scanchain_205/module_data_out[2] scanchain_205/module_data_out[3] scanchain_205/module_data_out[4]
+ scanchain_205/module_data_out[5] scanchain_205/module_data_out[6] scanchain_205/module_data_out[7]
+ scanchain_205/scan_select_in scanchain_206/scan_select_in vccd1 vssd1 scanchain
Xuser_module_361728533238569985_140 scanchain_140/module_data_in[0] scanchain_140/module_data_in[1]
+ scanchain_140/module_data_in[2] scanchain_140/module_data_in[3] scanchain_140/module_data_in[4]
+ scanchain_140/module_data_in[5] scanchain_140/module_data_in[6] scanchain_140/module_data_in[7]
+ scanchain_140/module_data_out[0] scanchain_140/module_data_out[1] scanchain_140/module_data_out[2]
+ scanchain_140/module_data_out[3] scanchain_140/module_data_out[4] scanchain_140/module_data_out[5]
+ scanchain_140/module_data_out[6] scanchain_140/module_data_out[7] vccd1 vssd1 user_module_361728533238569985
Xuser_module_361728533238569985_151 scanchain_151/module_data_in[0] scanchain_151/module_data_in[1]
+ scanchain_151/module_data_in[2] scanchain_151/module_data_in[3] scanchain_151/module_data_in[4]
+ scanchain_151/module_data_in[5] scanchain_151/module_data_in[6] scanchain_151/module_data_in[7]
+ scanchain_151/module_data_out[0] scanchain_151/module_data_out[1] scanchain_151/module_data_out[2]
+ scanchain_151/module_data_out[3] scanchain_151/module_data_out[4] scanchain_151/module_data_out[5]
+ scanchain_151/module_data_out[6] scanchain_151/module_data_out[7] vccd1 vssd1 user_module_361728533238569985
Xscanchain_024 scanchain_024/clk_in scanchain_025/clk_in scanchain_024/data_in scanchain_025/data_in
+ scanchain_024/latch_enable_in scanchain_025/latch_enable_in diferential_rvb3_024/io_in[0]
+ diferential_rvb3_024/io_in[1] diferential_rvb3_024/io_in[2] diferential_rvb3_024/io_in[3]
+ diferential_rvb3_024/io_in[4] diferential_rvb3_024/io_in[5] diferential_rvb3_024/io_in[6]
+ diferential_rvb3_024/io_in[7] diferential_rvb3_024/io_out[0] diferential_rvb3_024/io_out[1]
+ diferential_rvb3_024/io_out[2] diferential_rvb3_024/io_out[3] diferential_rvb3_024/io_out[4]
+ diferential_rvb3_024/io_out[5] diferential_rvb3_024/io_out[6] diferential_rvb3_024/io_out[7]
+ scanchain_024/scan_select_in scanchain_025/scan_select_in vccd1 vssd1 scanchain
Xscanchain_013 scanchain_013/clk_in scanchain_014/clk_in scanchain_013/data_in scanchain_014/data_in
+ scanchain_013/latch_enable_in scanchain_014/latch_enable_in greenstyle_lfsr_013/io_in[0]
+ greenstyle_lfsr_013/io_in[1] greenstyle_lfsr_013/io_in[2] greenstyle_lfsr_013/io_in[3]
+ greenstyle_lfsr_013/io_in[4] greenstyle_lfsr_013/io_in[5] greenstyle_lfsr_013/io_in[6]
+ greenstyle_lfsr_013/io_in[7] greenstyle_lfsr_013/io_out[0] greenstyle_lfsr_013/io_out[1]
+ greenstyle_lfsr_013/io_out[2] greenstyle_lfsr_013/io_out[3] greenstyle_lfsr_013/io_out[4]
+ greenstyle_lfsr_013/io_out[5] greenstyle_lfsr_013/io_out[6] greenstyle_lfsr_013/io_out[7]
+ scanchain_013/scan_select_in scanchain_014/scan_select_in vccd1 vssd1 scanchain
Xscanchain_002 scanchain_002/clk_in scanchain_003/clk_in scanchain_002/data_in scanchain_003/data_in
+ scanchain_002/latch_enable_in scanchain_003/latch_enable_in scanchain_002/module_data_in[0]
+ scanchain_002/module_data_in[1] scanchain_002/module_data_in[2] scanchain_002/module_data_in[3]
+ scanchain_002/module_data_in[4] scanchain_002/module_data_in[5] scanchain_002/module_data_in[6]
+ scanchain_002/module_data_in[7] scanchain_002/module_data_out[0] scanchain_002/module_data_out[1]
+ scanchain_002/module_data_out[2] scanchain_002/module_data_out[3] scanchain_002/module_data_out[4]
+ scanchain_002/module_data_out[5] scanchain_002/module_data_out[6] scanchain_002/module_data_out[7]
+ scanchain_002/scan_select_in scanchain_003/scan_select_in vccd1 vssd1 scanchain
Xscanchain_035 scanchain_035/clk_in scanchain_036/clk_in scanchain_035/data_in scanchain_036/data_in
+ scanchain_035/latch_enable_in scanchain_036/latch_enable_in nikor_clock_035/io_in[0]
+ nikor_clock_035/io_in[1] nikor_clock_035/io_in[2] nikor_clock_035/io_in[3] nikor_clock_035/io_in[4]
+ nikor_clock_035/io_in[5] nikor_clock_035/io_in[6] nikor_clock_035/io_in[7] nikor_clock_035/io_out[0]
+ nikor_clock_035/io_out[1] nikor_clock_035/io_out[2] nikor_clock_035/io_out[3] nikor_clock_035/io_out[4]
+ nikor_clock_035/io_out[5] nikor_clock_035/io_out[6] nikor_clock_035/io_out[7] scanchain_035/scan_select_in
+ scanchain_036/scan_select_in vccd1 vssd1 scanchain
Xscanchain_046 scanchain_046/clk_in scanchain_047/clk_in scanchain_046/data_in scanchain_047/data_in
+ scanchain_046/latch_enable_in scanchain_047/latch_enable_in scanchain_046/module_data_in[0]
+ scanchain_046/module_data_in[1] scanchain_046/module_data_in[2] scanchain_046/module_data_in[3]
+ scanchain_046/module_data_in[4] scanchain_046/module_data_in[5] scanchain_046/module_data_in[6]
+ scanchain_046/module_data_in[7] scanchain_046/module_data_out[0] scanchain_046/module_data_out[1]
+ scanchain_046/module_data_out[2] scanchain_046/module_data_out[3] scanchain_046/module_data_out[4]
+ scanchain_046/module_data_out[5] scanchain_046/module_data_out[6] scanchain_046/module_data_out[7]
+ scanchain_046/scan_select_in scanchain_047/scan_select_in vccd1 vssd1 scanchain
Xuser_module_361728533238569985_195 scanchain_195/module_data_in[0] scanchain_195/module_data_in[1]
+ scanchain_195/module_data_in[2] scanchain_195/module_data_in[3] scanchain_195/module_data_in[4]
+ scanchain_195/module_data_in[5] scanchain_195/module_data_in[6] scanchain_195/module_data_in[7]
+ scanchain_195/module_data_out[0] scanchain_195/module_data_out[1] scanchain_195/module_data_out[2]
+ scanchain_195/module_data_out[3] scanchain_195/module_data_out[4] scanchain_195/module_data_out[5]
+ scanchain_195/module_data_out[6] scanchain_195/module_data_out[7] vccd1 vssd1 user_module_361728533238569985
Xscanchain_057 scanchain_057/clk_in scanchain_058/clk_in scanchain_057/data_in scanchain_058/data_in
+ scanchain_057/latch_enable_in scanchain_058/latch_enable_in scanchain_057/module_data_in[0]
+ scanchain_057/module_data_in[1] scanchain_057/module_data_in[2] scanchain_057/module_data_in[3]
+ scanchain_057/module_data_in[4] scanchain_057/module_data_in[5] scanchain_057/module_data_in[6]
+ scanchain_057/module_data_in[7] scanchain_057/module_data_out[0] scanchain_057/module_data_out[1]
+ scanchain_057/module_data_out[2] scanchain_057/module_data_out[3] scanchain_057/module_data_out[4]
+ scanchain_057/module_data_out[5] scanchain_057/module_data_out[6] scanchain_057/module_data_out[7]
+ scanchain_057/scan_select_in scanchain_058/scan_select_in vccd1 vssd1 scanchain
Xuser_module_361728533238569985_184 scanchain_184/module_data_in[0] scanchain_184/module_data_in[1]
+ scanchain_184/module_data_in[2] scanchain_184/module_data_in[3] scanchain_184/module_data_in[4]
+ scanchain_184/module_data_in[5] scanchain_184/module_data_in[6] scanchain_184/module_data_in[7]
+ scanchain_184/module_data_out[0] scanchain_184/module_data_out[1] scanchain_184/module_data_out[2]
+ scanchain_184/module_data_out[3] scanchain_184/module_data_out[4] scanchain_184/module_data_out[5]
+ scanchain_184/module_data_out[6] scanchain_184/module_data_out[7] vccd1 vssd1 user_module_361728533238569985
Xuser_module_361728533238569985_173 scanchain_173/module_data_in[0] scanchain_173/module_data_in[1]
+ scanchain_173/module_data_in[2] scanchain_173/module_data_in[3] scanchain_173/module_data_in[4]
+ scanchain_173/module_data_in[5] scanchain_173/module_data_in[6] scanchain_173/module_data_in[7]
+ scanchain_173/module_data_out[0] scanchain_173/module_data_out[1] scanchain_173/module_data_out[2]
+ scanchain_173/module_data_out[3] scanchain_173/module_data_out[4] scanchain_173/module_data_out[5]
+ scanchain_173/module_data_out[6] scanchain_173/module_data_out[7] vccd1 vssd1 user_module_361728533238569985
Xuser_module_361728533238569985_162 scanchain_162/module_data_in[0] scanchain_162/module_data_in[1]
+ scanchain_162/module_data_in[2] scanchain_162/module_data_in[3] scanchain_162/module_data_in[4]
+ scanchain_162/module_data_in[5] scanchain_162/module_data_in[6] scanchain_162/module_data_in[7]
+ scanchain_162/module_data_out[0] scanchain_162/module_data_out[1] scanchain_162/module_data_out[2]
+ scanchain_162/module_data_out[3] scanchain_162/module_data_out[4] scanchain_162/module_data_out[5]
+ scanchain_162/module_data_out[6] scanchain_162/module_data_out[7] vccd1 vssd1 user_module_361728533238569985
Xuser_module_359357227471086593_011 scanchain_011/module_data_in[0] scanchain_011/module_data_in[1]
+ scanchain_011/module_data_in[2] scanchain_011/module_data_in[3] scanchain_011/module_data_in[4]
+ scanchain_011/module_data_in[5] scanchain_011/module_data_in[6] scanchain_011/module_data_in[7]
+ scanchain_011/module_data_out[0] scanchain_011/module_data_out[1] scanchain_011/module_data_out[2]
+ scanchain_011/module_data_out[3] scanchain_011/module_data_out[4] scanchain_011/module_data_out[5]
+ scanchain_011/module_data_out[6] scanchain_011/module_data_out[7] vccd1 vssd1 user_module_359357227471086593
Xscanchain_068 scanchain_068/clk_in scanchain_069/clk_in scanchain_068/data_in scanchain_069/data_in
+ scanchain_068/latch_enable_in scanchain_069/latch_enable_in scanchain_068/module_data_in[0]
+ scanchain_068/module_data_in[1] scanchain_068/module_data_in[2] scanchain_068/module_data_in[3]
+ scanchain_068/module_data_in[4] scanchain_068/module_data_in[5] scanchain_068/module_data_in[6]
+ scanchain_068/module_data_in[7] scanchain_068/module_data_out[0] scanchain_068/module_data_out[1]
+ scanchain_068/module_data_out[2] scanchain_068/module_data_out[3] scanchain_068/module_data_out[4]
+ scanchain_068/module_data_out[5] scanchain_068/module_data_out[6] scanchain_068/module_data_out[7]
+ scanchain_068/scan_select_in scanchain_069/scan_select_in vccd1 vssd1 scanchain
Xscanchain_079 scanchain_079/clk_in scanchain_080/clk_in scanchain_079/data_in scanchain_080/data_in
+ scanchain_079/latch_enable_in scanchain_080/latch_enable_in scanchain_079/module_data_in[0]
+ scanchain_079/module_data_in[1] scanchain_079/module_data_in[2] scanchain_079/module_data_in[3]
+ scanchain_079/module_data_in[4] scanchain_079/module_data_in[5] scanchain_079/module_data_in[6]
+ scanchain_079/module_data_in[7] scanchain_079/module_data_out[0] scanchain_079/module_data_out[1]
+ scanchain_079/module_data_out[2] scanchain_079/module_data_out[3] scanchain_079/module_data_out[4]
+ scanchain_079/module_data_out[5] scanchain_079/module_data_out[6] scanchain_079/module_data_out[7]
+ scanchain_079/scan_select_in scanchain_080/scan_select_in vccd1 vssd1 scanchain
Xscanchain_239 scanchain_239/clk_in scanchain_240/clk_in scanchain_239/data_in scanchain_240/data_in
+ scanchain_239/latch_enable_in scanchain_240/latch_enable_in scanchain_239/module_data_in[0]
+ scanchain_239/module_data_in[1] scanchain_239/module_data_in[2] scanchain_239/module_data_in[3]
+ scanchain_239/module_data_in[4] scanchain_239/module_data_in[5] scanchain_239/module_data_in[6]
+ scanchain_239/module_data_in[7] scanchain_239/module_data_out[0] scanchain_239/module_data_out[1]
+ scanchain_239/module_data_out[2] scanchain_239/module_data_out[3] scanchain_239/module_data_out[4]
+ scanchain_239/module_data_out[5] scanchain_239/module_data_out[6] scanchain_239/module_data_out[7]
+ scanchain_239/scan_select_in scanchain_240/scan_select_in vccd1 vssd1 scanchain
Xscanchain_228 scanchain_228/clk_in scanchain_229/clk_in scanchain_228/data_in scanchain_229/data_in
+ scanchain_228/latch_enable_in scanchain_229/latch_enable_in scanchain_228/module_data_in[0]
+ scanchain_228/module_data_in[1] scanchain_228/module_data_in[2] scanchain_228/module_data_in[3]
+ scanchain_228/module_data_in[4] scanchain_228/module_data_in[5] scanchain_228/module_data_in[6]
+ scanchain_228/module_data_in[7] scanchain_228/module_data_out[0] scanchain_228/module_data_out[1]
+ scanchain_228/module_data_out[2] scanchain_228/module_data_out[3] scanchain_228/module_data_out[4]
+ scanchain_228/module_data_out[5] scanchain_228/module_data_out[6] scanchain_228/module_data_out[7]
+ scanchain_228/scan_select_in scanchain_229/scan_select_in vccd1 vssd1 scanchain
Xscanchain_217 scanchain_217/clk_in scanchain_218/clk_in scanchain_217/data_in scanchain_218/data_in
+ scanchain_217/latch_enable_in scanchain_218/latch_enable_in scanchain_217/module_data_in[0]
+ scanchain_217/module_data_in[1] scanchain_217/module_data_in[2] scanchain_217/module_data_in[3]
+ scanchain_217/module_data_in[4] scanchain_217/module_data_in[5] scanchain_217/module_data_in[6]
+ scanchain_217/module_data_in[7] scanchain_217/module_data_out[0] scanchain_217/module_data_out[1]
+ scanchain_217/module_data_out[2] scanchain_217/module_data_out[3] scanchain_217/module_data_out[4]
+ scanchain_217/module_data_out[5] scanchain_217/module_data_out[6] scanchain_217/module_data_out[7]
+ scanchain_217/scan_select_in scanchain_218/scan_select_in vccd1 vssd1 scanchain
Xscanchain_206 scanchain_206/clk_in scanchain_207/clk_in scanchain_206/data_in scanchain_207/data_in
+ scanchain_206/latch_enable_in scanchain_207/latch_enable_in scanchain_206/module_data_in[0]
+ scanchain_206/module_data_in[1] scanchain_206/module_data_in[2] scanchain_206/module_data_in[3]
+ scanchain_206/module_data_in[4] scanchain_206/module_data_in[5] scanchain_206/module_data_in[6]
+ scanchain_206/module_data_in[7] scanchain_206/module_data_out[0] scanchain_206/module_data_out[1]
+ scanchain_206/module_data_out[2] scanchain_206/module_data_out[3] scanchain_206/module_data_out[4]
+ scanchain_206/module_data_out[5] scanchain_206/module_data_out[6] scanchain_206/module_data_out[7]
+ scanchain_206/scan_select_in scanchain_207/scan_select_in vccd1 vssd1 scanchain
Xuser_module_361728533238569985_130 scanchain_130/module_data_in[0] scanchain_130/module_data_in[1]
+ scanchain_130/module_data_in[2] scanchain_130/module_data_in[3] scanchain_130/module_data_in[4]
+ scanchain_130/module_data_in[5] scanchain_130/module_data_in[6] scanchain_130/module_data_in[7]
+ scanchain_130/module_data_out[0] scanchain_130/module_data_out[1] scanchain_130/module_data_out[2]
+ scanchain_130/module_data_out[3] scanchain_130/module_data_out[4] scanchain_130/module_data_out[5]
+ scanchain_130/module_data_out[6] scanchain_130/module_data_out[7] vccd1 vssd1 user_module_361728533238569985
Xuser_module_361728533238569985_141 scanchain_141/module_data_in[0] scanchain_141/module_data_in[1]
+ scanchain_141/module_data_in[2] scanchain_141/module_data_in[3] scanchain_141/module_data_in[4]
+ scanchain_141/module_data_in[5] scanchain_141/module_data_in[6] scanchain_141/module_data_in[7]
+ scanchain_141/module_data_out[0] scanchain_141/module_data_out[1] scanchain_141/module_data_out[2]
+ scanchain_141/module_data_out[3] scanchain_141/module_data_out[4] scanchain_141/module_data_out[5]
+ scanchain_141/module_data_out[6] scanchain_141/module_data_out[7] vccd1 vssd1 user_module_361728533238569985
Xuser_module_361728533238569985_152 scanchain_152/module_data_in[0] scanchain_152/module_data_in[1]
+ scanchain_152/module_data_in[2] scanchain_152/module_data_in[3] scanchain_152/module_data_in[4]
+ scanchain_152/module_data_in[5] scanchain_152/module_data_in[6] scanchain_152/module_data_in[7]
+ scanchain_152/module_data_out[0] scanchain_152/module_data_out[1] scanchain_152/module_data_out[2]
+ scanchain_152/module_data_out[3] scanchain_152/module_data_out[4] scanchain_152/module_data_out[5]
+ scanchain_152/module_data_out[6] scanchain_152/module_data_out[7] vccd1 vssd1 user_module_361728533238569985
Xuser_module_361728533238569985_163 scanchain_163/module_data_in[0] scanchain_163/module_data_in[1]
+ scanchain_163/module_data_in[2] scanchain_163/module_data_in[3] scanchain_163/module_data_in[4]
+ scanchain_163/module_data_in[5] scanchain_163/module_data_in[6] scanchain_163/module_data_in[7]
+ scanchain_163/module_data_out[0] scanchain_163/module_data_out[1] scanchain_163/module_data_out[2]
+ scanchain_163/module_data_out[3] scanchain_163/module_data_out[4] scanchain_163/module_data_out[5]
+ scanchain_163/module_data_out[6] scanchain_163/module_data_out[7] vccd1 vssd1 user_module_361728533238569985
Xscanchain_025 scanchain_025/clk_in scanchain_026/clk_in scanchain_025/data_in scanchain_026/data_in
+ scanchain_025/latch_enable_in scanchain_026/latch_enable_in diferential_rvb4_025/io_in[0]
+ diferential_rvb4_025/io_in[1] diferential_rvb4_025/io_in[2] diferential_rvb4_025/io_in[3]
+ diferential_rvb4_025/io_in[4] diferential_rvb4_025/io_in[5] diferential_rvb4_025/io_in[6]
+ diferential_rvb4_025/io_in[7] diferential_rvb4_025/io_out[0] diferential_rvb4_025/io_out[1]
+ diferential_rvb4_025/io_out[2] diferential_rvb4_025/io_out[3] diferential_rvb4_025/io_out[4]
+ diferential_rvb4_025/io_out[5] diferential_rvb4_025/io_out[6] diferential_rvb4_025/io_out[7]
+ scanchain_025/scan_select_in scanchain_026/scan_select_in vccd1 vssd1 scanchain
Xscanchain_014 scanchain_014/clk_in scanchain_015/clk_in scanchain_014/data_in scanchain_015/data_in
+ scanchain_014/latch_enable_in scanchain_015/latch_enable_in scanchain_014/module_data_in[0]
+ scanchain_014/module_data_in[1] scanchain_014/module_data_in[2] scanchain_014/module_data_in[3]
+ scanchain_014/module_data_in[4] scanchain_014/module_data_in[5] scanchain_014/module_data_in[6]
+ scanchain_014/module_data_in[7] scanchain_014/module_data_out[0] scanchain_014/module_data_out[1]
+ scanchain_014/module_data_out[2] scanchain_014/module_data_out[3] scanchain_014/module_data_out[4]
+ scanchain_014/module_data_out[5] scanchain_014/module_data_out[6] scanchain_014/module_data_out[7]
+ scanchain_014/scan_select_in scanchain_015/scan_select_in vccd1 vssd1 scanchain
Xscanchain_003 scanchain_003/clk_in scanchain_004/clk_in scanchain_003/data_in scanchain_004/data_in
+ scanchain_003/latch_enable_in scanchain_004/latch_enable_in meiniki_pi_003/io_in[0]
+ meiniki_pi_003/io_in[1] meiniki_pi_003/io_in[2] meiniki_pi_003/io_in[3] meiniki_pi_003/io_in[4]
+ meiniki_pi_003/io_in[5] meiniki_pi_003/io_in[6] meiniki_pi_003/io_in[7] meiniki_pi_003/io_out[0]
+ meiniki_pi_003/io_out[1] meiniki_pi_003/io_out[2] meiniki_pi_003/io_out[3] meiniki_pi_003/io_out[4]
+ meiniki_pi_003/io_out[5] meiniki_pi_003/io_out[6] meiniki_pi_003/io_out[7] scanchain_003/scan_select_in
+ scanchain_004/scan_select_in vccd1 vssd1 scanchain
Xscanchain_036 scanchain_036/clk_in scanchain_037/clk_in scanchain_036/data_in scanchain_037/data_in
+ scanchain_036/latch_enable_in scanchain_037/latch_enable_in scanchain_036/module_data_in[0]
+ scanchain_036/module_data_in[1] scanchain_036/module_data_in[2] scanchain_036/module_data_in[3]
+ scanchain_036/module_data_in[4] scanchain_036/module_data_in[5] scanchain_036/module_data_in[6]
+ scanchain_036/module_data_in[7] scanchain_036/module_data_out[0] scanchain_036/module_data_out[1]
+ scanchain_036/module_data_out[2] scanchain_036/module_data_out[3] scanchain_036/module_data_out[4]
+ scanchain_036/module_data_out[5] scanchain_036/module_data_out[6] scanchain_036/module_data_out[7]
+ scanchain_036/scan_select_in scanchain_037/scan_select_in vccd1 vssd1 scanchain
Xscanchain_047 scanchain_047/clk_in scanchain_048/clk_in scanchain_047/data_in scanchain_048/data_in
+ scanchain_047/latch_enable_in scanchain_048/latch_enable_in my_design_047/io_in[0]
+ my_design_047/io_in[1] my_design_047/io_in[2] my_design_047/io_in[3] my_design_047/io_in[4]
+ my_design_047/io_in[5] my_design_047/io_in[6] my_design_047/io_in[7] my_design_047/io_out[0]
+ my_design_047/io_out[1] my_design_047/io_out[2] my_design_047/io_out[3] my_design_047/io_out[4]
+ my_design_047/io_out[5] my_design_047/io_out[6] my_design_047/io_out[7] scanchain_047/scan_select_in
+ scanchain_048/scan_select_in vccd1 vssd1 scanchain
Xuser_module_361728533238569985_196 scanchain_196/module_data_in[0] scanchain_196/module_data_in[1]
+ scanchain_196/module_data_in[2] scanchain_196/module_data_in[3] scanchain_196/module_data_in[4]
+ scanchain_196/module_data_in[5] scanchain_196/module_data_in[6] scanchain_196/module_data_in[7]
+ scanchain_196/module_data_out[0] scanchain_196/module_data_out[1] scanchain_196/module_data_out[2]
+ scanchain_196/module_data_out[3] scanchain_196/module_data_out[4] scanchain_196/module_data_out[5]
+ scanchain_196/module_data_out[6] scanchain_196/module_data_out[7] vccd1 vssd1 user_module_361728533238569985
Xscanchain_058 scanchain_058/clk_in scanchain_059/clk_in scanchain_058/data_in scanchain_059/data_in
+ scanchain_058/latch_enable_in scanchain_059/latch_enable_in BenAtUvu_combo_058/io_in[0]
+ BenAtUvu_combo_058/io_in[1] BenAtUvu_combo_058/io_in[2] BenAtUvu_combo_058/io_in[3]
+ BenAtUvu_combo_058/io_in[4] BenAtUvu_combo_058/io_in[5] BenAtUvu_combo_058/io_in[6]
+ BenAtUvu_combo_058/io_in[7] BenAtUvu_combo_058/io_out[0] BenAtUvu_combo_058/io_out[1]
+ BenAtUvu_combo_058/io_out[2] BenAtUvu_combo_058/io_out[3] BenAtUvu_combo_058/io_out[4]
+ BenAtUvu_combo_058/io_out[5] BenAtUvu_combo_058/io_out[6] BenAtUvu_combo_058/io_out[7]
+ scanchain_058/scan_select_in scanchain_059/scan_select_in vccd1 vssd1 scanchain
Xuser_module_361728533238569985_185 scanchain_185/module_data_in[0] scanchain_185/module_data_in[1]
+ scanchain_185/module_data_in[2] scanchain_185/module_data_in[3] scanchain_185/module_data_in[4]
+ scanchain_185/module_data_in[5] scanchain_185/module_data_in[6] scanchain_185/module_data_in[7]
+ scanchain_185/module_data_out[0] scanchain_185/module_data_out[1] scanchain_185/module_data_out[2]
+ scanchain_185/module_data_out[3] scanchain_185/module_data_out[4] scanchain_185/module_data_out[5]
+ scanchain_185/module_data_out[6] scanchain_185/module_data_out[7] vccd1 vssd1 user_module_361728533238569985
Xscanchain_069 scanchain_069/clk_in scanchain_070/clk_in scanchain_069/data_in scanchain_070/data_in
+ scanchain_069/latch_enable_in scanchain_070/latch_enable_in scanchain_069/module_data_in[0]
+ scanchain_069/module_data_in[1] scanchain_069/module_data_in[2] scanchain_069/module_data_in[3]
+ scanchain_069/module_data_in[4] scanchain_069/module_data_in[5] scanchain_069/module_data_in[6]
+ scanchain_069/module_data_in[7] scanchain_069/module_data_out[0] scanchain_069/module_data_out[1]
+ scanchain_069/module_data_out[2] scanchain_069/module_data_out[3] scanchain_069/module_data_out[4]
+ scanchain_069/module_data_out[5] scanchain_069/module_data_out[6] scanchain_069/module_data_out[7]
+ scanchain_069/scan_select_in scanchain_070/scan_select_in vccd1 vssd1 scanchain
Xuser_module_361728533238569985_174 scanchain_174/module_data_in[0] scanchain_174/module_data_in[1]
+ scanchain_174/module_data_in[2] scanchain_174/module_data_in[3] scanchain_174/module_data_in[4]
+ scanchain_174/module_data_in[5] scanchain_174/module_data_in[6] scanchain_174/module_data_in[7]
+ scanchain_174/module_data_out[0] scanchain_174/module_data_out[1] scanchain_174/module_data_out[2]
+ scanchain_174/module_data_out[3] scanchain_174/module_data_out[4] scanchain_174/module_data_out[5]
+ scanchain_174/module_data_out[6] scanchain_174/module_data_out[7] vccd1 vssd1 user_module_361728533238569985
Xuser_module_362592986761938945_076 scanchain_076/module_data_in[0] scanchain_076/module_data_in[1]
+ scanchain_076/module_data_in[2] scanchain_076/module_data_in[3] scanchain_076/module_data_in[4]
+ scanchain_076/module_data_in[5] scanchain_076/module_data_in[6] scanchain_076/module_data_in[7]
+ scanchain_076/module_data_out[0] scanchain_076/module_data_out[1] scanchain_076/module_data_out[2]
+ scanchain_076/module_data_out[3] scanchain_076/module_data_out[4] scanchain_076/module_data_out[5]
+ scanchain_076/module_data_out[6] scanchain_076/module_data_out[7] vccd1 vssd1 user_module_362592986761938945
Xscanchain_229 scanchain_229/clk_in scanchain_230/clk_in scanchain_229/data_in scanchain_230/data_in
+ scanchain_229/latch_enable_in scanchain_230/latch_enable_in scanchain_229/module_data_in[0]
+ scanchain_229/module_data_in[1] scanchain_229/module_data_in[2] scanchain_229/module_data_in[3]
+ scanchain_229/module_data_in[4] scanchain_229/module_data_in[5] scanchain_229/module_data_in[6]
+ scanchain_229/module_data_in[7] scanchain_229/module_data_out[0] scanchain_229/module_data_out[1]
+ scanchain_229/module_data_out[2] scanchain_229/module_data_out[3] scanchain_229/module_data_out[4]
+ scanchain_229/module_data_out[5] scanchain_229/module_data_out[6] scanchain_229/module_data_out[7]
+ scanchain_229/scan_select_in scanchain_230/scan_select_in vccd1 vssd1 scanchain
Xscanchain_218 scanchain_218/clk_in scanchain_219/clk_in scanchain_218/data_in scanchain_219/data_in
+ scanchain_218/latch_enable_in scanchain_219/latch_enable_in scanchain_218/module_data_in[0]
+ scanchain_218/module_data_in[1] scanchain_218/module_data_in[2] scanchain_218/module_data_in[3]
+ scanchain_218/module_data_in[4] scanchain_218/module_data_in[5] scanchain_218/module_data_in[6]
+ scanchain_218/module_data_in[7] scanchain_218/module_data_out[0] scanchain_218/module_data_out[1]
+ scanchain_218/module_data_out[2] scanchain_218/module_data_out[3] scanchain_218/module_data_out[4]
+ scanchain_218/module_data_out[5] scanchain_218/module_data_out[6] scanchain_218/module_data_out[7]
+ scanchain_218/scan_select_in scanchain_219/scan_select_in vccd1 vssd1 scanchain
Xscanchain_207 scanchain_207/clk_in scanchain_208/clk_in scanchain_207/data_in scanchain_208/data_in
+ scanchain_207/latch_enable_in scanchain_208/latch_enable_in scanchain_207/module_data_in[0]
+ scanchain_207/module_data_in[1] scanchain_207/module_data_in[2] scanchain_207/module_data_in[3]
+ scanchain_207/module_data_in[4] scanchain_207/module_data_in[5] scanchain_207/module_data_in[6]
+ scanchain_207/module_data_in[7] scanchain_207/module_data_out[0] scanchain_207/module_data_out[1]
+ scanchain_207/module_data_out[2] scanchain_207/module_data_out[3] scanchain_207/module_data_out[4]
+ scanchain_207/module_data_out[5] scanchain_207/module_data_out[6] scanchain_207/module_data_out[7]
+ scanchain_207/scan_select_in scanchain_208/scan_select_in vccd1 vssd1 scanchain
Xuser_module_361728533238569985_131 scanchain_131/module_data_in[0] scanchain_131/module_data_in[1]
+ scanchain_131/module_data_in[2] scanchain_131/module_data_in[3] scanchain_131/module_data_in[4]
+ scanchain_131/module_data_in[5] scanchain_131/module_data_in[6] scanchain_131/module_data_in[7]
+ scanchain_131/module_data_out[0] scanchain_131/module_data_out[1] scanchain_131/module_data_out[2]
+ scanchain_131/module_data_out[3] scanchain_131/module_data_out[4] scanchain_131/module_data_out[5]
+ scanchain_131/module_data_out[6] scanchain_131/module_data_out[7] vccd1 vssd1 user_module_361728533238569985
Xuser_module_361728533238569985_120 scanchain_120/module_data_in[0] scanchain_120/module_data_in[1]
+ scanchain_120/module_data_in[2] scanchain_120/module_data_in[3] scanchain_120/module_data_in[4]
+ scanchain_120/module_data_in[5] scanchain_120/module_data_in[6] scanchain_120/module_data_in[7]
+ scanchain_120/module_data_out[0] scanchain_120/module_data_out[1] scanchain_120/module_data_out[2]
+ scanchain_120/module_data_out[3] scanchain_120/module_data_out[4] scanchain_120/module_data_out[5]
+ scanchain_120/module_data_out[6] scanchain_120/module_data_out[7] vccd1 vssd1 user_module_361728533238569985
Xuser_module_361728533238569985_142 scanchain_142/module_data_in[0] scanchain_142/module_data_in[1]
+ scanchain_142/module_data_in[2] scanchain_142/module_data_in[3] scanchain_142/module_data_in[4]
+ scanchain_142/module_data_in[5] scanchain_142/module_data_in[6] scanchain_142/module_data_in[7]
+ scanchain_142/module_data_out[0] scanchain_142/module_data_out[1] scanchain_142/module_data_out[2]
+ scanchain_142/module_data_out[3] scanchain_142/module_data_out[4] scanchain_142/module_data_out[5]
+ scanchain_142/module_data_out[6] scanchain_142/module_data_out[7] vccd1 vssd1 user_module_361728533238569985
Xscanchain_026 scanchain_026/clk_in scanchain_027/clk_in scanchain_026/data_in scanchain_027/data_in
+ scanchain_026/latch_enable_in scanchain_027/latch_enable_in scanchain_026/module_data_in[0]
+ scanchain_026/module_data_in[1] scanchain_026/module_data_in[2] scanchain_026/module_data_in[3]
+ scanchain_026/module_data_in[4] scanchain_026/module_data_in[5] scanchain_026/module_data_in[6]
+ scanchain_026/module_data_in[7] scanchain_026/module_data_out[0] scanchain_026/module_data_out[1]
+ scanchain_026/module_data_out[2] scanchain_026/module_data_out[3] scanchain_026/module_data_out[4]
+ scanchain_026/module_data_out[5] scanchain_026/module_data_out[6] scanchain_026/module_data_out[7]
+ scanchain_026/scan_select_in scanchain_027/scan_select_in vccd1 vssd1 scanchain
Xscanchain_015 scanchain_015/clk_in scanchain_016/clk_in scanchain_015/data_in scanchain_016/data_in
+ scanchain_015/latch_enable_in scanchain_016/latch_enable_in scanchain_015/module_data_in[0]
+ scanchain_015/module_data_in[1] scanchain_015/module_data_in[2] scanchain_015/module_data_in[3]
+ scanchain_015/module_data_in[4] scanchain_015/module_data_in[5] scanchain_015/module_data_in[6]
+ scanchain_015/module_data_in[7] scanchain_015/module_data_out[0] scanchain_015/module_data_out[1]
+ scanchain_015/module_data_out[2] scanchain_015/module_data_out[3] scanchain_015/module_data_out[4]
+ scanchain_015/module_data_out[5] scanchain_015/module_data_out[6] scanchain_015/module_data_out[7]
+ scanchain_015/scan_select_in scanchain_016/scan_select_in vccd1 vssd1 scanchain
Xscanchain_004 scanchain_004/clk_in scanchain_005/clk_in scanchain_004/data_in scanchain_005/data_in
+ scanchain_004/latch_enable_in scanchain_005/latch_enable_in wormy_top_004/io_in[0]
+ wormy_top_004/io_in[1] wormy_top_004/io_in[2] wormy_top_004/io_in[3] wormy_top_004/io_in[4]
+ wormy_top_004/io_in[5] wormy_top_004/io_in[6] wormy_top_004/io_in[7] wormy_top_004/io_out[0]
+ wormy_top_004/io_out[1] wormy_top_004/io_out[2] wormy_top_004/io_out[3] wormy_top_004/io_out[4]
+ wormy_top_004/io_out[5] wormy_top_004/io_out[6] wormy_top_004/io_out[7] scanchain_004/scan_select_in
+ scanchain_005/scan_select_in vccd1 vssd1 scanchain
Xscanchain_037 scanchain_037/clk_in scanchain_038/clk_in scanchain_037/data_in scanchain_038/data_in
+ scanchain_037/latch_enable_in scanchain_038/latch_enable_in scanchain_037/module_data_in[0]
+ scanchain_037/module_data_in[1] scanchain_037/module_data_in[2] scanchain_037/module_data_in[3]
+ scanchain_037/module_data_in[4] scanchain_037/module_data_in[5] scanchain_037/module_data_in[6]
+ scanchain_037/module_data_in[7] scanchain_037/module_data_out[0] scanchain_037/module_data_out[1]
+ scanchain_037/module_data_out[2] scanchain_037/module_data_out[3] scanchain_037/module_data_out[4]
+ scanchain_037/module_data_out[5] scanchain_037/module_data_out[6] scanchain_037/module_data_out[7]
+ scanchain_037/scan_select_in scanchain_038/scan_select_in vccd1 vssd1 scanchain
Xuser_module_361728533238569985_197 scanchain_197/module_data_in[0] scanchain_197/module_data_in[1]
+ scanchain_197/module_data_in[2] scanchain_197/module_data_in[3] scanchain_197/module_data_in[4]
+ scanchain_197/module_data_in[5] scanchain_197/module_data_in[6] scanchain_197/module_data_in[7]
+ scanchain_197/module_data_out[0] scanchain_197/module_data_out[1] scanchain_197/module_data_out[2]
+ scanchain_197/module_data_out[3] scanchain_197/module_data_out[4] scanchain_197/module_data_out[5]
+ scanchain_197/module_data_out[6] scanchain_197/module_data_out[7] vccd1 vssd1 user_module_361728533238569985
Xscanchain_048 scanchain_048/clk_in scanchain_049/clk_in scanchain_048/data_in scanchain_049/data_in
+ scanchain_048/latch_enable_in scanchain_049/latch_enable_in scanchain_048/module_data_in[0]
+ scanchain_048/module_data_in[1] scanchain_048/module_data_in[2] scanchain_048/module_data_in[3]
+ scanchain_048/module_data_in[4] scanchain_048/module_data_in[5] scanchain_048/module_data_in[6]
+ scanchain_048/module_data_in[7] scanchain_048/module_data_out[0] scanchain_048/module_data_out[1]
+ scanchain_048/module_data_out[2] scanchain_048/module_data_out[3] scanchain_048/module_data_out[4]
+ scanchain_048/module_data_out[5] scanchain_048/module_data_out[6] scanchain_048/module_data_out[7]
+ scanchain_048/scan_select_in scanchain_049/scan_select_in vccd1 vssd1 scanchain
Xscanchain_059 scanchain_059/clk_in scanchain_060/clk_in scanchain_059/data_in scanchain_060/data_in
+ scanchain_059/latch_enable_in scanchain_060/latch_enable_in top_tt03_059/io_in[0]
+ top_tt03_059/io_in[1] top_tt03_059/io_in[2] top_tt03_059/io_in[3] top_tt03_059/io_in[4]
+ top_tt03_059/io_in[5] top_tt03_059/io_in[6] top_tt03_059/io_in[7] top_tt03_059/io_out[0]
+ top_tt03_059/io_out[1] top_tt03_059/io_out[2] top_tt03_059/io_out[3] top_tt03_059/io_out[4]
+ top_tt03_059/io_out[5] top_tt03_059/io_out[6] top_tt03_059/io_out[7] scanchain_059/scan_select_in
+ scanchain_060/scan_select_in vccd1 vssd1 scanchain
Xuser_module_361728533238569985_186 scanchain_186/module_data_in[0] scanchain_186/module_data_in[1]
+ scanchain_186/module_data_in[2] scanchain_186/module_data_in[3] scanchain_186/module_data_in[4]
+ scanchain_186/module_data_in[5] scanchain_186/module_data_in[6] scanchain_186/module_data_in[7]
+ scanchain_186/module_data_out[0] scanchain_186/module_data_out[1] scanchain_186/module_data_out[2]
+ scanchain_186/module_data_out[3] scanchain_186/module_data_out[4] scanchain_186/module_data_out[5]
+ scanchain_186/module_data_out[6] scanchain_186/module_data_out[7] vccd1 vssd1 user_module_361728533238569985
Xuser_module_361728533238569985_175 scanchain_175/module_data_in[0] scanchain_175/module_data_in[1]
+ scanchain_175/module_data_in[2] scanchain_175/module_data_in[3] scanchain_175/module_data_in[4]
+ scanchain_175/module_data_in[5] scanchain_175/module_data_in[6] scanchain_175/module_data_in[7]
+ scanchain_175/module_data_out[0] scanchain_175/module_data_out[1] scanchain_175/module_data_out[2]
+ scanchain_175/module_data_out[3] scanchain_175/module_data_out[4] scanchain_175/module_data_out[5]
+ scanchain_175/module_data_out[6] scanchain_175/module_data_out[7] vccd1 vssd1 user_module_361728533238569985
Xuser_module_361728533238569985_164 scanchain_164/module_data_in[0] scanchain_164/module_data_in[1]
+ scanchain_164/module_data_in[2] scanchain_164/module_data_in[3] scanchain_164/module_data_in[4]
+ scanchain_164/module_data_in[5] scanchain_164/module_data_in[6] scanchain_164/module_data_in[7]
+ scanchain_164/module_data_out[0] scanchain_164/module_data_out[1] scanchain_164/module_data_out[2]
+ scanchain_164/module_data_out[3] scanchain_164/module_data_out[4] scanchain_164/module_data_out[5]
+ scanchain_164/module_data_out[6] scanchain_164/module_data_out[7] vccd1 vssd1 user_module_361728533238569985
Xuser_module_361728533238569985_153 scanchain_153/module_data_in[0] scanchain_153/module_data_in[1]
+ scanchain_153/module_data_in[2] scanchain_153/module_data_in[3] scanchain_153/module_data_in[4]
+ scanchain_153/module_data_in[5] scanchain_153/module_data_in[6] scanchain_153/module_data_in[7]
+ scanchain_153/module_data_out[0] scanchain_153/module_data_out[1] scanchain_153/module_data_out[2]
+ scanchain_153/module_data_out[3] scanchain_153/module_data_out[4] scanchain_153/module_data_out[5]
+ scanchain_153/module_data_out[6] scanchain_153/module_data_out[7] vccd1 vssd1 user_module_361728533238569985
Xdiferential_rvb4_025 diferential_rvb4_025/io_in[0] diferential_rvb4_025/io_in[1]
+ diferential_rvb4_025/io_in[2] diferential_rvb4_025/io_in[3] diferential_rvb4_025/io_in[4]
+ diferential_rvb4_025/io_in[5] diferential_rvb4_025/io_in[6] diferential_rvb4_025/io_in[7]
+ diferential_rvb4_025/io_out[0] diferential_rvb4_025/io_out[1] diferential_rvb4_025/io_out[2]
+ diferential_rvb4_025/io_out[3] diferential_rvb4_025/io_out[4] diferential_rvb4_025/io_out[5]
+ diferential_rvb4_025/io_out[6] diferential_rvb4_025/io_out[7] vccd1 vssd1 diferential_rvb4
Xscanchain_219 scanchain_219/clk_in scanchain_220/clk_in scanchain_219/data_in scanchain_220/data_in
+ scanchain_219/latch_enable_in scanchain_220/latch_enable_in scanchain_219/module_data_in[0]
+ scanchain_219/module_data_in[1] scanchain_219/module_data_in[2] scanchain_219/module_data_in[3]
+ scanchain_219/module_data_in[4] scanchain_219/module_data_in[5] scanchain_219/module_data_in[6]
+ scanchain_219/module_data_in[7] scanchain_219/module_data_out[0] scanchain_219/module_data_out[1]
+ scanchain_219/module_data_out[2] scanchain_219/module_data_out[3] scanchain_219/module_data_out[4]
+ scanchain_219/module_data_out[5] scanchain_219/module_data_out[6] scanchain_219/module_data_out[7]
+ scanchain_219/scan_select_in scanchain_220/scan_select_in vccd1 vssd1 scanchain
Xscanchain_208 scanchain_208/clk_in scanchain_209/clk_in scanchain_208/data_in scanchain_209/data_in
+ scanchain_208/latch_enable_in scanchain_209/latch_enable_in scanchain_208/module_data_in[0]
+ scanchain_208/module_data_in[1] scanchain_208/module_data_in[2] scanchain_208/module_data_in[3]
+ scanchain_208/module_data_in[4] scanchain_208/module_data_in[5] scanchain_208/module_data_in[6]
+ scanchain_208/module_data_in[7] scanchain_208/module_data_out[0] scanchain_208/module_data_out[1]
+ scanchain_208/module_data_out[2] scanchain_208/module_data_out[3] scanchain_208/module_data_out[4]
+ scanchain_208/module_data_out[5] scanchain_208/module_data_out[6] scanchain_208/module_data_out[7]
+ scanchain_208/scan_select_in scanchain_209/scan_select_in vccd1 vssd1 scanchain
Xtiny_bnn_072 tiny_bnn_072/io_in[0] tiny_bnn_072/io_in[1] tiny_bnn_072/io_in[2] tiny_bnn_072/io_in[3]
+ tiny_bnn_072/io_in[4] tiny_bnn_072/io_in[5] tiny_bnn_072/io_in[6] tiny_bnn_072/io_in[7]
+ tiny_bnn_072/io_out[0] tiny_bnn_072/io_out[1] tiny_bnn_072/io_out[2] tiny_bnn_072/io_out[3]
+ tiny_bnn_072/io_out[4] tiny_bnn_072/io_out[5] tiny_bnn_072/io_out[6] tiny_bnn_072/io_out[7]
+ vccd1 vssd1 tiny_bnn
Xuser_module_361728533238569985_121 scanchain_121/module_data_in[0] scanchain_121/module_data_in[1]
+ scanchain_121/module_data_in[2] scanchain_121/module_data_in[3] scanchain_121/module_data_in[4]
+ scanchain_121/module_data_in[5] scanchain_121/module_data_in[6] scanchain_121/module_data_in[7]
+ scanchain_121/module_data_out[0] scanchain_121/module_data_out[1] scanchain_121/module_data_out[2]
+ scanchain_121/module_data_out[3] scanchain_121/module_data_out[4] scanchain_121/module_data_out[5]
+ scanchain_121/module_data_out[6] scanchain_121/module_data_out[7] vccd1 vssd1 user_module_361728533238569985
Xuser_module_361728533238569985_132 scanchain_132/module_data_in[0] scanchain_132/module_data_in[1]
+ scanchain_132/module_data_in[2] scanchain_132/module_data_in[3] scanchain_132/module_data_in[4]
+ scanchain_132/module_data_in[5] scanchain_132/module_data_in[6] scanchain_132/module_data_in[7]
+ scanchain_132/module_data_out[0] scanchain_132/module_data_out[1] scanchain_132/module_data_out[2]
+ scanchain_132/module_data_out[3] scanchain_132/module_data_out[4] scanchain_132/module_data_out[5]
+ scanchain_132/module_data_out[6] scanchain_132/module_data_out[7] vccd1 vssd1 user_module_361728533238569985
Xuser_module_361728533238569985_143 scanchain_143/module_data_in[0] scanchain_143/module_data_in[1]
+ scanchain_143/module_data_in[2] scanchain_143/module_data_in[3] scanchain_143/module_data_in[4]
+ scanchain_143/module_data_in[5] scanchain_143/module_data_in[6] scanchain_143/module_data_in[7]
+ scanchain_143/module_data_out[0] scanchain_143/module_data_out[1] scanchain_143/module_data_out[2]
+ scanchain_143/module_data_out[3] scanchain_143/module_data_out[4] scanchain_143/module_data_out[5]
+ scanchain_143/module_data_out[6] scanchain_143/module_data_out[7] vccd1 vssd1 user_module_361728533238569985
Xuser_module_361728533238569985_110 scanchain_110/module_data_in[0] scanchain_110/module_data_in[1]
+ scanchain_110/module_data_in[2] scanchain_110/module_data_in[3] scanchain_110/module_data_in[4]
+ scanchain_110/module_data_in[5] scanchain_110/module_data_in[6] scanchain_110/module_data_in[7]
+ scanchain_110/module_data_out[0] scanchain_110/module_data_out[1] scanchain_110/module_data_out[2]
+ scanchain_110/module_data_out[3] scanchain_110/module_data_out[4] scanchain_110/module_data_out[5]
+ scanchain_110/module_data_out[6] scanchain_110/module_data_out[7] vccd1 vssd1 user_module_361728533238569985
Xscanchain_016 scanchain_016/clk_in scanchain_017/clk_in scanchain_016/data_in scanchain_017/data_in
+ scanchain_016/latch_enable_in scanchain_017/latch_enable_in shadow1229_player_016/io_in[0]
+ shadow1229_player_016/io_in[1] shadow1229_player_016/io_in[2] shadow1229_player_016/io_in[3]
+ shadow1229_player_016/io_in[4] shadow1229_player_016/io_in[5] shadow1229_player_016/io_in[6]
+ shadow1229_player_016/io_in[7] shadow1229_player_016/io_out[0] shadow1229_player_016/io_out[1]
+ shadow1229_player_016/io_out[2] shadow1229_player_016/io_out[3] shadow1229_player_016/io_out[4]
+ shadow1229_player_016/io_out[5] shadow1229_player_016/io_out[6] shadow1229_player_016/io_out[7]
+ scanchain_016/scan_select_in scanchain_017/scan_select_in vccd1 vssd1 scanchain
Xscanchain_005 scanchain_005/clk_in scanchain_006/clk_in scanchain_005/data_in scanchain_006/data_in
+ scanchain_005/latch_enable_in scanchain_006/latch_enable_in scanchain_005/module_data_in[0]
+ scanchain_005/module_data_in[1] scanchain_005/module_data_in[2] scanchain_005/module_data_in[3]
+ scanchain_005/module_data_in[4] scanchain_005/module_data_in[5] scanchain_005/module_data_in[6]
+ scanchain_005/module_data_in[7] scanchain_005/module_data_out[0] scanchain_005/module_data_out[1]
+ scanchain_005/module_data_out[2] scanchain_005/module_data_out[3] scanchain_005/module_data_out[4]
+ scanchain_005/module_data_out[5] scanchain_005/module_data_out[6] scanchain_005/module_data_out[7]
+ scanchain_005/scan_select_in scanchain_006/scan_select_in vccd1 vssd1 scanchain
Xscanchain_027 scanchain_027/clk_in scanchain_028/clk_in scanchain_027/data_in scanchain_028/data_in
+ scanchain_027/latch_enable_in scanchain_028/latch_enable_in scanchain_027/module_data_in[0]
+ scanchain_027/module_data_in[1] scanchain_027/module_data_in[2] scanchain_027/module_data_in[3]
+ scanchain_027/module_data_in[4] scanchain_027/module_data_in[5] scanchain_027/module_data_in[6]
+ scanchain_027/module_data_in[7] scanchain_027/module_data_out[0] scanchain_027/module_data_out[1]
+ scanchain_027/module_data_out[2] scanchain_027/module_data_out[3] scanchain_027/module_data_out[4]
+ scanchain_027/module_data_out[5] scanchain_027/module_data_out[6] scanchain_027/module_data_out[7]
+ scanchain_027/scan_select_in scanchain_028/scan_select_in vccd1 vssd1 scanchain
Xscanchain_038 scanchain_038/clk_in scanchain_039/clk_in scanchain_038/data_in scanchain_039/data_in
+ scanchain_038/latch_enable_in scanchain_039/latch_enable_in scanchain_038/module_data_in[0]
+ scanchain_038/module_data_in[1] scanchain_038/module_data_in[2] scanchain_038/module_data_in[3]
+ scanchain_038/module_data_in[4] scanchain_038/module_data_in[5] scanchain_038/module_data_in[6]
+ scanchain_038/module_data_in[7] scanchain_038/module_data_out[0] scanchain_038/module_data_out[1]
+ scanchain_038/module_data_out[2] scanchain_038/module_data_out[3] scanchain_038/module_data_out[4]
+ scanchain_038/module_data_out[5] scanchain_038/module_data_out[6] scanchain_038/module_data_out[7]
+ scanchain_038/scan_select_in scanchain_039/scan_select_in vccd1 vssd1 scanchain
Xuser_module_361728533238569985_198 scanchain_198/module_data_in[0] scanchain_198/module_data_in[1]
+ scanchain_198/module_data_in[2] scanchain_198/module_data_in[3] scanchain_198/module_data_in[4]
+ scanchain_198/module_data_in[5] scanchain_198/module_data_in[6] scanchain_198/module_data_in[7]
+ scanchain_198/module_data_out[0] scanchain_198/module_data_out[1] scanchain_198/module_data_out[2]
+ scanchain_198/module_data_out[3] scanchain_198/module_data_out[4] scanchain_198/module_data_out[5]
+ scanchain_198/module_data_out[6] scanchain_198/module_data_out[7] vccd1 vssd1 user_module_361728533238569985
Xscanchain_049 scanchain_049/clk_in scanchain_050/clk_in scanchain_049/data_in scanchain_050/data_in
+ scanchain_049/latch_enable_in scanchain_050/latch_enable_in dsp_4bits_seq_alu_049/io_in[0]
+ dsp_4bits_seq_alu_049/io_in[1] dsp_4bits_seq_alu_049/io_in[2] dsp_4bits_seq_alu_049/io_in[3]
+ dsp_4bits_seq_alu_049/io_in[4] dsp_4bits_seq_alu_049/io_in[5] dsp_4bits_seq_alu_049/io_in[6]
+ dsp_4bits_seq_alu_049/io_in[7] dsp_4bits_seq_alu_049/io_out[0] dsp_4bits_seq_alu_049/io_out[1]
+ dsp_4bits_seq_alu_049/io_out[2] dsp_4bits_seq_alu_049/io_out[3] dsp_4bits_seq_alu_049/io_out[4]
+ dsp_4bits_seq_alu_049/io_out[5] dsp_4bits_seq_alu_049/io_out[6] dsp_4bits_seq_alu_049/io_out[7]
+ scanchain_049/scan_select_in scanchain_050/scan_select_in vccd1 vssd1 scanchain
Xuser_module_361728533238569985_187 scanchain_187/module_data_in[0] scanchain_187/module_data_in[1]
+ scanchain_187/module_data_in[2] scanchain_187/module_data_in[3] scanchain_187/module_data_in[4]
+ scanchain_187/module_data_in[5] scanchain_187/module_data_in[6] scanchain_187/module_data_in[7]
+ scanchain_187/module_data_out[0] scanchain_187/module_data_out[1] scanchain_187/module_data_out[2]
+ scanchain_187/module_data_out[3] scanchain_187/module_data_out[4] scanchain_187/module_data_out[5]
+ scanchain_187/module_data_out[6] scanchain_187/module_data_out[7] vccd1 vssd1 user_module_361728533238569985
Xuser_module_361728533238569985_176 scanchain_176/module_data_in[0] scanchain_176/module_data_in[1]
+ scanchain_176/module_data_in[2] scanchain_176/module_data_in[3] scanchain_176/module_data_in[4]
+ scanchain_176/module_data_in[5] scanchain_176/module_data_in[6] scanchain_176/module_data_in[7]
+ scanchain_176/module_data_out[0] scanchain_176/module_data_out[1] scanchain_176/module_data_out[2]
+ scanchain_176/module_data_out[3] scanchain_176/module_data_out[4] scanchain_176/module_data_out[5]
+ scanchain_176/module_data_out[6] scanchain_176/module_data_out[7] vccd1 vssd1 user_module_361728533238569985
Xuser_module_361728533238569985_165 scanchain_165/module_data_in[0] scanchain_165/module_data_in[1]
+ scanchain_165/module_data_in[2] scanchain_165/module_data_in[3] scanchain_165/module_data_in[4]
+ scanchain_165/module_data_in[5] scanchain_165/module_data_in[6] scanchain_165/module_data_in[7]
+ scanchain_165/module_data_out[0] scanchain_165/module_data_out[1] scanchain_165/module_data_out[2]
+ scanchain_165/module_data_out[3] scanchain_165/module_data_out[4] scanchain_165/module_data_out[5]
+ scanchain_165/module_data_out[6] scanchain_165/module_data_out[7] vccd1 vssd1 user_module_361728533238569985
Xuser_module_361728533238569985_154 scanchain_154/module_data_in[0] scanchain_154/module_data_in[1]
+ scanchain_154/module_data_in[2] scanchain_154/module_data_in[3] scanchain_154/module_data_in[4]
+ scanchain_154/module_data_in[5] scanchain_154/module_data_in[6] scanchain_154/module_data_in[7]
+ scanchain_154/module_data_out[0] scanchain_154/module_data_out[1] scanchain_154/module_data_out[2]
+ scanchain_154/module_data_out[3] scanchain_154/module_data_out[4] scanchain_154/module_data_out[5]
+ scanchain_154/module_data_out[6] scanchain_154/module_data_out[7] vccd1 vssd1 user_module_361728533238569985
Xuser_module_358970514554149889_006 scanchain_006/module_data_in[0] scanchain_006/module_data_in[1]
+ scanchain_006/module_data_in[2] scanchain_006/module_data_in[3] scanchain_006/module_data_in[4]
+ scanchain_006/module_data_in[5] scanchain_006/module_data_in[6] scanchain_006/module_data_in[7]
+ scanchain_006/module_data_out[0] scanchain_006/module_data_out[1] scanchain_006/module_data_out[2]
+ scanchain_006/module_data_out[3] scanchain_006/module_data_out[4] scanchain_006/module_data_out[5]
+ scanchain_006/module_data_out[6] scanchain_006/module_data_out[7] vccd1 vssd1 user_module_358970514554149889
XFSM_LAT_060 FSM_LAT_060/io_in[0] FSM_LAT_060/io_in[1] FSM_LAT_060/io_in[2] FSM_LAT_060/io_in[3]
+ FSM_LAT_060/io_in[4] FSM_LAT_060/io_in[5] FSM_LAT_060/io_in[6] FSM_LAT_060/io_in[7]
+ FSM_LAT_060/io_out[0] FSM_LAT_060/io_out[1] FSM_LAT_060/io_out[2] FSM_LAT_060/io_out[3]
+ FSM_LAT_060/io_out[4] FSM_LAT_060/io_out[5] FSM_LAT_060/io_out[6] FSM_LAT_060/io_out[7]
+ vccd1 vssd1 FSM_LAT
Xpwm_050 pwm_050/io_in[0] pwm_050/io_in[1] pwm_050/io_in[2] pwm_050/io_in[3] pwm_050/io_in[4]
+ pwm_050/io_in[5] pwm_050/io_in[6] pwm_050/io_in[7] pwm_050/io_out[0] pwm_050/io_out[1]
+ pwm_050/io_out[2] pwm_050/io_out[3] pwm_050/io_out[4] pwm_050/io_out[5] pwm_050/io_out[6]
+ pwm_050/io_out[7] vccd1 vssd1 pwm
Xscanchain_209 scanchain_209/clk_in scanchain_210/clk_in scanchain_209/data_in scanchain_210/data_in
+ scanchain_209/latch_enable_in scanchain_210/latch_enable_in scanchain_209/module_data_in[0]
+ scanchain_209/module_data_in[1] scanchain_209/module_data_in[2] scanchain_209/module_data_in[3]
+ scanchain_209/module_data_in[4] scanchain_209/module_data_in[5] scanchain_209/module_data_in[6]
+ scanchain_209/module_data_in[7] scanchain_209/module_data_out[0] scanchain_209/module_data_out[1]
+ scanchain_209/module_data_out[2] scanchain_209/module_data_out[3] scanchain_209/module_data_out[4]
+ scanchain_209/module_data_out[5] scanchain_209/module_data_out[6] scanchain_209/module_data_out[7]
+ scanchain_209/scan_select_in scanchain_210/scan_select_in vccd1 vssd1 scanchain
Xuser_module_361728533238569985_122 scanchain_122/module_data_in[0] scanchain_122/module_data_in[1]
+ scanchain_122/module_data_in[2] scanchain_122/module_data_in[3] scanchain_122/module_data_in[4]
+ scanchain_122/module_data_in[5] scanchain_122/module_data_in[6] scanchain_122/module_data_in[7]
+ scanchain_122/module_data_out[0] scanchain_122/module_data_out[1] scanchain_122/module_data_out[2]
+ scanchain_122/module_data_out[3] scanchain_122/module_data_out[4] scanchain_122/module_data_out[5]
+ scanchain_122/module_data_out[6] scanchain_122/module_data_out[7] vccd1 vssd1 user_module_361728533238569985
Xuser_module_361728533238569985_133 scanchain_133/module_data_in[0] scanchain_133/module_data_in[1]
+ scanchain_133/module_data_in[2] scanchain_133/module_data_in[3] scanchain_133/module_data_in[4]
+ scanchain_133/module_data_in[5] scanchain_133/module_data_in[6] scanchain_133/module_data_in[7]
+ scanchain_133/module_data_out[0] scanchain_133/module_data_out[1] scanchain_133/module_data_out[2]
+ scanchain_133/module_data_out[3] scanchain_133/module_data_out[4] scanchain_133/module_data_out[5]
+ scanchain_133/module_data_out[6] scanchain_133/module_data_out[7] vccd1 vssd1 user_module_361728533238569985
Xuser_module_361728533238569985_111 scanchain_111/module_data_in[0] scanchain_111/module_data_in[1]
+ scanchain_111/module_data_in[2] scanchain_111/module_data_in[3] scanchain_111/module_data_in[4]
+ scanchain_111/module_data_in[5] scanchain_111/module_data_in[6] scanchain_111/module_data_in[7]
+ scanchain_111/module_data_out[0] scanchain_111/module_data_out[1] scanchain_111/module_data_out[2]
+ scanchain_111/module_data_out[3] scanchain_111/module_data_out[4] scanchain_111/module_data_out[5]
+ scanchain_111/module_data_out[6] scanchain_111/module_data_out[7] vccd1 vssd1 user_module_361728533238569985
Xuser_module_361728533238569985_144 scanchain_144/module_data_in[0] scanchain_144/module_data_in[1]
+ scanchain_144/module_data_in[2] scanchain_144/module_data_in[3] scanchain_144/module_data_in[4]
+ scanchain_144/module_data_in[5] scanchain_144/module_data_in[6] scanchain_144/module_data_in[7]
+ scanchain_144/module_data_out[0] scanchain_144/module_data_out[1] scanchain_144/module_data_out[2]
+ scanchain_144/module_data_out[3] scanchain_144/module_data_out[4] scanchain_144/module_data_out[5]
+ scanchain_144/module_data_out[6] scanchain_144/module_data_out[7] vccd1 vssd1 user_module_361728533238569985
Xuser_module_361728533238569985_100 scanchain_100/module_data_in[0] scanchain_100/module_data_in[1]
+ scanchain_100/module_data_in[2] scanchain_100/module_data_in[3] scanchain_100/module_data_in[4]
+ scanchain_100/module_data_in[5] scanchain_100/module_data_in[6] scanchain_100/module_data_in[7]
+ scanchain_100/module_data_out[0] scanchain_100/module_data_out[1] scanchain_100/module_data_out[2]
+ scanchain_100/module_data_out[3] scanchain_100/module_data_out[4] scanchain_100/module_data_out[5]
+ scanchain_100/module_data_out[6] scanchain_100/module_data_out[7] vccd1 vssd1 user_module_361728533238569985
Xscanchain_017 scanchain_017/clk_in scanchain_018/clk_in scanchain_017/data_in scanchain_018/data_in
+ scanchain_017/latch_enable_in scanchain_018/latch_enable_in scanchain_017/module_data_in[0]
+ scanchain_017/module_data_in[1] scanchain_017/module_data_in[2] scanchain_017/module_data_in[3]
+ scanchain_017/module_data_in[4] scanchain_017/module_data_in[5] scanchain_017/module_data_in[6]
+ scanchain_017/module_data_in[7] scanchain_017/module_data_out[0] scanchain_017/module_data_out[1]
+ scanchain_017/module_data_out[2] scanchain_017/module_data_out[3] scanchain_017/module_data_out[4]
+ scanchain_017/module_data_out[5] scanchain_017/module_data_out[6] scanchain_017/module_data_out[7]
+ scanchain_017/scan_select_in scanchain_018/scan_select_in vccd1 vssd1 scanchain
Xscanchain_006 scanchain_006/clk_in scanchain_007/clk_in scanchain_006/data_in scanchain_007/data_in
+ scanchain_006/latch_enable_in scanchain_007/latch_enable_in scanchain_006/module_data_in[0]
+ scanchain_006/module_data_in[1] scanchain_006/module_data_in[2] scanchain_006/module_data_in[3]
+ scanchain_006/module_data_in[4] scanchain_006/module_data_in[5] scanchain_006/module_data_in[6]
+ scanchain_006/module_data_in[7] scanchain_006/module_data_out[0] scanchain_006/module_data_out[1]
+ scanchain_006/module_data_out[2] scanchain_006/module_data_out[3] scanchain_006/module_data_out[4]
+ scanchain_006/module_data_out[5] scanchain_006/module_data_out[6] scanchain_006/module_data_out[7]
+ scanchain_006/scan_select_in scanchain_007/scan_select_in vccd1 vssd1 scanchain
Xscanchain_028 scanchain_028/clk_in scanchain_029/clk_in scanchain_028/data_in scanchain_029/data_in
+ scanchain_028/latch_enable_in scanchain_029/latch_enable_in scanchain_028/module_data_in[0]
+ scanchain_028/module_data_in[1] scanchain_028/module_data_in[2] scanchain_028/module_data_in[3]
+ scanchain_028/module_data_in[4] scanchain_028/module_data_in[5] scanchain_028/module_data_in[6]
+ scanchain_028/module_data_in[7] scanchain_028/module_data_out[0] scanchain_028/module_data_out[1]
+ scanchain_028/module_data_out[2] scanchain_028/module_data_out[3] scanchain_028/module_data_out[4]
+ scanchain_028/module_data_out[5] scanchain_028/module_data_out[6] scanchain_028/module_data_out[7]
+ scanchain_028/scan_select_in scanchain_029/scan_select_in vccd1 vssd1 scanchain
Xscanchain_039 scanchain_039/clk_in scanchain_040/clk_in scanchain_039/data_in scanchain_040/data_in
+ scanchain_039/latch_enable_in scanchain_040/latch_enable_in tinysat_039/io_in[0]
+ tinysat_039/io_in[1] tinysat_039/io_in[2] tinysat_039/io_in[3] tinysat_039/io_in[4]
+ tinysat_039/io_in[5] tinysat_039/io_in[6] tinysat_039/io_in[7] tinysat_039/io_out[0]
+ tinysat_039/io_out[1] tinysat_039/io_out[2] tinysat_039/io_out[3] tinysat_039/io_out[4]
+ tinysat_039/io_out[5] tinysat_039/io_out[6] tinysat_039/io_out[7] scanchain_039/scan_select_in
+ scanchain_040/scan_select_in vccd1 vssd1 scanchain
Xuser_module_361728533238569985_199 scanchain_199/module_data_in[0] scanchain_199/module_data_in[1]
+ scanchain_199/module_data_in[2] scanchain_199/module_data_in[3] scanchain_199/module_data_in[4]
+ scanchain_199/module_data_in[5] scanchain_199/module_data_in[6] scanchain_199/module_data_in[7]
+ scanchain_199/module_data_out[0] scanchain_199/module_data_out[1] scanchain_199/module_data_out[2]
+ scanchain_199/module_data_out[3] scanchain_199/module_data_out[4] scanchain_199/module_data_out[5]
+ scanchain_199/module_data_out[6] scanchain_199/module_data_out[7] vccd1 vssd1 user_module_361728533238569985
Xuser_module_361728533238569985_188 scanchain_188/module_data_in[0] scanchain_188/module_data_in[1]
+ scanchain_188/module_data_in[2] scanchain_188/module_data_in[3] scanchain_188/module_data_in[4]
+ scanchain_188/module_data_in[5] scanchain_188/module_data_in[6] scanchain_188/module_data_in[7]
+ scanchain_188/module_data_out[0] scanchain_188/module_data_out[1] scanchain_188/module_data_out[2]
+ scanchain_188/module_data_out[3] scanchain_188/module_data_out[4] scanchain_188/module_data_out[5]
+ scanchain_188/module_data_out[6] scanchain_188/module_data_out[7] vccd1 vssd1 user_module_361728533238569985
Xuser_module_361728533238569985_177 scanchain_177/module_data_in[0] scanchain_177/module_data_in[1]
+ scanchain_177/module_data_in[2] scanchain_177/module_data_in[3] scanchain_177/module_data_in[4]
+ scanchain_177/module_data_in[5] scanchain_177/module_data_in[6] scanchain_177/module_data_in[7]
+ scanchain_177/module_data_out[0] scanchain_177/module_data_out[1] scanchain_177/module_data_out[2]
+ scanchain_177/module_data_out[3] scanchain_177/module_data_out[4] scanchain_177/module_data_out[5]
+ scanchain_177/module_data_out[6] scanchain_177/module_data_out[7] vccd1 vssd1 user_module_361728533238569985
Xuser_module_361728533238569985_166 scanchain_166/module_data_in[0] scanchain_166/module_data_in[1]
+ scanchain_166/module_data_in[2] scanchain_166/module_data_in[3] scanchain_166/module_data_in[4]
+ scanchain_166/module_data_in[5] scanchain_166/module_data_in[6] scanchain_166/module_data_in[7]
+ scanchain_166/module_data_out[0] scanchain_166/module_data_out[1] scanchain_166/module_data_out[2]
+ scanchain_166/module_data_out[3] scanchain_166/module_data_out[4] scanchain_166/module_data_out[5]
+ scanchain_166/module_data_out[6] scanchain_166/module_data_out[7] vccd1 vssd1 user_module_361728533238569985
Xuser_module_361728533238569985_155 scanchain_155/module_data_in[0] scanchain_155/module_data_in[1]
+ scanchain_155/module_data_in[2] scanchain_155/module_data_in[3] scanchain_155/module_data_in[4]
+ scanchain_155/module_data_in[5] scanchain_155/module_data_in[6] scanchain_155/module_data_in[7]
+ scanchain_155/module_data_out[0] scanchain_155/module_data_out[1] scanchain_155/module_data_out[2]
+ scanchain_155/module_data_out[3] scanchain_155/module_data_out[4] scanchain_155/module_data_out[5]
+ scanchain_155/module_data_out[6] scanchain_155/module_data_out[7] vccd1 vssd1 user_module_361728533238569985
Xuser_module_361728533238569985_123 scanchain_123/module_data_in[0] scanchain_123/module_data_in[1]
+ scanchain_123/module_data_in[2] scanchain_123/module_data_in[3] scanchain_123/module_data_in[4]
+ scanchain_123/module_data_in[5] scanchain_123/module_data_in[6] scanchain_123/module_data_in[7]
+ scanchain_123/module_data_out[0] scanchain_123/module_data_out[1] scanchain_123/module_data_out[2]
+ scanchain_123/module_data_out[3] scanchain_123/module_data_out[4] scanchain_123/module_data_out[5]
+ scanchain_123/module_data_out[6] scanchain_123/module_data_out[7] vccd1 vssd1 user_module_361728533238569985
Xuser_module_361728533238569985_134 scanchain_134/module_data_in[0] scanchain_134/module_data_in[1]
+ scanchain_134/module_data_in[2] scanchain_134/module_data_in[3] scanchain_134/module_data_in[4]
+ scanchain_134/module_data_in[5] scanchain_134/module_data_in[6] scanchain_134/module_data_in[7]
+ scanchain_134/module_data_out[0] scanchain_134/module_data_out[1] scanchain_134/module_data_out[2]
+ scanchain_134/module_data_out[3] scanchain_134/module_data_out[4] scanchain_134/module_data_out[5]
+ scanchain_134/module_data_out[6] scanchain_134/module_data_out[7] vccd1 vssd1 user_module_361728533238569985
Xuser_module_361728533238569985_112 scanchain_112/module_data_in[0] scanchain_112/module_data_in[1]
+ scanchain_112/module_data_in[2] scanchain_112/module_data_in[3] scanchain_112/module_data_in[4]
+ scanchain_112/module_data_in[5] scanchain_112/module_data_in[6] scanchain_112/module_data_in[7]
+ scanchain_112/module_data_out[0] scanchain_112/module_data_out[1] scanchain_112/module_data_out[2]
+ scanchain_112/module_data_out[3] scanchain_112/module_data_out[4] scanchain_112/module_data_out[5]
+ scanchain_112/module_data_out[6] scanchain_112/module_data_out[7] vccd1 vssd1 user_module_361728533238569985
Xuser_module_361728533238569985_145 scanchain_145/module_data_in[0] scanchain_145/module_data_in[1]
+ scanchain_145/module_data_in[2] scanchain_145/module_data_in[3] scanchain_145/module_data_in[4]
+ scanchain_145/module_data_in[5] scanchain_145/module_data_in[6] scanchain_145/module_data_in[7]
+ scanchain_145/module_data_out[0] scanchain_145/module_data_out[1] scanchain_145/module_data_out[2]
+ scanchain_145/module_data_out[3] scanchain_145/module_data_out[4] scanchain_145/module_data_out[5]
+ scanchain_145/module_data_out[6] scanchain_145/module_data_out[7] vccd1 vssd1 user_module_361728533238569985
Xuser_module_361728533238569985_101 scanchain_101/module_data_in[0] scanchain_101/module_data_in[1]
+ scanchain_101/module_data_in[2] scanchain_101/module_data_in[3] scanchain_101/module_data_in[4]
+ scanchain_101/module_data_in[5] scanchain_101/module_data_in[6] scanchain_101/module_data_in[7]
+ scanchain_101/module_data_out[0] scanchain_101/module_data_out[1] scanchain_101/module_data_out[2]
+ scanchain_101/module_data_out[3] scanchain_101/module_data_out[4] scanchain_101/module_data_out[5]
+ scanchain_101/module_data_out[6] scanchain_101/module_data_out[7] vccd1 vssd1 user_module_361728533238569985
Xscanchain_018 scanchain_018/clk_in scanchain_019/clk_in scanchain_018/data_in scanchain_019/data_in
+ scanchain_018/latch_enable_in scanchain_019/latch_enable_in scanchain_018/module_data_in[0]
+ scanchain_018/module_data_in[1] scanchain_018/module_data_in[2] scanchain_018/module_data_in[3]
+ scanchain_018/module_data_in[4] scanchain_018/module_data_in[5] scanchain_018/module_data_in[6]
+ scanchain_018/module_data_in[7] scanchain_018/module_data_out[0] scanchain_018/module_data_out[1]
+ scanchain_018/module_data_out[2] scanchain_018/module_data_out[3] scanchain_018/module_data_out[4]
+ scanchain_018/module_data_out[5] scanchain_018/module_data_out[6] scanchain_018/module_data_out[7]
+ scanchain_018/scan_select_in scanchain_019/scan_select_in vccd1 vssd1 scanchain
Xscanchain_007 scanchain_007/clk_in scanchain_008/clk_in scanchain_007/data_in scanchain_008/data_in
+ scanchain_007/latch_enable_in scanchain_008/latch_enable_in scanchain_007/module_data_in[0]
+ scanchain_007/module_data_in[1] scanchain_007/module_data_in[2] scanchain_007/module_data_in[3]
+ scanchain_007/module_data_in[4] scanchain_007/module_data_in[5] scanchain_007/module_data_in[6]
+ scanchain_007/module_data_in[7] scanchain_007/module_data_out[0] scanchain_007/module_data_out[1]
+ scanchain_007/module_data_out[2] scanchain_007/module_data_out[3] scanchain_007/module_data_out[4]
+ scanchain_007/module_data_out[5] scanchain_007/module_data_out[6] scanchain_007/module_data_out[7]
+ scanchain_007/scan_select_in scanchain_008/scan_select_in vccd1 vssd1 scanchain
Xscanchain_029 scanchain_029/clk_in scanchain_030/clk_in scanchain_029/data_in scanchain_030/data_in
+ scanchain_029/latch_enable_in scanchain_030/latch_enable_in scanchain_029/module_data_in[0]
+ scanchain_029/module_data_in[1] scanchain_029/module_data_in[2] scanchain_029/module_data_in[3]
+ scanchain_029/module_data_in[4] scanchain_029/module_data_in[5] scanchain_029/module_data_in[6]
+ scanchain_029/module_data_in[7] scanchain_029/module_data_out[0] scanchain_029/module_data_out[1]
+ scanchain_029/module_data_out[2] scanchain_029/module_data_out[3] scanchain_029/module_data_out[4]
+ scanchain_029/module_data_out[5] scanchain_029/module_data_out[6] scanchain_029/module_data_out[7]
+ scanchain_029/scan_select_in scanchain_030/scan_select_in vccd1 vssd1 scanchain
Xuser_module_361728533238569985_189 scanchain_189/module_data_in[0] scanchain_189/module_data_in[1]
+ scanchain_189/module_data_in[2] scanchain_189/module_data_in[3] scanchain_189/module_data_in[4]
+ scanchain_189/module_data_in[5] scanchain_189/module_data_in[6] scanchain_189/module_data_in[7]
+ scanchain_189/module_data_out[0] scanchain_189/module_data_out[1] scanchain_189/module_data_out[2]
+ scanchain_189/module_data_out[3] scanchain_189/module_data_out[4] scanchain_189/module_data_out[5]
+ scanchain_189/module_data_out[6] scanchain_189/module_data_out[7] vccd1 vssd1 user_module_361728533238569985
Xuser_module_361728533238569985_178 scanchain_178/module_data_in[0] scanchain_178/module_data_in[1]
+ scanchain_178/module_data_in[2] scanchain_178/module_data_in[3] scanchain_178/module_data_in[4]
+ scanchain_178/module_data_in[5] scanchain_178/module_data_in[6] scanchain_178/module_data_in[7]
+ scanchain_178/module_data_out[0] scanchain_178/module_data_out[1] scanchain_178/module_data_out[2]
+ scanchain_178/module_data_out[3] scanchain_178/module_data_out[4] scanchain_178/module_data_out[5]
+ scanchain_178/module_data_out[6] scanchain_178/module_data_out[7] vccd1 vssd1 user_module_361728533238569985
Xuser_module_361728533238569985_167 scanchain_167/module_data_in[0] scanchain_167/module_data_in[1]
+ scanchain_167/module_data_in[2] scanchain_167/module_data_in[3] scanchain_167/module_data_in[4]
+ scanchain_167/module_data_in[5] scanchain_167/module_data_in[6] scanchain_167/module_data_in[7]
+ scanchain_167/module_data_out[0] scanchain_167/module_data_out[1] scanchain_167/module_data_out[2]
+ scanchain_167/module_data_out[3] scanchain_167/module_data_out[4] scanchain_167/module_data_out[5]
+ scanchain_167/module_data_out[6] scanchain_167/module_data_out[7] vccd1 vssd1 user_module_361728533238569985
Xuser_module_361728533238569985_156 scanchain_156/module_data_in[0] scanchain_156/module_data_in[1]
+ scanchain_156/module_data_in[2] scanchain_156/module_data_in[3] scanchain_156/module_data_in[4]
+ scanchain_156/module_data_in[5] scanchain_156/module_data_in[6] scanchain_156/module_data_in[7]
+ scanchain_156/module_data_out[0] scanchain_156/module_data_out[1] scanchain_156/module_data_out[2]
+ scanchain_156/module_data_out[3] scanchain_156/module_data_out[4] scanchain_156/module_data_out[5]
+ scanchain_156/module_data_out[6] scanchain_156/module_data_out[7] vccd1 vssd1 user_module_361728533238569985
Xscan_controller io_in[12] io_in[13] io_in[14] io_in[15] io_in[16] io_in[17] io_in[18]
+ io_in[19] io_in[20] wb_clk_i io_in[8] io_in[9] io_in[21] io_in[22] io_in[23] io_in[24]
+ io_in[25] io_in[26] io_in[27] io_in[28] la_data_in[0] la_data_in[1] la_data_out[0]
+ la_data_in[3] la_data_in[2] io_oeb[0] io_oeb[10] io_oeb[11] io_oeb[12] io_oeb[13]
+ io_oeb[14] io_oeb[15] io_oeb[16] io_oeb[17] io_oeb[18] io_oeb[19] io_oeb[1] io_oeb[20]
+ io_oeb[21] io_oeb[22] io_oeb[23] io_oeb[24] io_oeb[25] io_oeb[26] io_oeb[27] io_oeb[28]
+ io_oeb[29] io_oeb[2] io_oeb[30] io_oeb[31] io_oeb[32] io_oeb[33] io_oeb[34] io_oeb[35]
+ io_oeb[36] io_oeb[37] io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7] io_oeb[8]
+ io_oeb[9] io_out[29] io_out[30] io_out[31] io_out[32] io_out[33] io_out[34] io_out[35]
+ io_out[36] io_out[37] wb_rst_i scanchain_249/clk_out scanchain_000/clk_in scanchain_249/data_out
+ scanchain_000/data_in scanchain_000/latch_enable_in scan_controller/scan_select
+ io_in[11] io_out[10] vccd1 vssd1 scan_controller
Xuser_module_362379207695863809_082 scanchain_082/module_data_in[0] scanchain_082/module_data_in[1]
+ scanchain_082/module_data_in[2] scanchain_082/module_data_in[3] scanchain_082/module_data_in[4]
+ scanchain_082/module_data_in[5] scanchain_082/module_data_in[6] scanchain_082/module_data_in[7]
+ scanchain_082/module_data_out[0] scanchain_082/module_data_out[1] scanchain_082/module_data_out[2]
+ scanchain_082/module_data_out[3] scanchain_082/module_data_out[4] scanchain_082/module_data_out[5]
+ scanchain_082/module_data_out[6] scanchain_082/module_data_out[7] vccd1 vssd1 user_module_362379207695863809
Xuser_module_359387860730498049_015 scanchain_015/module_data_in[0] scanchain_015/module_data_in[1]
+ scanchain_015/module_data_in[2] scanchain_015/module_data_in[3] scanchain_015/module_data_in[4]
+ scanchain_015/module_data_in[5] scanchain_015/module_data_in[6] scanchain_015/module_data_in[7]
+ scanchain_015/module_data_out[0] scanchain_015/module_data_out[1] scanchain_015/module_data_out[2]
+ scanchain_015/module_data_out[3] scanchain_015/module_data_out[4] scanchain_015/module_data_out[5]
+ scanchain_015/module_data_out[6] scanchain_015/module_data_out[7] vccd1 vssd1 user_module_359387860730498049
Xscanchain_190 scanchain_190/clk_in scanchain_191/clk_in scanchain_190/data_in scanchain_191/data_in
+ scanchain_190/latch_enable_in scanchain_191/latch_enable_in scanchain_190/module_data_in[0]
+ scanchain_190/module_data_in[1] scanchain_190/module_data_in[2] scanchain_190/module_data_in[3]
+ scanchain_190/module_data_in[4] scanchain_190/module_data_in[5] scanchain_190/module_data_in[6]
+ scanchain_190/module_data_in[7] scanchain_190/module_data_out[0] scanchain_190/module_data_out[1]
+ scanchain_190/module_data_out[2] scanchain_190/module_data_out[3] scanchain_190/module_data_out[4]
+ scanchain_190/module_data_out[5] scanchain_190/module_data_out[6] scanchain_190/module_data_out[7]
+ scanchain_190/scan_select_in scanchain_191/scan_select_in vccd1 vssd1 scanchain
Xnikor_clock_035 nikor_clock_035/io_in[0] nikor_clock_035/io_in[1] nikor_clock_035/io_in[2]
+ nikor_clock_035/io_in[3] nikor_clock_035/io_in[4] nikor_clock_035/io_in[5] nikor_clock_035/io_in[6]
+ nikor_clock_035/io_in[7] nikor_clock_035/io_out[0] nikor_clock_035/io_out[1] nikor_clock_035/io_out[2]
+ nikor_clock_035/io_out[3] nikor_clock_035/io_out[4] nikor_clock_035/io_out[5] nikor_clock_035/io_out[6]
+ nikor_clock_035/io_out[7] vccd1 vssd1 nikor_clock
Xgranth_crc_decelerator_034 scanchain_034/module_data_in[0] scanchain_034/module_data_in[1]
+ scanchain_034/module_data_in[2] scanchain_034/module_data_in[3] scanchain_034/module_data_in[4]
+ scanchain_034/module_data_in[5] scanchain_034/module_data_in[6] scanchain_034/module_data_in[7]
+ scanchain_034/module_data_out[0] scanchain_034/module_data_out[1] scanchain_034/module_data_out[2]
+ scanchain_034/module_data_out[3] scanchain_034/module_data_out[4] scanchain_034/module_data_out[5]
+ scanchain_034/module_data_out[6] scanchain_034/module_data_out[7] vccd1 vssd1 granth_crc_decelerator
Xuser_module_361728533238569985_124 scanchain_124/module_data_in[0] scanchain_124/module_data_in[1]
+ scanchain_124/module_data_in[2] scanchain_124/module_data_in[3] scanchain_124/module_data_in[4]
+ scanchain_124/module_data_in[5] scanchain_124/module_data_in[6] scanchain_124/module_data_in[7]
+ scanchain_124/module_data_out[0] scanchain_124/module_data_out[1] scanchain_124/module_data_out[2]
+ scanchain_124/module_data_out[3] scanchain_124/module_data_out[4] scanchain_124/module_data_out[5]
+ scanchain_124/module_data_out[6] scanchain_124/module_data_out[7] vccd1 vssd1 user_module_361728533238569985
Xuser_module_361728533238569985_135 scanchain_135/module_data_in[0] scanchain_135/module_data_in[1]
+ scanchain_135/module_data_in[2] scanchain_135/module_data_in[3] scanchain_135/module_data_in[4]
+ scanchain_135/module_data_in[5] scanchain_135/module_data_in[6] scanchain_135/module_data_in[7]
+ scanchain_135/module_data_out[0] scanchain_135/module_data_out[1] scanchain_135/module_data_out[2]
+ scanchain_135/module_data_out[3] scanchain_135/module_data_out[4] scanchain_135/module_data_out[5]
+ scanchain_135/module_data_out[6] scanchain_135/module_data_out[7] vccd1 vssd1 user_module_361728533238569985
Xuser_module_361728533238569985_113 scanchain_113/module_data_in[0] scanchain_113/module_data_in[1]
+ scanchain_113/module_data_in[2] scanchain_113/module_data_in[3] scanchain_113/module_data_in[4]
+ scanchain_113/module_data_in[5] scanchain_113/module_data_in[6] scanchain_113/module_data_in[7]
+ scanchain_113/module_data_out[0] scanchain_113/module_data_out[1] scanchain_113/module_data_out[2]
+ scanchain_113/module_data_out[3] scanchain_113/module_data_out[4] scanchain_113/module_data_out[5]
+ scanchain_113/module_data_out[6] scanchain_113/module_data_out[7] vccd1 vssd1 user_module_361728533238569985
Xuser_module_361728533238569985_146 scanchain_146/module_data_in[0] scanchain_146/module_data_in[1]
+ scanchain_146/module_data_in[2] scanchain_146/module_data_in[3] scanchain_146/module_data_in[4]
+ scanchain_146/module_data_in[5] scanchain_146/module_data_in[6] scanchain_146/module_data_in[7]
+ scanchain_146/module_data_out[0] scanchain_146/module_data_out[1] scanchain_146/module_data_out[2]
+ scanchain_146/module_data_out[3] scanchain_146/module_data_out[4] scanchain_146/module_data_out[5]
+ scanchain_146/module_data_out[6] scanchain_146/module_data_out[7] vccd1 vssd1 user_module_361728533238569985
Xuser_module_361728533238569985_102 scanchain_102/module_data_in[0] scanchain_102/module_data_in[1]
+ scanchain_102/module_data_in[2] scanchain_102/module_data_in[3] scanchain_102/module_data_in[4]
+ scanchain_102/module_data_in[5] scanchain_102/module_data_in[6] scanchain_102/module_data_in[7]
+ scanchain_102/module_data_out[0] scanchain_102/module_data_out[1] scanchain_102/module_data_out[2]
+ scanchain_102/module_data_out[3] scanchain_102/module_data_out[4] scanchain_102/module_data_out[5]
+ scanchain_102/module_data_out[6] scanchain_102/module_data_out[7] vccd1 vssd1 user_module_361728533238569985
Xuser_module_361728533238569985_179 scanchain_179/module_data_in[0] scanchain_179/module_data_in[1]
+ scanchain_179/module_data_in[2] scanchain_179/module_data_in[3] scanchain_179/module_data_in[4]
+ scanchain_179/module_data_in[5] scanchain_179/module_data_in[6] scanchain_179/module_data_in[7]
+ scanchain_179/module_data_out[0] scanchain_179/module_data_out[1] scanchain_179/module_data_out[2]
+ scanchain_179/module_data_out[3] scanchain_179/module_data_out[4] scanchain_179/module_data_out[5]
+ scanchain_179/module_data_out[6] scanchain_179/module_data_out[7] vccd1 vssd1 user_module_361728533238569985
Xuser_module_361728533238569985_168 scanchain_168/module_data_in[0] scanchain_168/module_data_in[1]
+ scanchain_168/module_data_in[2] scanchain_168/module_data_in[3] scanchain_168/module_data_in[4]
+ scanchain_168/module_data_in[5] scanchain_168/module_data_in[6] scanchain_168/module_data_in[7]
+ scanchain_168/module_data_out[0] scanchain_168/module_data_out[1] scanchain_168/module_data_out[2]
+ scanchain_168/module_data_out[3] scanchain_168/module_data_out[4] scanchain_168/module_data_out[5]
+ scanchain_168/module_data_out[6] scanchain_168/module_data_out[7] vccd1 vssd1 user_module_361728533238569985
Xuser_module_361728533238569985_157 scanchain_157/module_data_in[0] scanchain_157/module_data_in[1]
+ scanchain_157/module_data_in[2] scanchain_157/module_data_in[3] scanchain_157/module_data_in[4]
+ scanchain_157/module_data_in[5] scanchain_157/module_data_in[6] scanchain_157/module_data_in[7]
+ scanchain_157/module_data_out[0] scanchain_157/module_data_out[1] scanchain_157/module_data_out[2]
+ scanchain_157/module_data_out[3] scanchain_157/module_data_out[4] scanchain_157/module_data_out[5]
+ scanchain_157/module_data_out[6] scanchain_157/module_data_out[7] vccd1 vssd1 user_module_361728533238569985
Xscanchain_019 scanchain_019/clk_in scanchain_020/clk_in scanchain_019/data_in scanchain_020/data_in
+ scanchain_019/latch_enable_in scanchain_020/latch_enable_in moonbase_pdp8_019/io_in[0]
+ moonbase_pdp8_019/io_in[1] moonbase_pdp8_019/io_in[2] moonbase_pdp8_019/io_in[3]
+ moonbase_pdp8_019/io_in[4] moonbase_pdp8_019/io_in[5] moonbase_pdp8_019/io_in[6]
+ moonbase_pdp8_019/io_in[7] moonbase_pdp8_019/io_out[0] moonbase_pdp8_019/io_out[1]
+ moonbase_pdp8_019/io_out[2] moonbase_pdp8_019/io_out[3] moonbase_pdp8_019/io_out[4]
+ moonbase_pdp8_019/io_out[5] moonbase_pdp8_019/io_out[6] moonbase_pdp8_019/io_out[7]
+ scanchain_019/scan_select_in scanchain_020/scan_select_in vccd1 vssd1 scanchain
Xscanchain_008 scanchain_008/clk_in scanchain_009/clk_in scanchain_008/data_in scanchain_009/data_in
+ scanchain_008/latch_enable_in scanchain_009/latch_enable_in scanchain_008/module_data_in[0]
+ scanchain_008/module_data_in[1] scanchain_008/module_data_in[2] scanchain_008/module_data_in[3]
+ scanchain_008/module_data_in[4] scanchain_008/module_data_in[5] scanchain_008/module_data_in[6]
+ scanchain_008/module_data_in[7] scanchain_008/module_data_out[0] scanchain_008/module_data_out[1]
+ scanchain_008/module_data_out[2] scanchain_008/module_data_out[3] scanchain_008/module_data_out[4]
+ scanchain_008/module_data_out[5] scanchain_008/module_data_out[6] scanchain_008/module_data_out[7]
+ scanchain_008/scan_select_in scanchain_009/scan_select_in vccd1 vssd1 scanchain
Xuser_module_359360834113498113_012 scanchain_012/module_data_in[0] scanchain_012/module_data_in[1]
+ scanchain_012/module_data_in[2] scanchain_012/module_data_in[3] scanchain_012/module_data_in[4]
+ scanchain_012/module_data_in[5] scanchain_012/module_data_in[6] scanchain_012/module_data_in[7]
+ scanchain_012/module_data_out[0] scanchain_012/module_data_out[1] scanchain_012/module_data_out[2]
+ scanchain_012/module_data_out[3] scanchain_012/module_data_out[4] scanchain_012/module_data_out[5]
+ scanchain_012/module_data_out[6] scanchain_012/module_data_out[7] vccd1 vssd1 user_module_359360834113498113
Xyannickreiss_dot_op_021 scanchain_021/module_data_in[0] scanchain_021/module_data_in[1]
+ scanchain_021/module_data_in[2] scanchain_021/module_data_in[3] scanchain_021/module_data_in[4]
+ scanchain_021/module_data_in[5] scanchain_021/module_data_in[6] scanchain_021/module_data_in[7]
+ scanchain_021/module_data_out[0] scanchain_021/module_data_out[1] scanchain_021/module_data_out[2]
+ scanchain_021/module_data_out[3] scanchain_021/module_data_out[4] scanchain_021/module_data_out[5]
+ scanchain_021/module_data_out[6] scanchain_021/module_data_out[7] vccd1 vssd1 yannickreiss_dot_op
Xscanchain_191 scanchain_191/clk_in scanchain_192/clk_in scanchain_191/data_in scanchain_192/data_in
+ scanchain_191/latch_enable_in scanchain_192/latch_enable_in scanchain_191/module_data_in[0]
+ scanchain_191/module_data_in[1] scanchain_191/module_data_in[2] scanchain_191/module_data_in[3]
+ scanchain_191/module_data_in[4] scanchain_191/module_data_in[5] scanchain_191/module_data_in[6]
+ scanchain_191/module_data_in[7] scanchain_191/module_data_out[0] scanchain_191/module_data_out[1]
+ scanchain_191/module_data_out[2] scanchain_191/module_data_out[3] scanchain_191/module_data_out[4]
+ scanchain_191/module_data_out[5] scanchain_191/module_data_out[6] scanchain_191/module_data_out[7]
+ scanchain_191/scan_select_in scanchain_192/scan_select_in vccd1 vssd1 scanchain
Xscanchain_180 scanchain_180/clk_in scanchain_181/clk_in scanchain_180/data_in scanchain_181/data_in
+ scanchain_180/latch_enable_in scanchain_181/latch_enable_in scanchain_180/module_data_in[0]
+ scanchain_180/module_data_in[1] scanchain_180/module_data_in[2] scanchain_180/module_data_in[3]
+ scanchain_180/module_data_in[4] scanchain_180/module_data_in[5] scanchain_180/module_data_in[6]
+ scanchain_180/module_data_in[7] scanchain_180/module_data_out[0] scanchain_180/module_data_out[1]
+ scanchain_180/module_data_out[2] scanchain_180/module_data_out[3] scanchain_180/module_data_out[4]
+ scanchain_180/module_data_out[5] scanchain_180/module_data_out[6] scanchain_180/module_data_out[7]
+ scanchain_180/scan_select_in scanchain_181/scan_select_in vccd1 vssd1 scanchain
Xuser_module_361728533238569985_125 scanchain_125/module_data_in[0] scanchain_125/module_data_in[1]
+ scanchain_125/module_data_in[2] scanchain_125/module_data_in[3] scanchain_125/module_data_in[4]
+ scanchain_125/module_data_in[5] scanchain_125/module_data_in[6] scanchain_125/module_data_in[7]
+ scanchain_125/module_data_out[0] scanchain_125/module_data_out[1] scanchain_125/module_data_out[2]
+ scanchain_125/module_data_out[3] scanchain_125/module_data_out[4] scanchain_125/module_data_out[5]
+ scanchain_125/module_data_out[6] scanchain_125/module_data_out[7] vccd1 vssd1 user_module_361728533238569985
Xuser_module_361728533238569985_114 scanchain_114/module_data_in[0] scanchain_114/module_data_in[1]
+ scanchain_114/module_data_in[2] scanchain_114/module_data_in[3] scanchain_114/module_data_in[4]
+ scanchain_114/module_data_in[5] scanchain_114/module_data_in[6] scanchain_114/module_data_in[7]
+ scanchain_114/module_data_out[0] scanchain_114/module_data_out[1] scanchain_114/module_data_out[2]
+ scanchain_114/module_data_out[3] scanchain_114/module_data_out[4] scanchain_114/module_data_out[5]
+ scanchain_114/module_data_out[6] scanchain_114/module_data_out[7] vccd1 vssd1 user_module_361728533238569985
Xuser_module_361728533238569985_136 scanchain_136/module_data_in[0] scanchain_136/module_data_in[1]
+ scanchain_136/module_data_in[2] scanchain_136/module_data_in[3] scanchain_136/module_data_in[4]
+ scanchain_136/module_data_in[5] scanchain_136/module_data_in[6] scanchain_136/module_data_in[7]
+ scanchain_136/module_data_out[0] scanchain_136/module_data_out[1] scanchain_136/module_data_out[2]
+ scanchain_136/module_data_out[3] scanchain_136/module_data_out[4] scanchain_136/module_data_out[5]
+ scanchain_136/module_data_out[6] scanchain_136/module_data_out[7] vccd1 vssd1 user_module_361728533238569985
Xuser_module_361728533238569985_103 scanchain_103/module_data_in[0] scanchain_103/module_data_in[1]
+ scanchain_103/module_data_in[2] scanchain_103/module_data_in[3] scanchain_103/module_data_in[4]
+ scanchain_103/module_data_in[5] scanchain_103/module_data_in[6] scanchain_103/module_data_in[7]
+ scanchain_103/module_data_out[0] scanchain_103/module_data_out[1] scanchain_103/module_data_out[2]
+ scanchain_103/module_data_out[3] scanchain_103/module_data_out[4] scanchain_103/module_data_out[5]
+ scanchain_103/module_data_out[6] scanchain_103/module_data_out[7] vccd1 vssd1 user_module_361728533238569985
Xuser_module_361728533238569985_147 scanchain_147/module_data_in[0] scanchain_147/module_data_in[1]
+ scanchain_147/module_data_in[2] scanchain_147/module_data_in[3] scanchain_147/module_data_in[4]
+ scanchain_147/module_data_in[5] scanchain_147/module_data_in[6] scanchain_147/module_data_in[7]
+ scanchain_147/module_data_out[0] scanchain_147/module_data_out[1] scanchain_147/module_data_out[2]
+ scanchain_147/module_data_out[3] scanchain_147/module_data_out[4] scanchain_147/module_data_out[5]
+ scanchain_147/module_data_out[6] scanchain_147/module_data_out[7] vccd1 vssd1 user_module_361728533238569985
Xscanchain_009 scanchain_009/clk_in scanchain_010/clk_in scanchain_009/data_in scanchain_010/data_in
+ scanchain_009/latch_enable_in scanchain_010/latch_enable_in scanchain_009/module_data_in[0]
+ scanchain_009/module_data_in[1] scanchain_009/module_data_in[2] scanchain_009/module_data_in[3]
+ scanchain_009/module_data_in[4] scanchain_009/module_data_in[5] scanchain_009/module_data_in[6]
+ scanchain_009/module_data_in[7] scanchain_009/module_data_out[0] scanchain_009/module_data_out[1]
+ scanchain_009/module_data_out[2] scanchain_009/module_data_out[3] scanchain_009/module_data_out[4]
+ scanchain_009/module_data_out[5] scanchain_009/module_data_out[6] scanchain_009/module_data_out[7]
+ scanchain_009/scan_select_in scanchain_010/scan_select_in vccd1 vssd1 scanchain
Xlucaz97_tt_top_073 lucaz97_tt_top_073/io_in[0] lucaz97_tt_top_073/io_in[1] lucaz97_tt_top_073/io_in[2]
+ lucaz97_tt_top_073/io_in[3] lucaz97_tt_top_073/io_in[4] lucaz97_tt_top_073/io_in[5]
+ lucaz97_tt_top_073/io_in[6] lucaz97_tt_top_073/io_in[7] lucaz97_tt_top_073/io_out[0]
+ lucaz97_tt_top_073/io_out[1] lucaz97_tt_top_073/io_out[2] lucaz97_tt_top_073/io_out[3]
+ lucaz97_tt_top_073/io_out[4] lucaz97_tt_top_073/io_out[5] lucaz97_tt_top_073/io_out[6]
+ lucaz97_tt_top_073/io_out[7] vccd1 vssd1 lucaz97_tt_top
Xuser_module_361728533238569985_169 scanchain_169/module_data_in[0] scanchain_169/module_data_in[1]
+ scanchain_169/module_data_in[2] scanchain_169/module_data_in[3] scanchain_169/module_data_in[4]
+ scanchain_169/module_data_in[5] scanchain_169/module_data_in[6] scanchain_169/module_data_in[7]
+ scanchain_169/module_data_out[0] scanchain_169/module_data_out[1] scanchain_169/module_data_out[2]
+ scanchain_169/module_data_out[3] scanchain_169/module_data_out[4] scanchain_169/module_data_out[5]
+ scanchain_169/module_data_out[6] scanchain_169/module_data_out[7] vccd1 vssd1 user_module_361728533238569985
Xuser_module_361728533238569985_158 scanchain_158/module_data_in[0] scanchain_158/module_data_in[1]
+ scanchain_158/module_data_in[2] scanchain_158/module_data_in[3] scanchain_158/module_data_in[4]
+ scanchain_158/module_data_in[5] scanchain_158/module_data_in[6] scanchain_158/module_data_in[7]
+ scanchain_158/module_data_out[0] scanchain_158/module_data_out[1] scanchain_158/module_data_out[2]
+ scanchain_158/module_data_out[3] scanchain_158/module_data_out[4] scanchain_158/module_data_out[5]
+ scanchain_158/module_data_out[6] scanchain_158/module_data_out[7] vccd1 vssd1 user_module_361728533238569985
Xyubex_tiny_logic_analyzer_031 scanchain_031/module_data_in[0] scanchain_031/module_data_in[1]
+ scanchain_031/module_data_in[2] scanchain_031/module_data_in[3] scanchain_031/module_data_in[4]
+ scanchain_031/module_data_in[5] scanchain_031/module_data_in[6] scanchain_031/module_data_in[7]
+ scanchain_031/module_data_out[0] scanchain_031/module_data_out[1] scanchain_031/module_data_out[2]
+ scanchain_031/module_data_out[3] scanchain_031/module_data_out[4] scanchain_031/module_data_out[5]
+ scanchain_031/module_data_out[6] scanchain_031/module_data_out[7] vccd1 vssd1 yubex_tiny_logic_analyzer
Xscanchain_181 scanchain_181/clk_in scanchain_182/clk_in scanchain_181/data_in scanchain_182/data_in
+ scanchain_181/latch_enable_in scanchain_182/latch_enable_in scanchain_181/module_data_in[0]
+ scanchain_181/module_data_in[1] scanchain_181/module_data_in[2] scanchain_181/module_data_in[3]
+ scanchain_181/module_data_in[4] scanchain_181/module_data_in[5] scanchain_181/module_data_in[6]
+ scanchain_181/module_data_in[7] scanchain_181/module_data_out[0] scanchain_181/module_data_out[1]
+ scanchain_181/module_data_out[2] scanchain_181/module_data_out[3] scanchain_181/module_data_out[4]
+ scanchain_181/module_data_out[5] scanchain_181/module_data_out[6] scanchain_181/module_data_out[7]
+ scanchain_181/scan_select_in scanchain_182/scan_select_in vccd1 vssd1 scanchain
Xscanchain_192 scanchain_192/clk_in scanchain_193/clk_in scanchain_192/data_in scanchain_193/data_in
+ scanchain_192/latch_enable_in scanchain_193/latch_enable_in scanchain_192/module_data_in[0]
+ scanchain_192/module_data_in[1] scanchain_192/module_data_in[2] scanchain_192/module_data_in[3]
+ scanchain_192/module_data_in[4] scanchain_192/module_data_in[5] scanchain_192/module_data_in[6]
+ scanchain_192/module_data_in[7] scanchain_192/module_data_out[0] scanchain_192/module_data_out[1]
+ scanchain_192/module_data_out[2] scanchain_192/module_data_out[3] scanchain_192/module_data_out[4]
+ scanchain_192/module_data_out[5] scanchain_192/module_data_out[6] scanchain_192/module_data_out[7]
+ scanchain_192/scan_select_in scanchain_193/scan_select_in vccd1 vssd1 scanchain
Xscanchain_170 scanchain_170/clk_in scanchain_171/clk_in scanchain_170/data_in scanchain_171/data_in
+ scanchain_170/latch_enable_in scanchain_171/latch_enable_in scanchain_170/module_data_in[0]
+ scanchain_170/module_data_in[1] scanchain_170/module_data_in[2] scanchain_170/module_data_in[3]
+ scanchain_170/module_data_in[4] scanchain_170/module_data_in[5] scanchain_170/module_data_in[6]
+ scanchain_170/module_data_in[7] scanchain_170/module_data_out[0] scanchain_170/module_data_out[1]
+ scanchain_170/module_data_out[2] scanchain_170/module_data_out[3] scanchain_170/module_data_out[4]
+ scanchain_170/module_data_out[5] scanchain_170/module_data_out[6] scanchain_170/module_data_out[7]
+ scanchain_170/scan_select_in scanchain_171/scan_select_in vccd1 vssd1 scanchain
Xuser_module_361728533238569985_126 scanchain_126/module_data_in[0] scanchain_126/module_data_in[1]
+ scanchain_126/module_data_in[2] scanchain_126/module_data_in[3] scanchain_126/module_data_in[4]
+ scanchain_126/module_data_in[5] scanchain_126/module_data_in[6] scanchain_126/module_data_in[7]
+ scanchain_126/module_data_out[0] scanchain_126/module_data_out[1] scanchain_126/module_data_out[2]
+ scanchain_126/module_data_out[3] scanchain_126/module_data_out[4] scanchain_126/module_data_out[5]
+ scanchain_126/module_data_out[6] scanchain_126/module_data_out[7] vccd1 vssd1 user_module_361728533238569985
Xuser_module_361728533238569985_115 scanchain_115/module_data_in[0] scanchain_115/module_data_in[1]
+ scanchain_115/module_data_in[2] scanchain_115/module_data_in[3] scanchain_115/module_data_in[4]
+ scanchain_115/module_data_in[5] scanchain_115/module_data_in[6] scanchain_115/module_data_in[7]
+ scanchain_115/module_data_out[0] scanchain_115/module_data_out[1] scanchain_115/module_data_out[2]
+ scanchain_115/module_data_out[3] scanchain_115/module_data_out[4] scanchain_115/module_data_out[5]
+ scanchain_115/module_data_out[6] scanchain_115/module_data_out[7] vccd1 vssd1 user_module_361728533238569985
Xuser_module_361728533238569985_137 scanchain_137/module_data_in[0] scanchain_137/module_data_in[1]
+ scanchain_137/module_data_in[2] scanchain_137/module_data_in[3] scanchain_137/module_data_in[4]
+ scanchain_137/module_data_in[5] scanchain_137/module_data_in[6] scanchain_137/module_data_in[7]
+ scanchain_137/module_data_out[0] scanchain_137/module_data_out[1] scanchain_137/module_data_out[2]
+ scanchain_137/module_data_out[3] scanchain_137/module_data_out[4] scanchain_137/module_data_out[5]
+ scanchain_137/module_data_out[6] scanchain_137/module_data_out[7] vccd1 vssd1 user_module_361728533238569985
Xuser_module_361728533238569985_104 scanchain_104/module_data_in[0] scanchain_104/module_data_in[1]
+ scanchain_104/module_data_in[2] scanchain_104/module_data_in[3] scanchain_104/module_data_in[4]
+ scanchain_104/module_data_in[5] scanchain_104/module_data_in[6] scanchain_104/module_data_in[7]
+ scanchain_104/module_data_out[0] scanchain_104/module_data_out[1] scanchain_104/module_data_out[2]
+ scanchain_104/module_data_out[3] scanchain_104/module_data_out[4] scanchain_104/module_data_out[5]
+ scanchain_104/module_data_out[6] scanchain_104/module_data_out[7] vccd1 vssd1 user_module_361728533238569985
Xuser_module_361728533238569985_148 scanchain_148/module_data_in[0] scanchain_148/module_data_in[1]
+ scanchain_148/module_data_in[2] scanchain_148/module_data_in[3] scanchain_148/module_data_in[4]
+ scanchain_148/module_data_in[5] scanchain_148/module_data_in[6] scanchain_148/module_data_in[7]
+ scanchain_148/module_data_out[0] scanchain_148/module_data_out[1] scanchain_148/module_data_out[2]
+ scanchain_148/module_data_out[3] scanchain_148/module_data_out[4] scanchain_148/module_data_out[5]
+ scanchain_148/module_data_out[6] scanchain_148/module_data_out[7] vccd1 vssd1 user_module_361728533238569985
Xuser_module_361728533238569985_159 scanchain_159/module_data_in[0] scanchain_159/module_data_in[1]
+ scanchain_159/module_data_in[2] scanchain_159/module_data_in[3] scanchain_159/module_data_in[4]
+ scanchain_159/module_data_in[5] scanchain_159/module_data_in[6] scanchain_159/module_data_in[7]
+ scanchain_159/module_data_out[0] scanchain_159/module_data_out[1] scanchain_159/module_data_out[2]
+ scanchain_159/module_data_out[3] scanchain_159/module_data_out[4] scanchain_159/module_data_out[5]
+ scanchain_159/module_data_out[6] scanchain_159/module_data_out[7] vccd1 vssd1 user_module_361728533238569985
Xuser_module_339501025136214612_057 scanchain_057/module_data_in[0] scanchain_057/module_data_in[1]
+ scanchain_057/module_data_in[2] scanchain_057/module_data_in[3] scanchain_057/module_data_in[4]
+ scanchain_057/module_data_in[5] scanchain_057/module_data_in[6] scanchain_057/module_data_in[7]
+ scanchain_057/module_data_out[0] scanchain_057/module_data_out[1] scanchain_057/module_data_out[2]
+ scanchain_057/module_data_out[3] scanchain_057/module_data_out[4] scanchain_057/module_data_out[5]
+ scanchain_057/module_data_out[6] scanchain_057/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xscanchain_182 scanchain_182/clk_in scanchain_183/clk_in scanchain_182/data_in scanchain_183/data_in
+ scanchain_182/latch_enable_in scanchain_183/latch_enable_in scanchain_182/module_data_in[0]
+ scanchain_182/module_data_in[1] scanchain_182/module_data_in[2] scanchain_182/module_data_in[3]
+ scanchain_182/module_data_in[4] scanchain_182/module_data_in[5] scanchain_182/module_data_in[6]
+ scanchain_182/module_data_in[7] scanchain_182/module_data_out[0] scanchain_182/module_data_out[1]
+ scanchain_182/module_data_out[2] scanchain_182/module_data_out[3] scanchain_182/module_data_out[4]
+ scanchain_182/module_data_out[5] scanchain_182/module_data_out[6] scanchain_182/module_data_out[7]
+ scanchain_182/scan_select_in scanchain_183/scan_select_in vccd1 vssd1 scanchain
Xscanchain_193 scanchain_193/clk_in scanchain_194/clk_in scanchain_193/data_in scanchain_194/data_in
+ scanchain_193/latch_enable_in scanchain_194/latch_enable_in scanchain_193/module_data_in[0]
+ scanchain_193/module_data_in[1] scanchain_193/module_data_in[2] scanchain_193/module_data_in[3]
+ scanchain_193/module_data_in[4] scanchain_193/module_data_in[5] scanchain_193/module_data_in[6]
+ scanchain_193/module_data_in[7] scanchain_193/module_data_out[0] scanchain_193/module_data_out[1]
+ scanchain_193/module_data_out[2] scanchain_193/module_data_out[3] scanchain_193/module_data_out[4]
+ scanchain_193/module_data_out[5] scanchain_193/module_data_out[6] scanchain_193/module_data_out[7]
+ scanchain_193/scan_select_in scanchain_194/scan_select_in vccd1 vssd1 scanchain
Xscanchain_171 scanchain_171/clk_in scanchain_172/clk_in scanchain_171/data_in scanchain_172/data_in
+ scanchain_171/latch_enable_in scanchain_172/latch_enable_in scanchain_171/module_data_in[0]
+ scanchain_171/module_data_in[1] scanchain_171/module_data_in[2] scanchain_171/module_data_in[3]
+ scanchain_171/module_data_in[4] scanchain_171/module_data_in[5] scanchain_171/module_data_in[6]
+ scanchain_171/module_data_in[7] scanchain_171/module_data_out[0] scanchain_171/module_data_out[1]
+ scanchain_171/module_data_out[2] scanchain_171/module_data_out[3] scanchain_171/module_data_out[4]
+ scanchain_171/module_data_out[5] scanchain_171/module_data_out[6] scanchain_171/module_data_out[7]
+ scanchain_171/scan_select_in scanchain_172/scan_select_in vccd1 vssd1 scanchain
Xscanchain_160 scanchain_160/clk_in scanchain_161/clk_in scanchain_160/data_in scanchain_161/data_in
+ scanchain_160/latch_enable_in scanchain_161/latch_enable_in scanchain_160/module_data_in[0]
+ scanchain_160/module_data_in[1] scanchain_160/module_data_in[2] scanchain_160/module_data_in[3]
+ scanchain_160/module_data_in[4] scanchain_160/module_data_in[5] scanchain_160/module_data_in[6]
+ scanchain_160/module_data_in[7] scanchain_160/module_data_out[0] scanchain_160/module_data_out[1]
+ scanchain_160/module_data_out[2] scanchain_160/module_data_out[3] scanchain_160/module_data_out[4]
+ scanchain_160/module_data_out[5] scanchain_160/module_data_out[6] scanchain_160/module_data_out[7]
+ scanchain_160/scan_select_in scanchain_161/scan_select_in vccd1 vssd1 scanchain
Xuser_module_361728533238569985_127 scanchain_127/module_data_in[0] scanchain_127/module_data_in[1]
+ scanchain_127/module_data_in[2] scanchain_127/module_data_in[3] scanchain_127/module_data_in[4]
+ scanchain_127/module_data_in[5] scanchain_127/module_data_in[6] scanchain_127/module_data_in[7]
+ scanchain_127/module_data_out[0] scanchain_127/module_data_out[1] scanchain_127/module_data_out[2]
+ scanchain_127/module_data_out[3] scanchain_127/module_data_out[4] scanchain_127/module_data_out[5]
+ scanchain_127/module_data_out[6] scanchain_127/module_data_out[7] vccd1 vssd1 user_module_361728533238569985
Xuser_module_361728533238569985_116 scanchain_116/module_data_in[0] scanchain_116/module_data_in[1]
+ scanchain_116/module_data_in[2] scanchain_116/module_data_in[3] scanchain_116/module_data_in[4]
+ scanchain_116/module_data_in[5] scanchain_116/module_data_in[6] scanchain_116/module_data_in[7]
+ scanchain_116/module_data_out[0] scanchain_116/module_data_out[1] scanchain_116/module_data_out[2]
+ scanchain_116/module_data_out[3] scanchain_116/module_data_out[4] scanchain_116/module_data_out[5]
+ scanchain_116/module_data_out[6] scanchain_116/module_data_out[7] vccd1 vssd1 user_module_361728533238569985
Xuser_module_361728533238569985_138 scanchain_138/module_data_in[0] scanchain_138/module_data_in[1]
+ scanchain_138/module_data_in[2] scanchain_138/module_data_in[3] scanchain_138/module_data_in[4]
+ scanchain_138/module_data_in[5] scanchain_138/module_data_in[6] scanchain_138/module_data_in[7]
+ scanchain_138/module_data_out[0] scanchain_138/module_data_out[1] scanchain_138/module_data_out[2]
+ scanchain_138/module_data_out[3] scanchain_138/module_data_out[4] scanchain_138/module_data_out[5]
+ scanchain_138/module_data_out[6] scanchain_138/module_data_out[7] vccd1 vssd1 user_module_361728533238569985
Xuser_module_361728533238569985_105 scanchain_105/module_data_in[0] scanchain_105/module_data_in[1]
+ scanchain_105/module_data_in[2] scanchain_105/module_data_in[3] scanchain_105/module_data_in[4]
+ scanchain_105/module_data_in[5] scanchain_105/module_data_in[6] scanchain_105/module_data_in[7]
+ scanchain_105/module_data_out[0] scanchain_105/module_data_out[1] scanchain_105/module_data_out[2]
+ scanchain_105/module_data_out[3] scanchain_105/module_data_out[4] scanchain_105/module_data_out[5]
+ scanchain_105/module_data_out[6] scanchain_105/module_data_out[7] vccd1 vssd1 user_module_361728533238569985
Xuser_module_361728533238569985_149 scanchain_149/module_data_in[0] scanchain_149/module_data_in[1]
+ scanchain_149/module_data_in[2] scanchain_149/module_data_in[3] scanchain_149/module_data_in[4]
+ scanchain_149/module_data_in[5] scanchain_149/module_data_in[6] scanchain_149/module_data_in[7]
+ scanchain_149/module_data_out[0] scanchain_149/module_data_out[1] scanchain_149/module_data_out[2]
+ scanchain_149/module_data_out[3] scanchain_149/module_data_out[4] scanchain_149/module_data_out[5]
+ scanchain_149/module_data_out[6] scanchain_149/module_data_out[7] vccd1 vssd1 user_module_361728533238569985
Xuser_module_347144898258928211_086 scanchain_086/module_data_in[0] scanchain_086/module_data_in[1]
+ scanchain_086/module_data_in[2] scanchain_086/module_data_in[3] scanchain_086/module_data_in[4]
+ scanchain_086/module_data_in[5] scanchain_086/module_data_in[6] scanchain_086/module_data_in[7]
+ scanchain_086/module_data_out[0] scanchain_086/module_data_out[1] scanchain_086/module_data_out[2]
+ scanchain_086/module_data_out[3] scanchain_086/module_data_out[4] scanchain_086/module_data_out[5]
+ scanchain_086/module_data_out[6] scanchain_086/module_data_out[7] vccd1 vssd1 user_module_347144898258928211
.ends

