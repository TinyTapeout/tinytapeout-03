

module meiniki_pi
(
  input  [7:0] io_in,
  output [7:0] io_out
);

wire       clk      = io_in[0];
wire       reset    = io_in[1];

reg  [11:0] index;
wire [3:0]  digit_tripple[0:2];
wire [3:0]  digit;
wire [3:0]  digit_out;
wire [1:0]  sel;
wire [9:0]  code;
reg         dot_done;

assign sel    = index[1:0];
assign digit  = digit_tripple[sel];
assign code   = f(index[11:2]);

assign digit_out = (index == 'b1) && ~dot_done ? 4'b1010 : digit;

always @(posedge clk) begin
  if (reset) begin
    index     <= 'b0;
    dot_done  <= 'b0;
  end else begin
    if (index[1:0] == 'b10) begin
      index <= index + 'd2;
    //end else if ((index[11:2] == 'd466) && (index[1:0] == 'b10)) begin
    //  index <= 'b0;
    end else begin
      if (dot_done | index != 'b1) begin
        index <= index + 'd1;
      end else begin
        dot_done <= 1'b1;
      end
    end
  end
end

decoder i_decoder (
  .code     ( digit_out ),
  .segments ( io_out    )
);

decode1000 i_dpd ( 
  .in_000 ( code[0]             ), 
  .in_001 ( code[1]             ), 
  .in_002 ( code[2]             ), 
  .in_003 ( code[3]             ), 
  .in_004 ( code[4]             ), 
  .in_005 ( code[5]             ), 
  .in_006 ( code[6]             ), 
  .in_007 ( code[7]             ), 
  .in_008 ( code[8]             ), 
  .in_009 ( code[9]             ), 
  .out000 ( digit_tripple[2][0] ),
  .out001 ( digit_tripple[2][1] ),
  .out002 ( digit_tripple[2][2] ),
  .out003 ( digit_tripple[2][3] ),
  .out004 ( digit_tripple[1][0] ),
  .out005 ( digit_tripple[1][1] ),
  .out006 ( digit_tripple[1][2] ),
  .out007 ( digit_tripple[1][3] ),
  .out008 ( digit_tripple[0][0] ),
  .out009 ( digit_tripple[0][1] ),
  .out010 ( digit_tripple[0][2] ),
  .out011 ( digit_tripple[0][3] )
);


function [9:0] f(input [9:0] index);
  case( index ) 
  0: f = 10'b0110010100;
  1: f = 10'b0011011001;
  2: f = 10'b0101100101;
  3: f = 10'b0111011000;
  4: f = 10'b1110111111;
  5: f = 10'b0110100011;
  6: f = 10'b1101001100;
  7: f = 10'b0101100100;
  8: f = 10'b0110111000;
  9: f = 10'b0110100111;
  10: f = 10'b0011011100;
  11: f = 10'b0101001110;
  12: f = 10'b1000011001;
  13: f = 10'b1110010110;
  14: f = 10'b0110111111;
  15: f = 10'b1110111101;
  16: f = 10'b1010010000;
  17: f = 10'b1010101010;
  18: f = 10'b0001111011;
  19: f = 10'b1001011010;
  20: f = 10'b1001011001;
  21: f = 10'b0100110000;
  22: f = 10'b1110001011;
  23: f = 10'b1101000000;
  24: f = 10'b1100101000;
  25: f = 10'b1100100000;
  26: f = 10'b1101111111;
  27: f = 10'b0101101100;
  28: f = 10'b0100001101;
  29: f = 10'b1000101010;
  30: f = 10'b1010110100;
  31: f = 10'b0100010001;
  32: f = 10'b1110000110;
  33: f = 10'b1111011110;
  34: f = 10'b0100010100;
  35: f = 10'b0000101110;
  36: f = 10'b1101010001;
  37: f = 10'b0110101000;
  38: f = 10'b0100110000;
  39: f = 10'b1101100100;
  40: f = 10'b1110001001;
  41: f = 10'b0111001010;
  42: f = 10'b1001100000;
  43: f = 10'b1011011101;
  44: f = 10'b0001011000;
  45: f = 10'b0100100011;
  46: f = 10'b0011110010;
  47: f = 10'b1010110101;
  48: f = 10'b0011001100;
  49: f = 10'b0100011100;
  50: f = 10'b1000101110;
  51: f = 10'b0010010001;
  52: f = 10'b1111000101;
  53: f = 10'b0000101000;
  54: f = 10'b1000010000;
  55: f = 10'b0101110000;
  56: f = 10'b0010111011;
  57: f = 10'b0101011100;
  58: f = 10'b0010010000;
  59: f = 10'b1011010101;
  60: f = 10'b1011101100;
  61: f = 10'b1001100010;
  62: f = 10'b0101011010;
  63: f = 10'b1000011111;
  64: f = 10'b1000111011;
  65: f = 10'b0000111000;
  66: f = 10'b0011111010;
  67: f = 10'b1001000010;
  68: f = 10'b0000001111;
  69: f = 10'b0001111011;
  70: f = 10'b1011100110;
  71: f = 10'b1010111011;
  72: f = 10'b0111000100;
  73: f = 10'b1100010010;
  74: f = 10'b1101001101;
  75: f = 10'b1011100100;
  76: f = 10'b0100101101;
  77: f = 10'b0111111000;
  78: f = 10'b1101111000;
  79: f = 10'b0110010110;
  80: f = 10'b1010100111;
  81: f = 10'b0010100000;
  82: f = 10'b0010011010;
  83: f = 10'b1010011100;
  84: f = 10'b1011100100;
  85: f = 10'b1101011100;
  86: f = 10'b1100111010;
  87: f = 10'b0111000110;
  88: f = 10'b0000110100;
  89: f = 10'b0001101101;
  90: f = 10'b0001000101;
  91: f = 10'b1000110010;
  92: f = 10'b1101100100;
  93: f = 10'b0000101101;
  94: f = 10'b0110111001;
  95: f = 10'b0111100000;
  96: f = 10'b1110100110;
  97: f = 10'b0000100100;
  98: f = 10'b1010011100;
  99: f = 10'b0010100111;
  100: f = 10'b0111110010;
  101: f = 10'b1001011000;
  102: f = 10'b1110000000;
  103: f = 10'b1101100000;
  104: f = 10'b1100110001;
  105: f = 10'b1011011000;
  106: f = 10'b1100011101;
  107: f = 10'b1001001110;
  108: f = 10'b0011010010;
  109: f = 10'b0000111010;
  110: f = 10'b0001111010;
  111: f = 10'b0100101010;
  112: f = 10'b1010101101;
  113: f = 10'b1000001001;
  114: f = 10'b0011110001;
  115: f = 10'b1010110110;
  116: f = 10'b1000110110;
  117: f = 10'b1111001111;
  118: f = 10'b0101011001;
  119: f = 10'b0000110110;
  120: f = 10'b0000000001;
  121: f = 10'b0010110011;
  122: f = 10'b0001010011;
  123: f = 10'b0001010100;
  124: f = 10'b0100001110;
  125: f = 10'b0001000110;
  126: f = 10'b1101010010;
  127: f = 10'b0010111000;
  128: f = 10'b1000010100;
  129: f = 10'b1101011011;
  130: f = 10'b0011011010;
  131: f = 10'b0011010001;
  132: f = 10'b0011100000;
  133: f = 10'b0111001101;
  134: f = 10'b0110000101;
  135: f = 10'b1110100111;
  136: f = 10'b0000110110;
  137: f = 10'b1011110101;
  138: f = 10'b1010111111;
  139: f = 10'b0011011011;
  140: f = 10'b0110001001;
  141: f = 10'b0100011000;
  142: f = 10'b1100010001;
  143: f = 10'b1110111000;
  144: f = 10'b0010111011;
  145: f = 10'b0101100001;
  146: f = 10'b0011111001;
  147: f = 10'b0110010000;
  148: f = 10'b1010010001;
  149: f = 10'b1001011100;
  150: f = 10'b1100001101;
  151: f = 10'b1001000110;
  152: f = 10'b0100110111;
  153: f = 10'b1110011110;
  154: f = 10'b0101110100;
  155: f = 10'b1111011100;
  156: f = 10'b1110110101;
  157: f = 10'b0011001110;
  158: f = 10'b1011110101;
  159: f = 10'b0101110010;
  160: f = 10'b1001001111;
  161: f = 10'b0010100010;
  162: f = 10'b1110111011;
  163: f = 10'b0000111110;
  164: f = 10'b0110000001;
  165: f = 10'b0011011010;
  166: f = 10'b0110011100;
  167: f = 10'b0110001111;
  168: f = 10'b0111100111;
  169: f = 10'b0110110110;
  170: f = 10'b0101000100;
  171: f = 10'b0001100101;
  172: f = 10'b1101100100;
  173: f = 10'b0110001000;
  174: f = 10'b1100000010;
  175: f = 10'b0010111001;
  176: f = 10'b1001011010;
  177: f = 10'b1100111001;
  178: f = 10'b1010100010;
  179: f = 10'b1001110011;
  180: f = 10'b1110011001;
  181: f = 10'b0001110000;
  182: f = 10'b0100010111;
  183: f = 10'b1110001110;
  184: f = 10'b0001011010;
  185: f = 10'b0111110000;
  186: f = 10'b0101110111;
  187: f = 10'b0001010011;
  188: f = 10'b0010101101;
  189: f = 10'b1110010111;
  190: f = 10'b1100101001;
  191: f = 10'b0110010111;
  192: f = 10'b1101110101;
  193: f = 10'b0100111000;
  194: f = 10'b1001100111;
  195: f = 10'b1000001011;
  196: f = 10'b1101001100;
  197: f = 10'b1111100110;
  198: f = 10'b0011001100;
  199: f = 10'b1010010011;
  200: f = 10'b0100000000;
  201: f = 10'b0001010110;
  202: f = 10'b0100011100;
  203: f = 10'b1110010100;
  204: f = 10'b1010100110;
  205: f = 10'b0111010110;
  206: f = 10'b0000101010;
  207: f = 10'b1111111000;
  208: f = 10'b1011110111;
  209: f = 10'b0010110100;
  210: f = 10'b0101110101;
  211: f = 10'b1111111000;
  212: f = 10'b0011101100;
  213: f = 10'b1110011101;
  214: f = 10'b0111100011;
  215: f = 10'b1110010111;
  216: f = 10'b0101111100;
  217: f = 10'b0011000110;
  218: f = 10'b1001001100;
  219: f = 10'b0000011010;
  220: f = 10'b0010100010;
  221: f = 10'b1001011011;
  222: f = 10'b0111000011;
  223: f = 10'b0000010100;
  224: f = 10'b1101010100;
  225: f = 10'b1010111110;
  226: f = 10'b1010110111;
  227: f = 10'b0010000101;
  228: f = 10'b0001111001;
  229: f = 10'b0100100111;
  230: f = 10'b1110101110;
  231: f = 10'b1010101101;
  232: f = 10'b0100011110;
  233: f = 10'b0111010100;
  234: f = 10'b0100000001;
  235: f = 10'b1010011111;
  236: f = 10'b1100010001;
  237: f = 10'b0100010010;
  238: f = 10'b0110001100;
  239: f = 10'b0011111010;
  240: f = 10'b0001101010;
  241: f = 10'b1000000011;
  242: f = 10'b1001000001;
  243: f = 10'b1000011101;
  244: f = 10'b0010001111;
  245: f = 10'b0111100010;
  246: f = 10'b1111111101;
  247: f = 10'b1001110111;
  248: f = 10'b0010110000;
  249: f = 10'b1110011110;
  250: f = 10'b0001010001;
  251: f = 10'b0001111100;
  252: f = 10'b1110100001;
  253: f = 10'b0010110100;
  254: f = 10'b1111111111;
  255: f = 10'b1111111111;
  256: f = 10'b1100111101;
  257: f = 10'b0101111011;
  258: f = 10'b1000001100;
  259: f = 10'b1010011111;
  260: f = 10'b0010000101;
  261: f = 10'b0111111101;
  262: f = 10'b0011110011;
  263: f = 10'b0100001011;
  264: f = 10'b1100001001;
  265: f = 10'b1100110001;
  266: f = 10'b1000111111;
  267: f = 10'b1010000010;
  268: f = 10'b1001000101;
  269: f = 10'b1011001101;
  270: f = 10'b1010110100;
  271: f = 10'b1100011010;
  272: f = 10'b0000111100;
  273: f = 10'b0101100100;
  274: f = 10'b0101010010;
  275: f = 10'b0100110000;
  276: f = 10'b1000101101;
  277: f = 10'b0110110100;
  278: f = 10'b1001101000;
  279: f = 10'b1010000011;
  280: f = 10'b1010100110;
  281: f = 10'b0010111011;
  282: f = 10'b0010011000;
  283: f = 10'b1100011101;
  284: f = 10'b0010000001;
  285: f = 10'b0000000000;
  286: f = 10'b0110010011;
  287: f = 10'b1110101011;
  288: f = 10'b1001111101;
  289: f = 10'b0101001110;
  290: f = 10'b1101011000;
  291: f = 10'b1111010011;
  292: f = 10'b0110100000;
  293: f = 10'b0100111110;
  294: f = 10'b0011000010;
  295: f = 10'b0001100001;
  296: f = 10'b1110010111;
  297: f = 10'b1111100110;
  298: f = 10'b1010011100;
  299: f = 10'b1110110000;
  300: f = 10'b0111011001;
  301: f = 10'b1000101101;
  302: f = 10'b0111001001;
  303: f = 10'b0001000010;
  304: f = 10'b1001111101;
  305: f = 10'b1011000110;
  306: f = 10'b0101111101;
  307: f = 10'b0010010101;
  308: f = 10'b1111011100;
  309: f = 10'b0101101010;
  310: f = 10'b0111001110;
  311: f = 10'b0100110101;
  312: f = 10'b0111111000;
  313: f = 10'b1111011001;
  314: f = 10'b0111110101;
  315: f = 10'b0011011011;
  316: f = 10'b1111111000;
  317: f = 10'b0011001011;
  318: f = 10'b1111111000;
  319: f = 10'b0001010011;
  320: f = 10'b0100010111;
  321: f = 10'b0010100010;
  322: f = 10'b1100001010;
  323: f = 10'b1101100001;
  324: f = 10'b0110000000;
  325: f = 10'b0010111010;
  326: f = 10'b1111101011;
  327: f = 10'b1101100001;
  328: f = 10'b0010011001;
  329: f = 10'b1010011010;
  330: f = 10'b0010101101;
  331: f = 10'b1101000010;
  332: f = 10'b0000011001;
  333: f = 10'b0100011111;
  334: f = 10'b0000101111;
  335: f = 10'b1010100101;
  336: f = 10'b1110100000;
  337: f = 10'b0010000110;
  338: f = 10'b1011001000;
  339: f = 10'b1011101010;
  340: f = 10'b0110100111;
  341: f = 10'b1100001110;
  342: f = 10'b1010111011;
  343: f = 10'b1100010101;
  344: f = 10'b0110111000;
  345: f = 10'b0010101010;
  346: f = 10'b1111111010;
  347: f = 10'b0100101101;
  348: f = 10'b0000110000;
  349: f = 10'b0011011011;
  350: f = 10'b0100000011;
  351: f = 10'b1010110000;
  352: f = 10'b0011001011;
  353: f = 10'b0101111010;
  354: f = 10'b1101111111;
  355: f = 10'b1011110111;
  356: f = 10'b0111100010;
  357: f = 10'b0101011001;
  358: f = 10'b0011001101;
  359: f = 10'b0111001111;
  360: f = 10'b0010100100;
  361: f = 10'b0111111100;
  362: f = 10'b0011110111;
  363: f = 10'b1010101000;
  364: f = 10'b0111000111;
  365: f = 10'b0110011101;
  366: f = 10'b0011010001;
  367: f = 10'b1011010111;
  368: f = 10'b1001001011;
  369: f = 10'b1110100100;
  370: f = 10'b0101000101;
  371: f = 10'b1000010101;
  372: f = 10'b0001101001;
  373: f = 10'b1011011011;
  374: f = 10'b0000101010;
  375: f = 10'b0111011101;
  376: f = 10'b0110010001;
  377: f = 10'b1101101010;
  378: f = 10'b0011110010;
  379: f = 10'b1111001011;
  380: f = 10'b1011001110;
  381: f = 10'b1110001101;
  382: f = 10'b1010001001;
  383: f = 10'b0100111110;
  384: f = 10'b0011110101;
  385: f = 10'b1001100011;
  386: f = 10'b1111000110;
  387: f = 10'b1000111011;
  388: f = 10'b0010111101;
  389: f = 10'b1010101101;
  390: f = 10'b1010000110;
  391: f = 10'b0001000000;
  392: f = 10'b0000111010;
  393: f = 10'b1111110000;
  394: f = 10'b0011100111;
  395: f = 10'b0010010011;
  396: f = 10'b0010001100;
  397: f = 10'b1010001110;
  398: f = 10'b0100001110;
  399: f = 10'b1000000001;
  400: f = 10'b0101001011;
  401: f = 10'b1100111100;
  402: f = 10'b0011100000;
  403: f = 10'b0111010110;
  404: f = 10'b0111110000;
  405: f = 10'b1111100110;
  406: f = 10'b0000010000;
  407: f = 10'b1001110001;
  408: f = 10'b0000011000;
  409: f = 10'b0011011010;
  410: f = 10'b0101011011;
  411: f = 10'b1011011001;
  412: f = 10'b1100011001;
  413: f = 10'b1000011110;
  414: f = 10'b1101110110;
  415: f = 10'b1110101011;
  416: f = 10'b1111000100;
  417: f = 10'b1011001100;
  418: f = 10'b1000101101;
  419: f = 10'b1010110111;
  420: f = 10'b1111111101;
  421: f = 10'b1001110010;
  422: f = 10'b1101001010;
  423: f = 10'b1110010000;
  424: f = 10'b1000000100;
  425: f = 10'b1111010011;
  426: f = 10'b1001100100;
  427: f = 10'b1100100000;
  428: f = 10'b1000001100;
  429: f = 10'b1101101000;
  430: f = 10'b1000100101;
  431: f = 10'b1110001100;
  432: f = 10'b1010101111;
  433: f = 10'b0010101001;
  434: f = 10'b0110110001;
  435: f = 10'b0111100111;
  436: f = 10'b1110000010;
  437: f = 10'b1101111110;
  438: f = 10'b1010011101;
  439: f = 10'b0100010000;
  440: f = 10'b1001110101;
  441: f = 10'b0100010110;
  442: f = 10'b0100000101;
  443: f = 10'b1101111010;
  444: f = 10'b1100000010;
  445: f = 10'b1000000101;
  446: f = 10'b0100001101;
  447: f = 10'b1000011101;
  448: f = 10'b0000011001;
  449: f = 10'b0111010001;
  450: f = 10'b0010100101;
  451: f = 10'b0110111000;
  452: f = 10'b0101000011;
  453: f = 10'b0000000011;
  454: f = 10'b1011011000;
  455: f = 10'b1111100100;
  456: f = 10'b0000100100;
  457: f = 10'b1111001001;
  458: f = 10'b1101000111;
  459: f = 10'b0110100110;
  460: f = 10'b0110011011;
  461: f = 10'b1000011001;
  462: f = 10'b1110101101;
  463: f = 10'b0101100000;
  464: f = 10'b1000100110;
  465: f = 10'b0110011110;
  466: f = 10'b0101111001;
  default: f = 10'bXXXXXXXXXX;
  endcase
endfunction


endmodule
