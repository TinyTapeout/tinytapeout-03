VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO MichaelBell_hovalaag
  CLASS BLOCK ;
  FOREIGN MichaelBell_hovalaag ;
  ORIGIN 0.000 0.000 ;
  SIZE 150.000 BY 170.000 ;
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 8.200 2.000 8.800 ;
    END
  END io_in[0]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 18.400 2.000 19.000 ;
    END
  END io_in[1]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 28.600 2.000 29.200 ;
    END
  END io_in[2]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 38.800 2.000 39.400 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 49.000 2.000 49.600 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 59.200 2.000 59.800 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 69.400 2.000 70.000 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 79.600 2.000 80.200 ;
    END
  END io_in[7]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 89.800 2.000 90.400 ;
    END
  END io_out[0]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 100.000 2.000 100.600 ;
    END
  END io_out[1]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 110.200 2.000 110.800 ;
    END
  END io_out[2]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 120.400 2.000 121.000 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 130.600 2.000 131.200 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 140.800 2.000 141.400 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 151.000 2.000 151.600 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 161.200 2.000 161.800 ;
    END
  END io_out[7]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 22.085 5.200 23.685 163.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 56.815 5.200 58.415 163.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 91.545 5.200 93.145 163.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 126.275 5.200 127.875 163.440 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 39.450 5.200 41.050 163.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 74.180 5.200 75.780 163.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 108.910 5.200 110.510 163.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 143.640 5.200 145.240 163.440 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 5.355 144.440 163.285 ;
      LAYER met1 ;
        RECT 2.370 0.720 149.890 168.600 ;
      LAYER met2 ;
        RECT 2.390 0.690 149.860 168.630 ;
      LAYER met3 ;
        RECT 2.000 162.200 145.755 163.365 ;
        RECT 2.400 160.800 145.755 162.200 ;
        RECT 2.000 152.000 145.755 160.800 ;
        RECT 2.400 150.600 145.755 152.000 ;
        RECT 2.000 141.800 145.755 150.600 ;
        RECT 2.400 140.400 145.755 141.800 ;
        RECT 2.000 131.600 145.755 140.400 ;
        RECT 2.400 130.200 145.755 131.600 ;
        RECT 2.000 121.400 145.755 130.200 ;
        RECT 2.400 120.000 145.755 121.400 ;
        RECT 2.000 111.200 145.755 120.000 ;
        RECT 2.400 109.800 145.755 111.200 ;
        RECT 2.000 101.000 145.755 109.800 ;
        RECT 2.400 99.600 145.755 101.000 ;
        RECT 2.000 90.800 145.755 99.600 ;
        RECT 2.400 89.400 145.755 90.800 ;
        RECT 2.000 80.600 145.755 89.400 ;
        RECT 2.400 79.200 145.755 80.600 ;
        RECT 2.000 70.400 145.755 79.200 ;
        RECT 2.400 69.000 145.755 70.400 ;
        RECT 2.000 60.200 145.755 69.000 ;
        RECT 2.400 58.800 145.755 60.200 ;
        RECT 2.000 50.000 145.755 58.800 ;
        RECT 2.400 48.600 145.755 50.000 ;
        RECT 2.000 39.800 145.755 48.600 ;
        RECT 2.400 38.400 145.755 39.800 ;
        RECT 2.000 29.600 145.755 38.400 ;
        RECT 2.400 28.200 145.755 29.600 ;
        RECT 2.000 19.400 145.755 28.200 ;
        RECT 2.400 18.000 145.755 19.400 ;
        RECT 2.000 9.200 145.755 18.000 ;
        RECT 2.400 7.800 145.755 9.200 ;
        RECT 2.000 0.855 145.755 7.800 ;
      LAYER met4 ;
        RECT 7.655 5.615 21.685 159.625 ;
        RECT 24.085 5.615 39.050 159.625 ;
        RECT 41.450 5.615 56.415 159.625 ;
        RECT 58.815 5.615 73.780 159.625 ;
        RECT 76.180 5.615 91.145 159.625 ;
        RECT 93.545 5.615 108.510 159.625 ;
        RECT 110.910 5.615 125.875 159.625 ;
        RECT 128.275 5.615 142.305 159.625 ;
  END
END MichaelBell_hovalaag
END LIBRARY

