magic
tech sky130A
magscale 1 2
timestamp 1678955295
<< metal1 >>
rect 31662 700816 31668 700868
rect 31720 700856 31726 700868
rect 105446 700856 105452 700868
rect 31720 700828 105452 700856
rect 31720 700816 31726 700828
rect 105446 700816 105452 700828
rect 105504 700816 105510 700868
rect 62022 700748 62028 700800
rect 62080 700788 62086 700800
rect 202782 700788 202788 700800
rect 62080 700760 202788 700788
rect 62080 700748 62086 700760
rect 202782 700748 202788 700760
rect 202840 700748 202846 700800
rect 71038 700680 71044 700732
rect 71096 700720 71102 700732
rect 267642 700720 267648 700732
rect 71096 700692 267648 700720
rect 71096 700680 71102 700692
rect 267642 700680 267648 700692
rect 267700 700680 267706 700732
rect 23382 700612 23388 700664
rect 23440 700652 23446 700664
rect 235166 700652 235172 700664
rect 23440 700624 235172 700652
rect 23440 700612 23446 700624
rect 235166 700612 235172 700624
rect 235224 700612 235230 700664
rect 64782 700544 64788 700596
rect 64840 700584 64846 700596
rect 332502 700584 332508 700596
rect 64840 700556 332508 700584
rect 64840 700544 64846 700556
rect 332502 700544 332508 700556
rect 332560 700544 332566 700596
rect 17862 700476 17868 700528
rect 17920 700516 17926 700528
rect 300118 700516 300124 700528
rect 17920 700488 300124 700516
rect 17920 700476 17926 700488
rect 300118 700476 300124 700488
rect 300176 700476 300182 700528
rect 68278 700408 68284 700460
rect 68336 700448 68342 700460
rect 364978 700448 364984 700460
rect 68336 700420 364984 700448
rect 68336 700408 68342 700420
rect 364978 700408 364984 700420
rect 365036 700408 365042 700460
rect 28902 700340 28908 700392
rect 28960 700380 28966 700392
rect 462314 700380 462320 700392
rect 28960 700352 462320 700380
rect 28960 700340 28966 700352
rect 462314 700340 462320 700352
rect 462372 700340 462378 700392
rect 50982 700272 50988 700324
rect 51040 700312 51046 700324
rect 494790 700312 494796 700324
rect 51040 700284 494796 700312
rect 51040 700272 51046 700284
rect 494790 700272 494796 700284
rect 494848 700272 494854 700324
rect 57882 696940 57888 696992
rect 57940 696980 57946 696992
rect 580166 696980 580172 696992
rect 57940 696952 580172 696980
rect 57940 696940 57946 696952
rect 580166 696940 580172 696952
rect 580224 696940 580230 696992
rect 3510 656888 3516 656940
rect 3568 656928 3574 656940
rect 19978 656928 19984 656940
rect 3568 656900 19984 656928
rect 3568 656888 3574 656900
rect 19978 656888 19984 656900
rect 20036 656888 20042 656940
rect 3510 632068 3516 632120
rect 3568 632108 3574 632120
rect 18598 632108 18604 632120
rect 3568 632080 18604 632108
rect 3568 632068 3574 632080
rect 18598 632068 18604 632080
rect 18656 632068 18662 632120
rect 68370 590656 68376 590708
rect 68428 590696 68434 590708
rect 580166 590696 580172 590708
rect 68428 590668 580172 590696
rect 68428 590656 68434 590668
rect 580166 590656 580172 590668
rect 580224 590656 580230 590708
rect 22002 563048 22008 563100
rect 22060 563088 22066 563100
rect 580166 563088 580172 563100
rect 22060 563060 580172 563088
rect 22060 563048 22066 563060
rect 580166 563048 580172 563060
rect 580224 563048 580230 563100
rect 3326 553392 3332 553444
rect 3384 553432 3390 553444
rect 24118 553432 24124 553444
rect 3384 553404 24124 553432
rect 3384 553392 3390 553404
rect 24118 553392 24124 553404
rect 24176 553392 24182 553444
rect 68462 536800 68468 536852
rect 68520 536840 68526 536852
rect 580166 536840 580172 536852
rect 68520 536812 580172 536840
rect 68520 536800 68526 536812
rect 580166 536800 580172 536812
rect 580224 536800 580230 536852
rect 2774 527144 2780 527196
rect 2832 527184 2838 527196
rect 6178 527184 6184 527196
rect 2832 527156 6184 527184
rect 2832 527144 2838 527156
rect 6178 527144 6184 527156
rect 6236 527144 6242 527196
rect 30282 510620 30288 510672
rect 30340 510660 30346 510672
rect 580166 510660 580172 510672
rect 30340 510632 580172 510660
rect 30340 510620 30346 510632
rect 580166 510620 580172 510632
rect 580224 510620 580230 510672
rect 68554 470568 68560 470620
rect 68612 470608 68618 470620
rect 579982 470608 579988 470620
rect 68612 470580 579988 470608
rect 68612 470568 68618 470580
rect 579982 470568 579988 470580
rect 580040 470568 580046 470620
rect 3142 448536 3148 448588
rect 3200 448576 3206 448588
rect 43438 448576 43444 448588
rect 3200 448548 43444 448576
rect 3200 448536 3206 448548
rect 43438 448536 43444 448548
rect 43496 448536 43502 448588
rect 17770 430584 17776 430636
rect 17828 430624 17834 430636
rect 579614 430624 579620 430636
rect 17828 430596 579620 430624
rect 17828 430584 17834 430596
rect 579614 430584 579620 430596
rect 579672 430584 579678 430636
rect 17678 404336 17684 404388
rect 17736 404376 17742 404388
rect 580166 404376 580172 404388
rect 17736 404348 580172 404376
rect 17736 404336 17742 404348
rect 580166 404336 580172 404348
rect 580224 404336 580230 404388
rect 68646 378156 68652 378208
rect 68704 378196 68710 378208
rect 580166 378196 580172 378208
rect 68704 378168 580172 378196
rect 68704 378156 68710 378168
rect 580166 378156 580172 378168
rect 580224 378156 580230 378208
rect 3326 357416 3332 357468
rect 3384 357456 3390 357468
rect 65334 357456 65340 357468
rect 3384 357428 65340 357456
rect 3384 357416 3390 357428
rect 65334 357416 65340 357428
rect 65392 357416 65398 357468
rect 3326 345040 3332 345092
rect 3384 345080 3390 345092
rect 13078 345080 13084 345092
rect 3384 345052 13084 345080
rect 3384 345040 3390 345052
rect 13078 345040 13084 345052
rect 13136 345040 13142 345092
rect 3326 292544 3332 292596
rect 3384 292584 3390 292596
rect 14458 292584 14464 292596
rect 3384 292556 14464 292584
rect 3384 292544 3390 292556
rect 14458 292544 14464 292556
rect 14516 292544 14522 292596
rect 3326 253920 3332 253972
rect 3384 253960 3390 253972
rect 33778 253960 33784 253972
rect 3384 253932 33784 253960
rect 3384 253920 3390 253932
rect 33778 253920 33784 253932
rect 33836 253920 33842 253972
rect 39942 231820 39948 231872
rect 40000 231860 40006 231872
rect 579798 231860 579804 231872
rect 40000 231832 579804 231860
rect 40000 231820 40006 231832
rect 579798 231820 579804 231832
rect 579856 231820 579862 231872
rect 3326 201492 3332 201544
rect 3384 201532 3390 201544
rect 65242 201532 65248 201544
rect 3384 201504 65248 201532
rect 3384 201492 3390 201504
rect 65242 201492 65248 201504
rect 65300 201492 65306 201544
rect 66162 191836 66168 191888
rect 66220 191876 66226 191888
rect 580166 191876 580172 191888
rect 66220 191848 580172 191876
rect 66220 191836 66226 191848
rect 580166 191836 580172 191848
rect 580224 191836 580230 191888
rect 56502 151784 56508 151836
rect 56560 151824 56566 151836
rect 579982 151824 579988 151836
rect 56560 151796 579988 151824
rect 56560 151784 56566 151796
rect 579982 151784 579988 151796
rect 580040 151784 580046 151836
rect 3326 136620 3332 136672
rect 3384 136660 3390 136672
rect 15838 136660 15844 136672
rect 3384 136632 15844 136660
rect 3384 136620 3390 136632
rect 15838 136620 15844 136632
rect 15896 136620 15902 136672
rect 36630 52572 36636 52624
rect 36688 52612 36694 52624
rect 249058 52612 249064 52624
rect 36688 52584 249064 52612
rect 36688 52572 36694 52584
rect 249058 52572 249064 52584
rect 249116 52572 249122 52624
rect 17586 52504 17592 52556
rect 17644 52544 17650 52556
rect 249150 52544 249156 52556
rect 17644 52516 249156 52544
rect 17644 52504 17650 52516
rect 249150 52504 249156 52516
rect 249208 52504 249214 52556
rect 33042 52436 33048 52488
rect 33100 52476 33106 52488
rect 287698 52476 287704 52488
rect 33100 52448 287704 52476
rect 33100 52436 33106 52448
rect 287698 52436 287704 52448
rect 287756 52436 287762 52488
rect 176562 51076 176568 51128
rect 176620 51116 176626 51128
rect 178126 51116 178132 51128
rect 176620 51088 178132 51116
rect 176620 51076 176626 51088
rect 178126 51076 178132 51088
rect 178184 51076 178190 51128
rect 216582 51076 216588 51128
rect 216640 51116 216646 51128
rect 218054 51116 218060 51128
rect 216640 51088 218060 51116
rect 216640 51076 216646 51088
rect 218054 51076 218060 51088
rect 218112 51076 218118 51128
rect 96522 48288 96528 48340
rect 96580 48328 96586 48340
rect 97442 48328 97448 48340
rect 96580 48300 97448 48328
rect 96580 48288 96586 48300
rect 97442 48288 97448 48300
rect 97500 48288 97506 48340
rect 176470 48288 176476 48340
rect 176528 48328 176534 48340
rect 178126 48328 178132 48340
rect 176528 48300 178132 48328
rect 176528 48288 176534 48300
rect 178126 48288 178132 48300
rect 178184 48288 178190 48340
rect 217318 48288 217324 48340
rect 217376 48328 217382 48340
rect 218054 48328 218060 48340
rect 217376 48300 218060 48328
rect 217376 48288 217382 48300
rect 218054 48288 218060 48300
rect 218112 48288 218118 48340
rect 96246 46928 96252 46980
rect 96304 46968 96310 46980
rect 97442 46968 97448 46980
rect 96304 46940 97448 46968
rect 96304 46928 96310 46940
rect 97442 46928 97448 46940
rect 97500 46928 97506 46980
rect 216490 46928 216496 46980
rect 216548 46968 216554 46980
rect 218054 46968 218060 46980
rect 216548 46940 218060 46968
rect 216548 46928 216554 46940
rect 218054 46928 218060 46940
rect 218112 46928 218118 46980
rect 257338 46928 257344 46980
rect 257396 46968 257402 46980
rect 258258 46968 258264 46980
rect 257396 46940 258264 46968
rect 257396 46928 257402 46940
rect 258258 46928 258264 46940
rect 258316 46928 258322 46980
rect 3418 46180 3424 46232
rect 3476 46220 3482 46232
rect 58618 46220 58624 46232
rect 3476 46192 58624 46220
rect 3476 46180 3482 46192
rect 58618 46180 58624 46192
rect 58676 46180 58682 46232
rect 3418 46044 3424 46096
rect 3476 46084 3482 46096
rect 3786 46084 3792 46096
rect 3476 46056 3792 46084
rect 3476 46044 3482 46056
rect 3786 46044 3792 46056
rect 3844 46044 3850 46096
rect 2958 44140 2964 44192
rect 3016 44180 3022 44192
rect 16482 44180 16488 44192
rect 3016 44152 16488 44180
rect 3016 44140 3022 44152
rect 16482 44140 16488 44152
rect 16540 44140 16546 44192
rect 96338 44140 96344 44192
rect 96396 44180 96402 44192
rect 97442 44180 97448 44192
rect 96396 44152 97448 44180
rect 96396 44140 96402 44152
rect 97442 44140 97448 44152
rect 97500 44140 97506 44192
rect 257246 44140 257252 44192
rect 257304 44180 257310 44192
rect 258258 44180 258264 44192
rect 257304 44152 258264 44180
rect 257304 44140 257310 44152
rect 258258 44140 258264 44152
rect 258316 44140 258322 44192
rect 216398 43052 216404 43104
rect 216456 43092 216462 43104
rect 217962 43092 217968 43104
rect 216456 43064 217968 43092
rect 216456 43052 216462 43064
rect 217962 43052 217968 43064
rect 218020 43052 218026 43104
rect 176286 42780 176292 42832
rect 176344 42820 176350 42832
rect 178126 42820 178132 42832
rect 176344 42792 178132 42820
rect 176344 42780 176350 42792
rect 178126 42780 178132 42792
rect 178184 42780 178190 42832
rect 19978 42712 19984 42764
rect 20036 42752 20042 42764
rect 26418 42752 26424 42764
rect 20036 42724 26424 42752
rect 20036 42712 20042 42724
rect 26418 42712 26424 42724
rect 26476 42712 26482 42764
rect 33778 42712 33784 42764
rect 33836 42752 33842 42764
rect 37366 42752 37372 42764
rect 33836 42724 37372 42752
rect 33836 42712 33842 42724
rect 37366 42712 37372 42724
rect 37424 42712 37430 42764
rect 43438 42712 43444 42764
rect 43496 42752 43502 42764
rect 45738 42752 45744 42764
rect 43496 42724 45744 42752
rect 43496 42712 43502 42724
rect 45738 42712 45744 42724
rect 45796 42712 45802 42764
rect 257154 42644 257160 42696
rect 257212 42684 257218 42696
rect 258166 42684 258172 42696
rect 257212 42656 258172 42684
rect 257212 42644 257218 42656
rect 258166 42644 258172 42656
rect 258224 42644 258230 42696
rect 18598 42372 18604 42424
rect 18656 42412 18662 42424
rect 24486 42412 24492 42424
rect 18656 42384 24492 42412
rect 18656 42372 18662 42384
rect 24486 42372 24492 42384
rect 24544 42372 24550 42424
rect 65150 42372 65156 42424
rect 65208 42412 65214 42424
rect 66162 42412 66168 42424
rect 65208 42384 66168 42412
rect 65208 42372 65214 42384
rect 66162 42372 66168 42384
rect 66220 42372 66226 42424
rect 24118 42168 24124 42220
rect 24176 42208 24182 42220
rect 34146 42208 34152 42220
rect 24176 42180 34152 42208
rect 24176 42168 24182 42180
rect 34146 42168 34152 42180
rect 34204 42168 34210 42220
rect 40494 42168 40500 42220
rect 40552 42208 40558 42220
rect 52178 42208 52184 42220
rect 40552 42180 52184 42208
rect 40552 42168 40558 42180
rect 52178 42168 52184 42180
rect 52236 42168 52242 42220
rect 3418 42100 3424 42152
rect 3476 42140 3482 42152
rect 42518 42140 42524 42152
rect 3476 42112 42524 42140
rect 3476 42100 3482 42112
rect 42518 42100 42524 42112
rect 42576 42100 42582 42152
rect 3786 42032 3792 42084
rect 3844 42072 3850 42084
rect 48958 42072 48964 42084
rect 3844 42044 48964 42072
rect 3844 42032 3850 42044
rect 48958 42032 48964 42044
rect 49016 42032 49022 42084
rect 91002 41964 91008 42016
rect 91060 42004 91066 42016
rect 95878 42004 95884 42016
rect 91060 41976 95884 42004
rect 91060 41964 91066 41976
rect 95878 41964 95884 41976
rect 95936 41964 95942 42016
rect 131022 41964 131028 42016
rect 131080 42004 131086 42016
rect 135898 42004 135904 42016
rect 131080 41976 135904 42004
rect 131080 41964 131086 41976
rect 135898 41964 135904 41976
rect 135956 41964 135962 42016
rect 171410 41964 171416 42016
rect 171468 42004 171474 42016
rect 175918 42004 175924 42016
rect 171468 41976 175924 42004
rect 171468 41964 171474 41976
rect 175918 41964 175924 41976
rect 175976 41964 175982 42016
rect 40678 41420 40684 41472
rect 40736 41460 40742 41472
rect 65518 41460 65524 41472
rect 40736 41432 65524 41460
rect 40736 41420 40742 41432
rect 65518 41420 65524 41432
rect 65576 41420 65582 41472
rect 366358 40672 366364 40724
rect 366416 40712 366422 40724
rect 580902 40712 580908 40724
rect 366416 40684 580908 40712
rect 366416 40672 366422 40684
rect 580902 40672 580908 40684
rect 580960 40672 580966 40724
rect 176378 40060 176384 40112
rect 176436 40100 176442 40112
rect 178126 40100 178132 40112
rect 176436 40072 178132 40100
rect 176436 40060 176442 40072
rect 178126 40060 178132 40072
rect 178184 40060 178190 40112
rect 17678 39992 17684 40044
rect 17736 40032 17742 40044
rect 19702 40032 19708 40044
rect 17736 40004 19708 40032
rect 17736 39992 17742 40004
rect 19702 39992 19708 40004
rect 19760 39992 19766 40044
rect 176562 39380 176568 39432
rect 176620 39420 176626 39432
rect 178034 39420 178040 39432
rect 176620 39392 178040 39420
rect 176620 39380 176626 39392
rect 178034 39380 178040 39392
rect 178092 39380 178098 39432
rect 176470 38632 176476 38684
rect 176528 38672 176534 38684
rect 178126 38672 178132 38684
rect 176528 38644 178132 38672
rect 176528 38632 176534 38644
rect 178126 38632 178132 38644
rect 178184 38632 178190 38684
rect 176746 37884 176752 37936
rect 176804 37924 176810 37936
rect 177850 37924 177856 37936
rect 176804 37896 177856 37924
rect 176804 37884 176810 37896
rect 177850 37884 177856 37896
rect 177908 37884 177914 37936
rect 216582 37884 216588 37936
rect 216640 37924 216646 37936
rect 218054 37924 218060 37936
rect 216640 37896 218060 37924
rect 216640 37884 216646 37896
rect 218054 37884 218060 37896
rect 218112 37884 218118 37936
rect 96338 37136 96344 37188
rect 96396 37176 96402 37188
rect 97442 37176 97448 37188
rect 96396 37148 97448 37176
rect 96396 37136 96402 37148
rect 97442 37136 97448 37148
rect 97500 37136 97506 37188
rect 257338 35912 257344 35964
rect 257396 35952 257402 35964
rect 258258 35952 258264 35964
rect 257396 35924 258264 35952
rect 257396 35912 257402 35924
rect 258258 35912 258264 35924
rect 258316 35912 258322 35964
rect 3234 35844 3240 35896
rect 3292 35884 3298 35896
rect 17862 35884 17868 35896
rect 3292 35856 17868 35884
rect 3292 35844 3298 35856
rect 17862 35844 17868 35856
rect 17920 35844 17926 35896
rect 176746 34484 176752 34536
rect 176804 34524 176810 34536
rect 177850 34524 177856 34536
rect 176804 34496 177856 34524
rect 176804 34484 176810 34496
rect 177850 34484 177856 34496
rect 177908 34484 177914 34536
rect 216858 34484 216864 34536
rect 216916 34524 216922 34536
rect 217962 34524 217968 34536
rect 216916 34496 217968 34524
rect 216916 34484 216922 34496
rect 217962 34484 217968 34496
rect 218020 34484 218026 34536
rect 257154 34484 257160 34536
rect 257212 34524 257218 34536
rect 258258 34524 258264 34536
rect 257212 34496 258264 34524
rect 257212 34484 257218 34496
rect 258258 34484 258264 34496
rect 258316 34484 258322 34536
rect 287698 33056 287704 33108
rect 287756 33096 287762 33108
rect 580166 33096 580172 33108
rect 287756 33068 580172 33096
rect 287756 33056 287762 33068
rect 580166 33056 580172 33068
rect 580224 33056 580230 33108
rect 96338 32920 96344 32972
rect 96396 32960 96402 32972
rect 97442 32960 97448 32972
rect 96396 32932 97448 32960
rect 96396 32920 96402 32932
rect 97442 32920 97448 32932
rect 97500 32920 97506 32972
rect 216490 32852 216496 32904
rect 216548 32892 216554 32904
rect 217962 32892 217968 32904
rect 216548 32864 217968 32892
rect 216548 32852 216554 32864
rect 217962 32852 217968 32864
rect 218020 32852 218026 32904
rect 176562 31900 176568 31952
rect 176620 31940 176626 31952
rect 178126 31940 178132 31952
rect 176620 31912 178132 31940
rect 176620 31900 176626 31912
rect 178126 31900 178132 31912
rect 178184 31900 178190 31952
rect 216582 31900 216588 31952
rect 216640 31940 216646 31952
rect 218054 31940 218060 31952
rect 216640 31912 218060 31940
rect 216640 31900 216646 31912
rect 218054 31900 218060 31912
rect 218112 31900 218118 31952
rect 67726 31424 67732 31476
rect 67784 31464 67790 31476
rect 71038 31464 71044 31476
rect 67784 31436 71044 31464
rect 67784 31424 67790 31436
rect 71038 31424 71044 31436
rect 71096 31424 71102 31476
rect 96338 28908 96344 28960
rect 96396 28948 96402 28960
rect 97534 28948 97540 28960
rect 96396 28920 97540 28948
rect 96396 28908 96402 28920
rect 97534 28908 97540 28920
rect 97592 28908 97598 28960
rect 176562 28908 176568 28960
rect 176620 28948 176626 28960
rect 178034 28948 178040 28960
rect 176620 28920 178040 28948
rect 176620 28908 176626 28920
rect 178034 28908 178040 28920
rect 178092 28908 178098 28960
rect 96522 27616 96528 27668
rect 96580 27656 96586 27668
rect 97442 27656 97448 27668
rect 96580 27628 97448 27656
rect 96580 27616 96586 27628
rect 97442 27616 97448 27628
rect 97500 27616 97506 27668
rect 176746 27616 176752 27668
rect 176804 27656 176810 27668
rect 177850 27656 177856 27668
rect 176804 27628 177856 27656
rect 176804 27616 176810 27628
rect 177850 27616 177856 27628
rect 177908 27616 177914 27668
rect 257338 27616 257344 27668
rect 257396 27656 257402 27668
rect 258258 27656 258264 27668
rect 257396 27628 258264 27656
rect 257396 27616 257402 27628
rect 258258 27616 258264 27628
rect 258316 27616 258322 27668
rect 13078 27548 13084 27600
rect 13136 27588 13142 27600
rect 17862 27588 17868 27600
rect 13136 27560 17868 27588
rect 13136 27548 13142 27560
rect 17862 27548 17868 27560
rect 17920 27548 17926 27600
rect 96338 27412 96344 27464
rect 96396 27452 96402 27464
rect 97350 27452 97356 27464
rect 96396 27424 97356 27452
rect 96396 27412 96402 27424
rect 97350 27412 97356 27424
rect 97408 27412 97414 27464
rect 176562 27412 176568 27464
rect 176620 27452 176626 27464
rect 178126 27452 178132 27464
rect 176620 27424 178132 27452
rect 176620 27412 176626 27424
rect 178126 27412 178132 27424
rect 178184 27412 178190 27464
rect 216582 27412 216588 27464
rect 216640 27452 216646 27464
rect 218054 27452 218060 27464
rect 216640 27424 218060 27452
rect 216640 27412 216646 27424
rect 218054 27412 218060 27424
rect 218112 27412 218118 27464
rect 96338 26528 96344 26580
rect 96396 26568 96402 26580
rect 97442 26568 97448 26580
rect 96396 26540 97448 26568
rect 96396 26528 96402 26540
rect 97442 26528 97448 26540
rect 97500 26528 97506 26580
rect 216858 26528 216864 26580
rect 216916 26568 216922 26580
rect 218054 26568 218060 26580
rect 216916 26540 218060 26568
rect 216916 26528 216922 26540
rect 218054 26528 218060 26540
rect 218112 26528 218118 26580
rect 257154 26256 257160 26308
rect 257212 26296 257218 26308
rect 258258 26296 258264 26308
rect 257212 26268 258264 26296
rect 257212 26256 257218 26268
rect 258258 26256 258264 26268
rect 258316 26256 258322 26308
rect 216858 25916 216864 25968
rect 216916 25956 216922 25968
rect 217962 25956 217968 25968
rect 216916 25928 217968 25956
rect 216916 25916 216922 25928
rect 217962 25916 217968 25928
rect 218020 25916 218026 25968
rect 288342 25508 288348 25560
rect 288400 25548 288406 25560
rect 580810 25548 580816 25560
rect 288400 25520 580816 25548
rect 288400 25508 288406 25520
rect 580810 25508 580816 25520
rect 580868 25508 580874 25560
rect 6178 24760 6184 24812
rect 6236 24800 6242 24812
rect 17862 24800 17868 24812
rect 6236 24772 17868 24800
rect 6236 24760 6242 24772
rect 17862 24760 17868 24772
rect 17920 24760 17926 24812
rect 65518 24760 65524 24812
rect 65576 24800 65582 24812
rect 87230 24800 87236 24812
rect 65576 24772 87236 24800
rect 65576 24760 65582 24772
rect 87230 24760 87236 24772
rect 87288 24760 87294 24812
rect 176746 24760 176752 24812
rect 176804 24800 176810 24812
rect 177850 24800 177856 24812
rect 176804 24772 177856 24800
rect 176804 24760 176810 24772
rect 177850 24760 177856 24772
rect 177908 24760 177914 24812
rect 257154 23808 257160 23860
rect 257212 23848 257218 23860
rect 258258 23848 258264 23860
rect 257212 23820 258264 23848
rect 257212 23808 257218 23820
rect 258258 23808 258264 23820
rect 258316 23808 258322 23860
rect 96338 22924 96344 22976
rect 96396 22964 96402 22976
rect 97442 22964 97448 22976
rect 96396 22936 97448 22964
rect 96396 22924 96402 22936
rect 97442 22924 97448 22936
rect 97500 22924 97506 22976
rect 176562 22924 176568 22976
rect 176620 22964 176626 22976
rect 178126 22964 178132 22976
rect 176620 22936 178132 22964
rect 176620 22924 176626 22936
rect 178126 22924 178132 22936
rect 178184 22924 178190 22976
rect 216582 22924 216588 22976
rect 216640 22964 216646 22976
rect 218054 22964 218060 22976
rect 216640 22936 218060 22964
rect 216640 22924 216646 22936
rect 218054 22924 218060 22936
rect 218112 22924 218118 22976
rect 257154 22108 257160 22160
rect 257212 22148 257218 22160
rect 258258 22148 258264 22160
rect 257212 22120 258264 22148
rect 257212 22108 257218 22120
rect 258258 22108 258264 22120
rect 258316 22108 258322 22160
rect 14458 22040 14464 22092
rect 14516 22080 14522 22092
rect 17770 22080 17776 22092
rect 14516 22052 17776 22080
rect 14516 22040 14522 22052
rect 17770 22040 17776 22052
rect 17828 22040 17834 22092
rect 96338 21428 96344 21480
rect 96396 21468 96402 21480
rect 97442 21468 97448 21480
rect 96396 21440 97448 21468
rect 96396 21428 96402 21440
rect 97442 21428 97448 21440
rect 97500 21428 97506 21480
rect 176562 21428 176568 21480
rect 176620 21468 176626 21480
rect 178126 21468 178132 21480
rect 176620 21440 178132 21468
rect 176620 21428 176626 21440
rect 178126 21428 178132 21440
rect 178184 21428 178190 21480
rect 216582 21428 216588 21480
rect 216640 21468 216646 21480
rect 218054 21468 218060 21480
rect 216640 21440 218060 21468
rect 216640 21428 216646 21440
rect 218054 21428 218060 21440
rect 218112 21428 218118 21480
rect 216582 20680 216588 20732
rect 216640 20720 216646 20732
rect 218054 20720 218060 20732
rect 216640 20692 218060 20720
rect 216640 20680 216646 20692
rect 218054 20680 218060 20692
rect 218112 20680 218118 20732
rect 3418 20612 3424 20664
rect 3476 20652 3482 20664
rect 19702 20652 19708 20664
rect 3476 20624 19708 20652
rect 3476 20612 3482 20624
rect 19702 20612 19708 20624
rect 19760 20612 19766 20664
rect 87414 20652 87420 20664
rect 19904 20624 87420 20652
rect 3234 20544 3240 20596
rect 3292 20584 3298 20596
rect 3292 20556 6914 20584
rect 3292 20544 3298 20556
rect 6886 20448 6914 20556
rect 17862 20476 17868 20528
rect 17920 20516 17926 20528
rect 19904 20516 19932 20624
rect 87414 20612 87420 20624
rect 87472 20612 87478 20664
rect 67634 20584 67640 20596
rect 17920 20488 19932 20516
rect 26206 20556 67640 20584
rect 17920 20476 17926 20488
rect 26206 20448 26234 20556
rect 67634 20544 67640 20556
rect 67692 20544 67698 20596
rect 6886 20420 26234 20448
rect 88150 19932 88156 19984
rect 88208 19972 88214 19984
rect 127526 19972 127532 19984
rect 88208 19944 127532 19972
rect 88208 19932 88214 19944
rect 127526 19932 127532 19944
rect 127584 19932 127590 19984
rect 169570 19932 169576 19984
rect 169628 19972 169634 19984
rect 208486 19972 208492 19984
rect 169628 19944 208492 19972
rect 169628 19932 169634 19944
rect 208486 19932 208492 19944
rect 208544 19932 208550 19984
rect 88058 19864 88064 19916
rect 88116 19904 88122 19916
rect 127618 19904 127624 19916
rect 88116 19876 127624 19904
rect 88116 19864 88122 19876
rect 127618 19864 127624 19876
rect 127676 19864 127682 19916
rect 169478 19864 169484 19916
rect 169536 19904 169542 19916
rect 209038 19904 209044 19916
rect 169536 19876 209044 19904
rect 169536 19864 169542 19876
rect 209038 19864 209044 19876
rect 209096 19864 209102 19916
rect 95878 19796 95884 19848
rect 95936 19836 95942 19848
rect 126974 19836 126980 19848
rect 95936 19808 126980 19836
rect 95936 19796 95942 19808
rect 126974 19796 126980 19808
rect 127032 19796 127038 19848
rect 175918 19796 175924 19848
rect 175976 19836 175982 19848
rect 208394 19836 208400 19848
rect 175976 19808 208400 19836
rect 175976 19796 175982 19808
rect 208394 19796 208400 19808
rect 208452 19796 208458 19848
rect 128262 19524 128268 19576
rect 128320 19564 128326 19576
rect 168374 19564 168380 19576
rect 128320 19536 168380 19564
rect 128320 19524 128326 19536
rect 168374 19524 168380 19536
rect 168432 19524 168438 19576
rect 127986 19456 127992 19508
rect 128044 19496 128050 19508
rect 169018 19496 169024 19508
rect 128044 19468 169024 19496
rect 128044 19456 128050 19468
rect 169018 19456 169024 19468
rect 169076 19456 169082 19508
rect 66162 19252 66168 19304
rect 66220 19292 66226 19304
rect 288342 19292 288348 19304
rect 66220 19264 288348 19292
rect 66220 19252 66226 19264
rect 288342 19252 288348 19264
rect 288400 19252 288406 19304
rect 42610 19184 42616 19236
rect 42668 19224 42674 19236
rect 87598 19224 87604 19236
rect 42668 19196 87604 19224
rect 42668 19184 42674 19196
rect 87598 19184 87604 19196
rect 87656 19184 87662 19236
rect 128170 19184 128176 19236
rect 128228 19224 128234 19236
rect 169110 19224 169116 19236
rect 128228 19196 169116 19224
rect 128228 19184 128234 19196
rect 169110 19184 169116 19196
rect 169168 19184 169174 19236
rect 209406 19184 209412 19236
rect 209464 19224 209470 19236
rect 249058 19224 249064 19236
rect 209464 19196 249064 19224
rect 209464 19184 209470 19196
rect 249058 19184 249064 19196
rect 249116 19184 249122 19236
rect 209682 19116 209688 19168
rect 209740 19156 209746 19168
rect 249702 19156 249708 19168
rect 209740 19128 249708 19156
rect 209740 19116 209746 19128
rect 249702 19116 249708 19128
rect 249760 19116 249766 19168
rect 209590 19048 209596 19100
rect 209648 19088 209654 19100
rect 248598 19088 248604 19100
rect 209648 19060 248604 19088
rect 209648 19048 209654 19060
rect 248598 19048 248604 19060
rect 248656 19048 248662 19100
rect 209498 18980 209504 19032
rect 209556 19020 209562 19032
rect 249150 19020 249156 19032
rect 209556 18992 249156 19020
rect 209556 18980 209562 18992
rect 249150 18980 249156 18992
rect 249208 18980 249214 19032
rect 4062 17892 4068 17944
rect 4120 17932 4126 17944
rect 29638 17932 29644 17944
rect 4120 17904 29644 17932
rect 4120 17892 4126 17904
rect 29638 17892 29644 17904
rect 29696 17892 29702 17944
rect 43898 17892 43904 17944
rect 43956 17932 43962 17944
rect 72970 17932 72976 17944
rect 43956 17904 72976 17932
rect 43956 17892 43962 17904
rect 72970 17892 72976 17904
rect 73028 17892 73034 17944
rect 3510 17824 3516 17876
rect 3568 17864 3574 17876
rect 34146 17864 34152 17876
rect 3568 17836 34152 17864
rect 3568 17824 3574 17836
rect 34146 17824 34152 17836
rect 34204 17824 34210 17876
rect 40678 17824 40684 17876
rect 40736 17864 40742 17876
rect 580534 17864 580540 17876
rect 40736 17836 580540 17864
rect 40736 17824 40742 17836
rect 580534 17824 580540 17836
rect 580592 17824 580598 17876
rect 47118 17756 47124 17808
rect 47176 17796 47182 17808
rect 580626 17796 580632 17808
rect 47176 17768 580632 17796
rect 47176 17756 47182 17768
rect 580626 17756 580632 17768
rect 580684 17756 580690 17808
rect 3970 17688 3976 17740
rect 4028 17728 4034 17740
rect 26418 17728 26424 17740
rect 4028 17700 26424 17728
rect 4028 17688 4034 17700
rect 26418 17688 26424 17700
rect 26476 17688 26482 17740
rect 49050 17688 49056 17740
rect 49108 17728 49114 17740
rect 580350 17728 580356 17740
rect 49108 17700 580356 17728
rect 49108 17688 49114 17700
rect 580350 17688 580356 17700
rect 580408 17688 580414 17740
rect 3602 17620 3608 17672
rect 3660 17660 3666 17672
rect 58618 17660 58624 17672
rect 3660 17632 58624 17660
rect 3660 17620 3666 17632
rect 58618 17620 58624 17632
rect 58676 17620 58682 17672
rect 63862 17620 63868 17672
rect 63920 17660 63926 17672
rect 580442 17660 580448 17672
rect 63920 17632 580448 17660
rect 63920 17620 63926 17632
rect 580442 17620 580448 17632
rect 580500 17620 580506 17672
rect 8110 17552 8116 17604
rect 8168 17592 8174 17604
rect 59906 17592 59912 17604
rect 8168 17564 59912 17592
rect 8168 17552 8174 17564
rect 59906 17552 59912 17564
rect 59964 17552 59970 17604
rect 65150 17552 65156 17604
rect 65208 17592 65214 17604
rect 580258 17592 580264 17604
rect 65208 17564 580264 17592
rect 65208 17552 65214 17564
rect 580258 17552 580264 17564
rect 580316 17552 580322 17604
rect 23290 17484 23296 17536
rect 23348 17524 23354 17536
rect 527174 17524 527180 17536
rect 23348 17496 527180 17524
rect 23348 17484 23354 17496
rect 527174 17484 527180 17496
rect 527232 17484 527238 17536
rect 3694 17416 3700 17468
rect 3752 17456 3758 17468
rect 55398 17456 55404 17468
rect 3752 17428 55404 17456
rect 3752 17416 3758 17428
rect 55398 17416 55404 17428
rect 55456 17416 55462 17468
rect 56778 17416 56784 17468
rect 56836 17456 56842 17468
rect 559650 17456 559656 17468
rect 56836 17428 559656 17456
rect 56836 17416 56842 17428
rect 559650 17416 559656 17428
rect 559708 17416 559714 17468
rect 45830 17348 45836 17400
rect 45888 17388 45894 17400
rect 429838 17388 429844 17400
rect 45888 17360 429844 17388
rect 45888 17348 45894 17360
rect 429838 17348 429844 17360
rect 429896 17348 429902 17400
rect 31018 17280 31024 17332
rect 31076 17320 31082 17332
rect 397454 17320 397460 17332
rect 31076 17292 397460 17320
rect 31076 17280 31082 17292
rect 397454 17280 397460 17292
rect 397512 17280 397518 17332
rect 36170 17212 36176 17264
rect 36228 17252 36234 17264
rect 366358 17252 366364 17264
rect 36228 17224 366364 17252
rect 36228 17212 36234 17224
rect 366358 17212 366364 17224
rect 366416 17212 366422 17264
rect 52270 17144 52276 17196
rect 52328 17184 52334 17196
rect 170306 17184 170312 17196
rect 52328 17156 170312 17184
rect 52328 17144 52334 17156
rect 170306 17144 170312 17156
rect 170364 17144 170370 17196
rect 27798 17076 27804 17128
rect 27856 17116 27862 17128
rect 137738 17116 137744 17128
rect 27856 17088 137744 17116
rect 27856 17076 27862 17088
rect 137738 17076 137744 17088
rect 137796 17076 137802 17128
rect 24578 17008 24584 17060
rect 24636 17048 24642 17060
rect 580718 17048 580724 17060
rect 24636 17020 580724 17048
rect 24636 17008 24642 17020
rect 580718 17008 580724 17020
rect 580776 17008 580782 17060
rect 1670 3544 1676 3596
rect 1728 3584 1734 3596
rect 37274 3584 37280 3596
rect 1728 3556 37280 3584
rect 1728 3544 1734 3556
rect 37274 3544 37280 3556
rect 37332 3544 37338 3596
rect 68462 3544 68468 3596
rect 68520 3584 68526 3596
rect 125870 3584 125876 3596
rect 68520 3556 125876 3584
rect 68520 3544 68526 3556
rect 125870 3544 125876 3556
rect 125928 3544 125934 3596
rect 17862 3476 17868 3528
rect 17920 3516 17926 3528
rect 129366 3516 129372 3528
rect 17920 3488 129372 3516
rect 17920 3476 17926 3488
rect 129366 3476 129372 3488
rect 129424 3476 129430 3528
rect 566 3408 572 3460
rect 624 3448 630 3460
rect 52454 3448 52460 3460
rect 624 3420 52460 3448
rect 624 3408 630 3420
rect 52454 3408 52460 3420
rect 52512 3408 52518 3460
rect 68370 3408 68376 3460
rect 68428 3448 68434 3460
rect 126974 3448 126980 3460
rect 68428 3420 126980 3448
rect 68428 3408 68434 3420
rect 126974 3408 126980 3420
rect 127032 3408 127038 3460
<< via1 >>
rect 31668 700816 31720 700868
rect 105452 700816 105504 700868
rect 62028 700748 62080 700800
rect 202788 700748 202840 700800
rect 71044 700680 71096 700732
rect 267648 700680 267700 700732
rect 23388 700612 23440 700664
rect 235172 700612 235224 700664
rect 64788 700544 64840 700596
rect 332508 700544 332560 700596
rect 17868 700476 17920 700528
rect 300124 700476 300176 700528
rect 68284 700408 68336 700460
rect 364984 700408 365036 700460
rect 28908 700340 28960 700392
rect 462320 700340 462372 700392
rect 50988 700272 51040 700324
rect 494796 700272 494848 700324
rect 57888 696940 57940 696992
rect 580172 696940 580224 696992
rect 3516 656888 3568 656940
rect 19984 656888 20036 656940
rect 3516 632068 3568 632120
rect 18604 632068 18656 632120
rect 68376 590656 68428 590708
rect 580172 590656 580224 590708
rect 22008 563048 22060 563100
rect 580172 563048 580224 563100
rect 3332 553392 3384 553444
rect 24124 553392 24176 553444
rect 68468 536800 68520 536852
rect 580172 536800 580224 536852
rect 2780 527144 2832 527196
rect 6184 527144 6236 527196
rect 30288 510620 30340 510672
rect 580172 510620 580224 510672
rect 68560 470568 68612 470620
rect 579988 470568 580040 470620
rect 3148 448536 3200 448588
rect 43444 448536 43496 448588
rect 17776 430584 17828 430636
rect 579620 430584 579672 430636
rect 17684 404336 17736 404388
rect 580172 404336 580224 404388
rect 68652 378156 68704 378208
rect 580172 378156 580224 378208
rect 3332 357416 3384 357468
rect 65340 357416 65392 357468
rect 3332 345040 3384 345092
rect 13084 345040 13136 345092
rect 3332 292544 3384 292596
rect 14464 292544 14516 292596
rect 3332 253920 3384 253972
rect 33784 253920 33836 253972
rect 39948 231820 40000 231872
rect 579804 231820 579856 231872
rect 3332 201492 3384 201544
rect 65248 201492 65300 201544
rect 66168 191836 66220 191888
rect 580172 191836 580224 191888
rect 56508 151784 56560 151836
rect 579988 151784 580040 151836
rect 3332 136620 3384 136672
rect 15844 136620 15896 136672
rect 36636 52572 36688 52624
rect 249064 52572 249116 52624
rect 17592 52504 17644 52556
rect 249156 52504 249208 52556
rect 33048 52436 33100 52488
rect 287704 52436 287756 52488
rect 176568 51076 176620 51128
rect 178132 51076 178184 51128
rect 216588 51076 216640 51128
rect 218060 51076 218112 51128
rect 96528 48288 96580 48340
rect 97448 48288 97500 48340
rect 176476 48288 176528 48340
rect 178132 48288 178184 48340
rect 217324 48288 217376 48340
rect 218060 48288 218112 48340
rect 96252 46928 96304 46980
rect 97448 46928 97500 46980
rect 216496 46928 216548 46980
rect 218060 46928 218112 46980
rect 257344 46928 257396 46980
rect 258264 46928 258316 46980
rect 3424 46180 3476 46232
rect 58624 46180 58676 46232
rect 3424 46044 3476 46096
rect 3792 46044 3844 46096
rect 2964 44140 3016 44192
rect 16488 44140 16540 44192
rect 96344 44140 96396 44192
rect 97448 44140 97500 44192
rect 257252 44140 257304 44192
rect 258264 44140 258316 44192
rect 216404 43052 216456 43104
rect 217968 43052 218020 43104
rect 176292 42780 176344 42832
rect 178132 42780 178184 42832
rect 19984 42712 20036 42764
rect 26424 42712 26476 42764
rect 33784 42712 33836 42764
rect 37372 42712 37424 42764
rect 43444 42712 43496 42764
rect 45744 42712 45796 42764
rect 257160 42644 257212 42696
rect 258172 42644 258224 42696
rect 18604 42372 18656 42424
rect 24492 42372 24544 42424
rect 65156 42372 65208 42424
rect 66168 42372 66220 42424
rect 24124 42168 24176 42220
rect 34152 42168 34204 42220
rect 40500 42168 40552 42220
rect 52184 42168 52236 42220
rect 3424 42100 3476 42152
rect 42524 42100 42576 42152
rect 3792 42032 3844 42084
rect 48964 42032 49016 42084
rect 91008 41964 91060 42016
rect 95884 41964 95936 42016
rect 131028 41964 131080 42016
rect 135904 41964 135956 42016
rect 171416 41964 171468 42016
rect 175924 41964 175976 42016
rect 40684 41420 40736 41472
rect 65524 41420 65576 41472
rect 366364 40672 366416 40724
rect 580908 40672 580960 40724
rect 176384 40060 176436 40112
rect 178132 40060 178184 40112
rect 17684 39992 17736 40044
rect 19708 39992 19760 40044
rect 176568 39380 176620 39432
rect 178040 39380 178092 39432
rect 176476 38632 176528 38684
rect 178132 38632 178184 38684
rect 176752 37884 176804 37936
rect 177856 37884 177908 37936
rect 216588 37884 216640 37936
rect 218060 37884 218112 37936
rect 96344 37136 96396 37188
rect 97448 37136 97500 37188
rect 257344 35912 257396 35964
rect 258264 35912 258316 35964
rect 3240 35844 3292 35896
rect 17868 35844 17920 35896
rect 176752 34484 176804 34536
rect 177856 34484 177908 34536
rect 216864 34484 216916 34536
rect 217968 34484 218020 34536
rect 257160 34484 257212 34536
rect 258264 34484 258316 34536
rect 287704 33056 287756 33108
rect 580172 33056 580224 33108
rect 96344 32920 96396 32972
rect 97448 32920 97500 32972
rect 216496 32852 216548 32904
rect 217968 32852 218020 32904
rect 176568 31900 176620 31952
rect 178132 31900 178184 31952
rect 216588 31900 216640 31952
rect 218060 31900 218112 31952
rect 67732 31424 67784 31476
rect 71044 31424 71096 31476
rect 96344 28908 96396 28960
rect 97540 28908 97592 28960
rect 176568 28908 176620 28960
rect 178040 28908 178092 28960
rect 96528 27616 96580 27668
rect 97448 27616 97500 27668
rect 176752 27616 176804 27668
rect 177856 27616 177908 27668
rect 257344 27616 257396 27668
rect 258264 27616 258316 27668
rect 13084 27548 13136 27600
rect 17868 27548 17920 27600
rect 96344 27412 96396 27464
rect 97356 27412 97408 27464
rect 176568 27412 176620 27464
rect 178132 27412 178184 27464
rect 216588 27412 216640 27464
rect 218060 27412 218112 27464
rect 96344 26528 96396 26580
rect 97448 26528 97500 26580
rect 216864 26528 216916 26580
rect 218060 26528 218112 26580
rect 257160 26256 257212 26308
rect 258264 26256 258316 26308
rect 216864 25916 216916 25968
rect 217968 25916 218020 25968
rect 288348 25508 288400 25560
rect 580816 25508 580868 25560
rect 6184 24760 6236 24812
rect 17868 24760 17920 24812
rect 65524 24760 65576 24812
rect 87236 24760 87288 24812
rect 176752 24760 176804 24812
rect 177856 24760 177908 24812
rect 257160 23808 257212 23860
rect 258264 23808 258316 23860
rect 96344 22924 96396 22976
rect 97448 22924 97500 22976
rect 176568 22924 176620 22976
rect 178132 22924 178184 22976
rect 216588 22924 216640 22976
rect 218060 22924 218112 22976
rect 257160 22108 257212 22160
rect 258264 22108 258316 22160
rect 14464 22040 14516 22092
rect 17776 22040 17828 22092
rect 96344 21428 96396 21480
rect 97448 21428 97500 21480
rect 176568 21428 176620 21480
rect 178132 21428 178184 21480
rect 216588 21428 216640 21480
rect 218060 21428 218112 21480
rect 216588 20680 216640 20732
rect 218060 20680 218112 20732
rect 3424 20612 3476 20664
rect 19708 20612 19760 20664
rect 3240 20544 3292 20596
rect 17868 20476 17920 20528
rect 87420 20612 87472 20664
rect 67640 20544 67692 20596
rect 88156 19932 88208 19984
rect 127532 19932 127584 19984
rect 169576 19932 169628 19984
rect 208492 19932 208544 19984
rect 88064 19864 88116 19916
rect 127624 19864 127676 19916
rect 169484 19864 169536 19916
rect 209044 19864 209096 19916
rect 95884 19796 95936 19848
rect 126980 19796 127032 19848
rect 175924 19796 175976 19848
rect 208400 19796 208452 19848
rect 128268 19524 128320 19576
rect 168380 19524 168432 19576
rect 127992 19456 128044 19508
rect 169024 19456 169076 19508
rect 66168 19252 66220 19304
rect 288348 19252 288400 19304
rect 42616 19184 42668 19236
rect 87604 19184 87656 19236
rect 128176 19184 128228 19236
rect 169116 19184 169168 19236
rect 209412 19184 209464 19236
rect 249064 19184 249116 19236
rect 209688 19116 209740 19168
rect 249708 19116 249760 19168
rect 209596 19048 209648 19100
rect 248604 19048 248656 19100
rect 209504 18980 209556 19032
rect 249156 18980 249208 19032
rect 4068 17892 4120 17944
rect 29644 17892 29696 17944
rect 43904 17892 43956 17944
rect 72976 17892 73028 17944
rect 3516 17824 3568 17876
rect 34152 17824 34204 17876
rect 40684 17824 40736 17876
rect 580540 17824 580592 17876
rect 47124 17756 47176 17808
rect 580632 17756 580684 17808
rect 3976 17688 4028 17740
rect 26424 17688 26476 17740
rect 49056 17688 49108 17740
rect 580356 17688 580408 17740
rect 3608 17620 3660 17672
rect 58624 17620 58676 17672
rect 63868 17620 63920 17672
rect 580448 17620 580500 17672
rect 8116 17552 8168 17604
rect 59912 17552 59964 17604
rect 65156 17552 65208 17604
rect 580264 17552 580316 17604
rect 23296 17484 23348 17536
rect 527180 17484 527232 17536
rect 3700 17416 3752 17468
rect 55404 17416 55456 17468
rect 56784 17416 56836 17468
rect 559656 17416 559708 17468
rect 45836 17348 45888 17400
rect 429844 17348 429896 17400
rect 31024 17280 31076 17332
rect 397460 17280 397512 17332
rect 36176 17212 36228 17264
rect 366364 17212 366416 17264
rect 52276 17144 52328 17196
rect 170312 17144 170364 17196
rect 27804 17076 27856 17128
rect 137744 17076 137796 17128
rect 24584 17008 24636 17060
rect 580724 17008 580776 17060
rect 1676 3544 1728 3596
rect 37280 3544 37332 3596
rect 68468 3544 68520 3596
rect 125876 3544 125928 3596
rect 17868 3476 17920 3528
rect 129372 3476 129424 3528
rect 572 3408 624 3460
rect 52460 3408 52512 3460
rect 68376 3408 68428 3460
rect 126980 3408 127032 3460
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 3422 684312 3478 684321
rect 3422 684247 3478 684256
rect 3330 553888 3386 553897
rect 3330 553823 3386 553832
rect 3344 553450 3372 553823
rect 3332 553444 3384 553450
rect 3332 553386 3384 553392
rect 2778 527912 2834 527921
rect 2778 527847 2834 527856
rect 2792 527202 2820 527847
rect 2780 527196 2832 527202
rect 2780 527138 2832 527144
rect 3146 449576 3202 449585
rect 3146 449511 3202 449520
rect 3160 448594 3188 449511
rect 3148 448588 3200 448594
rect 3148 448530 3200 448536
rect 3330 358456 3386 358465
rect 3330 358391 3386 358400
rect 3344 357474 3372 358391
rect 3332 357468 3384 357474
rect 3332 357410 3384 357416
rect 3330 345400 3386 345409
rect 3330 345335 3386 345344
rect 3344 345098 3372 345335
rect 3332 345092 3384 345098
rect 3332 345034 3384 345040
rect 3330 293176 3386 293185
rect 3330 293111 3386 293120
rect 3344 292602 3372 293111
rect 3332 292596 3384 292602
rect 3332 292538 3384 292544
rect 3330 254144 3386 254153
rect 3330 254079 3386 254088
rect 3344 253978 3372 254079
rect 3332 253972 3384 253978
rect 3332 253914 3384 253920
rect 3330 201920 3386 201929
rect 3330 201855 3386 201864
rect 3344 201550 3372 201855
rect 3332 201544 3384 201550
rect 3332 201486 3384 201492
rect 3330 136776 3386 136785
rect 3330 136711 3386 136720
rect 3344 136678 3372 136711
rect 3332 136672 3384 136678
rect 3332 136614 3384 136620
rect 3330 84688 3386 84697
rect 3330 84623 3386 84632
rect 3238 58576 3294 58585
rect 3238 58511 3294 58520
rect 2962 45520 3018 45529
rect 2962 45455 3018 45464
rect 2976 44198 3004 45455
rect 2964 44192 3016 44198
rect 2964 44134 3016 44140
rect 3252 35902 3280 58511
rect 3240 35896 3292 35902
rect 3344 35894 3372 84623
rect 3436 46238 3464 684247
rect 3514 658200 3570 658209
rect 3514 658135 3570 658144
rect 3528 656946 3556 658135
rect 3516 656940 3568 656946
rect 3516 656882 3568 656888
rect 3516 632120 3568 632126
rect 3514 632088 3516 632097
rect 3568 632088 3570 632097
rect 3514 632023 3570 632032
rect 6184 527196 6236 527202
rect 6184 527138 6236 527144
rect 3514 410544 3570 410553
rect 3514 410479 3570 410488
rect 3424 46232 3476 46238
rect 3424 46174 3476 46180
rect 3424 46096 3476 46102
rect 3424 46038 3476 46044
rect 3436 42158 3464 46038
rect 3424 42152 3476 42158
rect 3424 42094 3476 42100
rect 3344 35866 3464 35894
rect 3240 35838 3292 35844
rect 3436 20670 3464 35866
rect 3424 20664 3476 20670
rect 3424 20606 3476 20612
rect 3240 20596 3292 20602
rect 3240 20538 3292 20544
rect 3252 19417 3280 20538
rect 3238 19408 3294 19417
rect 3238 19343 3294 19352
rect 3528 17882 3556 410479
rect 3606 397488 3662 397497
rect 3606 397423 3662 397432
rect 3516 17876 3568 17882
rect 3516 17818 3568 17824
rect 3620 17678 3648 397423
rect 3698 306232 3754 306241
rect 3698 306167 3754 306176
rect 3608 17672 3660 17678
rect 3608 17614 3660 17620
rect 3712 17474 3740 306167
rect 3790 241088 3846 241097
rect 3790 241023 3846 241032
rect 3804 46102 3832 241023
rect 3882 188864 3938 188873
rect 3882 188799 3938 188808
rect 3792 46096 3844 46102
rect 3792 46038 3844 46044
rect 3896 45554 3924 188799
rect 3974 149832 4030 149841
rect 3974 149767 4030 149776
rect 3804 45526 3924 45554
rect 3804 42090 3832 45526
rect 3792 42084 3844 42090
rect 3792 42026 3844 42032
rect 3988 17746 4016 149767
rect 4066 97608 4122 97617
rect 4066 97543 4122 97552
rect 4080 17950 4108 97543
rect 6196 24818 6224 527138
rect 6184 24812 6236 24818
rect 6184 24754 6236 24760
rect 4068 17944 4120 17950
rect 4068 17886 4120 17892
rect 3976 17740 4028 17746
rect 3976 17682 4028 17688
rect 8128 17610 8156 703520
rect 31668 700868 31720 700874
rect 31668 700810 31720 700816
rect 23388 700664 23440 700670
rect 23388 700606 23440 700612
rect 17868 700528 17920 700534
rect 17868 700470 17920 700476
rect 17776 430636 17828 430642
rect 17776 430578 17828 430584
rect 17684 404388 17736 404394
rect 17684 404330 17736 404336
rect 13084 345092 13136 345098
rect 13084 345034 13136 345040
rect 13096 27606 13124 345034
rect 14464 292596 14516 292602
rect 14464 292538 14516 292544
rect 13084 27600 13136 27606
rect 13084 27542 13136 27548
rect 14476 22098 14504 292538
rect 15844 136672 15896 136678
rect 15844 136614 15896 136620
rect 15856 24177 15884 136614
rect 17592 52556 17644 52562
rect 17592 52498 17644 52504
rect 16488 44192 16540 44198
rect 16488 44134 16540 44140
rect 16500 37913 16528 44134
rect 16486 37904 16542 37913
rect 16486 37839 16542 37848
rect 17604 31657 17632 52498
rect 17696 40050 17724 404330
rect 17684 40044 17736 40050
rect 17684 39986 17736 39992
rect 17788 33697 17816 430578
rect 17880 37097 17908 700470
rect 19984 656940 20036 656946
rect 19984 656882 20036 656888
rect 18604 632120 18656 632126
rect 18604 632062 18656 632068
rect 18616 42430 18644 632062
rect 19996 42770 20024 656882
rect 22008 563100 22060 563106
rect 22008 563042 22060 563048
rect 22020 45554 22048 563042
rect 21744 45526 22048 45554
rect 19984 42764 20036 42770
rect 19984 42706 20036 42712
rect 18604 42424 18656 42430
rect 18604 42366 18656 42372
rect 19708 40044 19760 40050
rect 19708 39986 19760 39992
rect 19720 39930 19748 39986
rect 21744 39930 21772 45526
rect 23400 39930 23428 700606
rect 28908 700392 28960 700398
rect 28908 700334 28960 700340
rect 24124 553444 24176 553450
rect 24124 553386 24176 553392
rect 24136 42226 24164 553386
rect 28920 45554 28948 700334
rect 30288 510672 30340 510678
rect 30288 510614 30340 510620
rect 30300 45554 30328 510614
rect 31680 45554 31708 700810
rect 33784 253972 33836 253978
rect 33784 253914 33836 253920
rect 33048 52488 33100 52494
rect 33048 52430 33100 52436
rect 28184 45526 28948 45554
rect 30208 45526 30328 45554
rect 31496 45526 31708 45554
rect 26424 42764 26476 42770
rect 26424 42706 26476 42712
rect 24492 42424 24544 42430
rect 24492 42366 24544 42372
rect 24124 42220 24176 42226
rect 24124 42162 24176 42168
rect 19720 39902 20010 39930
rect 21390 39902 21772 39930
rect 23322 39902 23428 39930
rect 24504 39916 24532 42366
rect 26436 39916 26464 42706
rect 28184 39930 28212 45526
rect 30208 39930 30236 45526
rect 31496 39930 31524 45526
rect 33060 39930 33088 52430
rect 33796 42770 33824 253914
rect 39948 231872 40000 231878
rect 39948 231814 40000 231820
rect 36636 52624 36688 52630
rect 36636 52566 36688 52572
rect 33784 42764 33836 42770
rect 33784 42706 33836 42712
rect 34152 42220 34204 42226
rect 34152 42162 34204 42168
rect 27830 39902 28212 39930
rect 29762 39902 30236 39930
rect 31050 39902 31524 39930
rect 32982 39902 33088 39930
rect 34164 39916 34192 42162
rect 36648 39930 36676 52566
rect 39960 45554 39988 231814
rect 39776 45526 39988 45554
rect 37372 42764 37424 42770
rect 37372 42706 37424 42712
rect 36202 39902 36676 39930
rect 37384 39916 37412 42706
rect 39776 39930 39804 45526
rect 40512 42226 40540 703520
rect 62028 700800 62080 700806
rect 62028 700742 62080 700748
rect 50988 700324 51040 700330
rect 50988 700266 51040 700272
rect 43444 448588 43496 448594
rect 43444 448530 43496 448536
rect 43456 42770 43484 448530
rect 43444 42764 43496 42770
rect 43444 42706 43496 42712
rect 45744 42764 45796 42770
rect 45744 42706 45796 42712
rect 40500 42220 40552 42226
rect 40500 42162 40552 42168
rect 42524 42152 42576 42158
rect 42524 42094 42576 42100
rect 40684 41472 40736 41478
rect 40684 41414 40736 41420
rect 39422 39902 39804 39930
rect 40696 39916 40724 41414
rect 42536 39916 42564 42094
rect 45756 39916 45784 42706
rect 48964 42084 49016 42090
rect 48964 42026 49016 42032
rect 48976 39916 49004 42026
rect 51000 39916 51028 700266
rect 57888 696992 57940 696998
rect 57888 696934 57940 696940
rect 56508 151836 56560 151842
rect 56508 151778 56560 151784
rect 56520 45554 56548 151778
rect 57900 45554 57928 696934
rect 58624 46232 58676 46238
rect 58624 46174 58676 46180
rect 55968 45526 56548 45554
rect 57808 45526 57928 45554
rect 52184 42220 52236 42226
rect 52184 42162 52236 42168
rect 52196 39916 52224 42162
rect 55968 39930 55996 45526
rect 57808 39930 57836 45526
rect 55522 39902 55996 39930
rect 57454 39902 57836 39930
rect 58636 39916 58664 46174
rect 62040 39930 62068 700742
rect 71044 700732 71096 700738
rect 71044 700674 71096 700680
rect 64788 700596 64840 700602
rect 64788 700538 64840 700544
rect 64800 45554 64828 700538
rect 68284 700460 68336 700466
rect 68284 700402 68336 700408
rect 65340 357468 65392 357474
rect 65340 357410 65392 357416
rect 65248 201544 65300 201550
rect 65248 201486 65300 201492
rect 64248 45526 64828 45554
rect 64248 39930 64276 45526
rect 65156 42424 65208 42430
rect 65156 42366 65208 42372
rect 61962 39902 62068 39930
rect 63894 39902 64276 39930
rect 65168 39916 65196 42366
rect 43994 39400 44050 39409
rect 43930 39358 43994 39386
rect 43994 39335 44050 39344
rect 47306 39400 47362 39409
rect 54574 39400 54630 39409
rect 47362 39358 47702 39386
rect 54234 39358 54574 39386
rect 47306 39335 47362 39344
rect 54574 39335 54630 39344
rect 60545 39208 60554 39264
rect 60610 39208 60619 39264
rect 17866 37088 17922 37097
rect 17866 37023 17922 37032
rect 17868 35896 17920 35902
rect 65260 35894 65288 201486
rect 65352 38321 65380 357410
rect 66168 191888 66220 191894
rect 66168 191830 66220 191836
rect 66180 42430 66208 191830
rect 66168 42424 66220 42430
rect 66168 42366 66220 42372
rect 65524 41472 65576 41478
rect 65524 41414 65576 41420
rect 65338 38312 65394 38321
rect 65338 38247 65394 38256
rect 65260 35866 65380 35894
rect 17868 35838 17920 35844
rect 17880 35057 17908 35838
rect 17866 35048 17922 35057
rect 17866 34983 17922 34992
rect 17774 33688 17830 33697
rect 17774 33623 17830 33632
rect 17590 31648 17646 31657
rect 17590 31583 17646 31592
rect 17774 30288 17830 30297
rect 17774 30223 17830 30232
rect 17682 28248 17738 28257
rect 17682 28183 17738 28192
rect 15842 24168 15898 24177
rect 15842 24103 15898 24112
rect 14464 22092 14516 22098
rect 14464 22034 14516 22040
rect 8116 17604 8168 17610
rect 8116 17546 8168 17552
rect 3700 17468 3752 17474
rect 3700 17410 3752 17416
rect 17696 16574 17724 28183
rect 17788 23474 17816 30223
rect 17868 27600 17920 27606
rect 17868 27542 17920 27548
rect 17880 26897 17908 27542
rect 17866 26888 17922 26897
rect 17866 26823 17922 26832
rect 17866 24848 17922 24857
rect 17866 24783 17868 24792
rect 17920 24783 17922 24792
rect 17868 24754 17920 24760
rect 65352 24721 65380 35866
rect 65536 24818 65564 41414
rect 67732 31476 67784 31482
rect 67732 31418 67784 31424
rect 67744 30977 67772 31418
rect 67730 30968 67786 30977
rect 67730 30903 67786 30912
rect 68296 27577 68324 700402
rect 68376 590708 68428 590714
rect 68376 590650 68428 590656
rect 68388 35737 68416 590650
rect 68468 536852 68520 536858
rect 68468 536794 68520 536800
rect 68374 35728 68430 35737
rect 68374 35663 68430 35672
rect 68374 34368 68430 34377
rect 68374 34303 68430 34312
rect 68282 27568 68338 27577
rect 68282 27503 68338 27512
rect 67638 25528 67694 25537
rect 67638 25463 67694 25472
rect 65524 24812 65576 24818
rect 65524 24754 65576 24760
rect 65338 24712 65394 24721
rect 65338 24647 65394 24656
rect 17788 23446 17908 23474
rect 17776 22092 17828 22098
rect 17776 22034 17828 22040
rect 17788 21457 17816 22034
rect 17774 21448 17830 21457
rect 17774 21383 17830 21392
rect 17880 20534 17908 23446
rect 19708 20664 19760 20670
rect 21638 20632 21694 20641
rect 19760 20612 20010 20618
rect 19708 20606 20010 20612
rect 19720 20590 20010 20606
rect 21390 20590 21638 20618
rect 21638 20567 21694 20576
rect 66166 20632 66222 20641
rect 67652 20602 67680 25463
rect 66166 20567 66222 20576
rect 67640 20596 67692 20602
rect 17868 20528 17920 20534
rect 17868 20470 17920 20476
rect 23308 17542 23336 20060
rect 23296 17536 23348 17542
rect 23296 17478 23348 17484
rect 24596 17066 24624 20060
rect 26436 17746 26464 20060
rect 26424 17740 26476 17746
rect 26424 17682 26476 17688
rect 27816 17134 27844 20060
rect 29656 17950 29684 20060
rect 29644 17944 29696 17950
rect 29644 17886 29696 17892
rect 31036 17338 31064 20060
rect 32876 17513 32904 20060
rect 34164 17882 34192 20060
rect 34152 17876 34204 17882
rect 34152 17818 34204 17824
rect 32862 17504 32918 17513
rect 32862 17439 32918 17448
rect 31024 17332 31076 17338
rect 31024 17274 31076 17280
rect 36188 17270 36216 20060
rect 37292 20046 37398 20074
rect 36176 17264 36228 17270
rect 36176 17206 36228 17212
rect 27804 17128 27856 17134
rect 27804 17070 27856 17076
rect 24584 17060 24636 17066
rect 24584 17002 24636 17008
rect 17696 16546 17908 16574
rect 1676 3596 1728 3602
rect 1676 3538 1728 3544
rect 572 3460 624 3466
rect 572 3402 624 3408
rect 584 480 612 3402
rect 1688 480 1716 3538
rect 17880 3534 17908 16546
rect 37292 3602 37320 20046
rect 39316 17649 39344 20060
rect 40696 17882 40724 20060
rect 42628 19242 42656 20060
rect 42616 19236 42668 19242
rect 42616 19178 42668 19184
rect 43916 17950 43944 20060
rect 43904 17944 43956 17950
rect 43904 17886 43956 17892
rect 40684 17876 40736 17882
rect 40684 17818 40736 17824
rect 39302 17640 39358 17649
rect 39302 17575 39358 17584
rect 45848 17406 45876 20060
rect 47136 17814 47164 20060
rect 47124 17808 47176 17814
rect 47124 17750 47176 17756
rect 49068 17746 49096 20060
rect 50264 17785 50292 20060
rect 50250 17776 50306 17785
rect 49056 17740 49108 17746
rect 50250 17711 50306 17720
rect 49056 17682 49108 17688
rect 45836 17400 45888 17406
rect 45836 17342 45888 17348
rect 52288 17202 52316 20060
rect 52472 20046 53498 20074
rect 52276 17196 52328 17202
rect 52276 17138 52328 17144
rect 37280 3596 37332 3602
rect 37280 3538 37332 3544
rect 17868 3528 17920 3534
rect 17868 3470 17920 3476
rect 52472 3466 52500 20046
rect 55416 17474 55444 20060
rect 56796 17474 56824 20060
rect 58636 17678 58664 20060
rect 58624 17672 58676 17678
rect 58624 17614 58676 17620
rect 59924 17610 59952 20060
rect 59912 17604 59964 17610
rect 59912 17546 59964 17552
rect 55404 17468 55456 17474
rect 55404 17410 55456 17416
rect 56784 17468 56836 17474
rect 56784 17410 56836 17416
rect 61856 17377 61884 20060
rect 63880 17678 63908 20060
rect 63868 17672 63920 17678
rect 63868 17614 63920 17620
rect 65168 17610 65196 20060
rect 66180 19310 66208 20567
rect 67640 20538 67692 20544
rect 66168 19304 66220 19310
rect 66168 19246 66220 19252
rect 65156 17604 65208 17610
rect 65156 17546 65208 17552
rect 61842 17368 61898 17377
rect 61842 17303 61898 17312
rect 68388 3466 68416 34303
rect 68480 32337 68508 536794
rect 68560 470620 68612 470626
rect 68560 470562 68612 470568
rect 68466 32328 68522 32337
rect 68466 32263 68522 32272
rect 68466 28928 68522 28937
rect 68466 28863 68522 28872
rect 68480 3602 68508 28863
rect 68572 22137 68600 470562
rect 68652 378208 68704 378214
rect 68652 378150 68704 378156
rect 68664 39137 68692 378150
rect 68650 39128 68706 39137
rect 68650 39063 68706 39072
rect 71056 31482 71084 700674
rect 71044 31476 71096 31482
rect 71044 31418 71096 31424
rect 68558 22128 68614 22137
rect 68558 22063 68614 22072
rect 72988 17950 73016 703520
rect 105464 700874 105492 703520
rect 105452 700868 105504 700874
rect 105452 700810 105504 700816
rect 137848 683114 137876 703520
rect 137756 683086 137876 683114
rect 96802 51368 96858 51377
rect 96802 51303 96858 51312
rect 136546 51368 136602 51377
rect 136546 51303 136602 51312
rect 96528 48340 96580 48346
rect 96528 48282 96580 48288
rect 96252 46980 96304 46986
rect 96252 46922 96304 46928
rect 91008 42016 91060 42022
rect 91006 41984 91008 41993
rect 95884 42016 95936 42022
rect 91060 41984 91062 41993
rect 95884 41958 95936 41964
rect 91006 41919 91062 41928
rect 88246 38448 88302 38457
rect 88246 38383 88302 38392
rect 88154 35456 88210 35465
rect 88154 35391 88210 35400
rect 88062 32464 88118 32473
rect 88062 32399 88118 32408
rect 87602 29472 87658 29481
rect 87602 29407 87658 29416
rect 87418 26480 87474 26489
rect 87418 26415 87474 26424
rect 87236 24812 87288 24818
rect 87236 24754 87288 24760
rect 87248 23497 87276 24754
rect 87234 23488 87290 23497
rect 87234 23423 87290 23432
rect 87432 20670 87460 26415
rect 87420 20664 87472 20670
rect 87420 20606 87472 20612
rect 87616 19242 87644 29407
rect 88076 19922 88104 32399
rect 88168 19990 88196 35391
rect 88156 19984 88208 19990
rect 88156 19926 88208 19932
rect 88064 19916 88116 19922
rect 88064 19858 88116 19864
rect 88260 19553 88288 38383
rect 95896 19854 95924 41958
rect 96264 39409 96292 46922
rect 96344 44192 96396 44198
rect 96344 44134 96396 44140
rect 96250 39400 96306 39409
rect 96250 39335 96306 39344
rect 96356 37913 96384 44134
rect 96540 40769 96568 48282
rect 96816 42265 96844 51303
rect 97446 49328 97502 49337
rect 97446 49263 97502 49272
rect 97460 48346 97488 49263
rect 97448 48340 97500 48346
rect 97448 48282 97500 48288
rect 97446 47288 97502 47297
rect 97446 47223 97502 47232
rect 97460 46986 97488 47223
rect 97448 46980 97500 46986
rect 97448 46922 97500 46928
rect 97446 45248 97502 45257
rect 97446 45183 97502 45192
rect 97460 44198 97488 45183
rect 97448 44192 97500 44198
rect 97448 44134 97500 44140
rect 97446 43208 97502 43217
rect 97446 43143 97502 43152
rect 96802 42256 96858 42265
rect 96802 42191 96858 42200
rect 96802 41168 96858 41177
rect 96802 41103 96858 41112
rect 96526 40760 96582 40769
rect 96526 40695 96582 40704
rect 96618 39128 96674 39137
rect 96618 39063 96674 39072
rect 96342 37904 96398 37913
rect 96342 37839 96398 37848
rect 96344 37188 96396 37194
rect 96344 37130 96396 37136
rect 96356 36417 96384 37130
rect 96342 36408 96398 36417
rect 96342 36343 96398 36352
rect 96632 33289 96660 39063
rect 96816 34785 96844 41103
rect 97460 37194 97488 43143
rect 136560 42401 136588 51303
rect 136730 48648 136786 48657
rect 136730 48583 136786 48592
rect 136638 47016 136694 47025
rect 136638 46951 136694 46960
rect 136546 42392 136602 42401
rect 136546 42327 136602 42336
rect 131028 42016 131080 42022
rect 131026 41984 131028 41993
rect 135904 42016 135956 42022
rect 131080 41984 131082 41993
rect 135904 41958 135956 41964
rect 131026 41919 131082 41928
rect 128266 38448 128322 38457
rect 128266 38383 128322 38392
rect 97448 37188 97500 37194
rect 97448 37130 97500 37136
rect 97446 37088 97502 37097
rect 97446 37023 97502 37032
rect 96894 35048 96950 35057
rect 96894 34983 96950 34992
rect 96802 34776 96858 34785
rect 96802 34711 96858 34720
rect 96618 33280 96674 33289
rect 96618 33215 96674 33224
rect 96344 32972 96396 32978
rect 96344 32914 96396 32920
rect 96356 31929 96384 32914
rect 96342 31920 96398 31929
rect 96342 31855 96398 31864
rect 96908 30297 96936 34983
rect 97460 32978 97488 37023
rect 128174 35456 128230 35465
rect 128174 35391 128230 35400
rect 97448 32972 97500 32978
rect 97448 32914 97500 32920
rect 97538 32736 97594 32745
rect 97538 32671 97594 32680
rect 97354 30968 97410 30977
rect 97354 30903 97410 30912
rect 96894 30288 96950 30297
rect 96894 30223 96950 30232
rect 96344 28960 96396 28966
rect 96342 28928 96344 28937
rect 96396 28928 96398 28937
rect 96342 28863 96398 28872
rect 96528 27668 96580 27674
rect 96528 27610 96580 27616
rect 96344 27464 96396 27470
rect 96342 27432 96344 27441
rect 96396 27432 96398 27441
rect 96342 27367 96398 27376
rect 96344 26580 96396 26586
rect 96344 26522 96396 26528
rect 96356 24449 96384 26522
rect 96540 25809 96568 27610
rect 97368 27470 97396 30903
rect 97552 28966 97580 32671
rect 127990 32464 128046 32473
rect 127990 32399 128046 32408
rect 127622 29472 127678 29481
rect 127622 29407 127678 29416
rect 97540 28960 97592 28966
rect 97446 28928 97502 28937
rect 97540 28902 97592 28908
rect 97446 28863 97502 28872
rect 97460 27674 97488 28863
rect 97448 27668 97500 27674
rect 97448 27610 97500 27616
rect 97356 27464 97408 27470
rect 97356 27406 97408 27412
rect 97446 26888 97502 26897
rect 97446 26823 97502 26832
rect 97460 26586 97488 26823
rect 97448 26580 97500 26586
rect 97448 26522 97500 26528
rect 127530 26480 127586 26489
rect 127530 26415 127586 26424
rect 96526 25800 96582 25809
rect 96526 25735 96582 25744
rect 97446 24848 97502 24857
rect 97446 24783 97502 24792
rect 96342 24440 96398 24449
rect 96342 24375 96398 24384
rect 97460 22982 97488 24783
rect 127070 23488 127126 23497
rect 127070 23423 127126 23432
rect 96344 22976 96396 22982
rect 96342 22944 96344 22953
rect 97448 22976 97500 22982
rect 96396 22944 96398 22953
rect 97448 22918 97500 22924
rect 96342 22879 96398 22888
rect 97446 22808 97502 22817
rect 97446 22743 97502 22752
rect 97460 21486 97488 22743
rect 96344 21480 96396 21486
rect 96342 21448 96344 21457
rect 97448 21480 97500 21486
rect 96396 21448 96398 21457
rect 97448 21422 97500 21428
rect 96342 21383 96398 21392
rect 126978 20496 127034 20505
rect 126978 20431 127034 20440
rect 126992 19854 127020 20431
rect 95884 19848 95936 19854
rect 95884 19790 95936 19796
rect 126980 19848 127032 19854
rect 126980 19790 127032 19796
rect 127084 19553 127112 23423
rect 127544 19990 127572 26415
rect 127532 19984 127584 19990
rect 127532 19926 127584 19932
rect 127636 19922 127664 29407
rect 127624 19916 127676 19922
rect 127624 19858 127676 19864
rect 88246 19544 88302 19553
rect 88246 19479 88302 19488
rect 127070 19544 127126 19553
rect 128004 19514 128032 32399
rect 127070 19479 127126 19488
rect 127992 19508 128044 19514
rect 127992 19450 128044 19456
rect 128188 19242 128216 35391
rect 128280 19582 128308 38383
rect 135916 30274 135944 41958
rect 136362 40488 136418 40497
rect 136362 40423 136418 40432
rect 136270 35048 136326 35057
rect 136270 34983 136326 34992
rect 136284 30433 136312 34983
rect 136376 34921 136404 40423
rect 136652 39409 136680 46951
rect 136744 40769 136772 48583
rect 136822 44568 136878 44577
rect 136822 44503 136878 44512
rect 136730 40760 136786 40769
rect 136730 40695 136786 40704
rect 136638 39400 136694 39409
rect 136638 39335 136694 39344
rect 136454 38720 136510 38729
rect 136454 38655 136510 38664
rect 136362 34912 136418 34921
rect 136362 34847 136418 34856
rect 136468 33425 136496 38655
rect 136836 37777 136864 44503
rect 136914 42936 136970 42945
rect 136914 42871 136970 42880
rect 136822 37768 136878 37777
rect 136822 37703 136878 37712
rect 136638 36544 136694 36553
rect 136638 36479 136694 36488
rect 136454 33416 136510 33425
rect 136454 33351 136510 33360
rect 136652 32450 136680 36479
rect 136928 36281 136956 42871
rect 136914 36272 136970 36281
rect 136914 36207 136970 36216
rect 136560 32422 136680 32450
rect 136560 31929 136588 32422
rect 136638 32328 136694 32337
rect 136638 32263 136694 32272
rect 136546 31920 136602 31929
rect 136546 31855 136602 31864
rect 136270 30424 136326 30433
rect 136270 30359 136326 30368
rect 135916 30246 136588 30274
rect 136454 28248 136510 28257
rect 136454 28183 136510 28192
rect 136270 26616 136326 26625
rect 136270 26551 136326 26560
rect 136284 24449 136312 26551
rect 136468 25945 136496 28183
rect 136454 25936 136510 25945
rect 136454 25871 136510 25880
rect 136270 24440 136326 24449
rect 136270 24375 136326 24384
rect 136454 24440 136510 24449
rect 136454 24375 136510 24384
rect 136468 22953 136496 24375
rect 136454 22944 136510 22953
rect 136454 22879 136510 22888
rect 136560 19961 136588 30246
rect 136652 28937 136680 32263
rect 136730 30424 136786 30433
rect 136730 30359 136786 30368
rect 136638 28928 136694 28937
rect 136638 28863 136694 28872
rect 136744 27305 136772 30359
rect 136730 27296 136786 27305
rect 136730 27231 136786 27240
rect 136546 19952 136602 19961
rect 136546 19887 136602 19896
rect 128268 19576 128320 19582
rect 128268 19518 128320 19524
rect 87604 19236 87656 19242
rect 87604 19178 87656 19184
rect 128176 19236 128228 19242
rect 128176 19178 128228 19184
rect 72976 17944 73028 17950
rect 72976 17886 73028 17892
rect 137756 17134 137784 683086
rect 169666 38448 169722 38457
rect 169666 38383 169722 38392
rect 169574 35456 169630 35465
rect 169574 35391 169630 35400
rect 169482 32464 169538 32473
rect 169482 32399 169538 32408
rect 169022 29472 169078 29481
rect 169022 29407 169078 29416
rect 168378 23488 168434 23497
rect 168378 23423 168434 23432
rect 168392 19582 168420 23423
rect 168380 19576 168432 19582
rect 168380 19518 168432 19524
rect 169036 19514 169064 29407
rect 169114 26480 169170 26489
rect 169114 26415 169170 26424
rect 169024 19508 169076 19514
rect 169024 19450 169076 19456
rect 169128 19242 169156 26415
rect 169496 19922 169524 32399
rect 169588 19990 169616 35391
rect 169576 19984 169628 19990
rect 169576 19926 169628 19932
rect 169484 19916 169536 19922
rect 169484 19858 169536 19864
rect 169680 19553 169708 38383
rect 169666 19544 169722 19553
rect 169666 19479 169722 19488
rect 169116 19236 169168 19242
rect 169116 19178 169168 19184
rect 170324 17202 170352 703520
rect 202800 700806 202828 703520
rect 202788 700800 202840 700806
rect 202788 700742 202840 700748
rect 235184 700670 235212 703520
rect 267660 700738 267688 703520
rect 267648 700732 267700 700738
rect 267648 700674 267700 700680
rect 235172 700664 235224 700670
rect 235172 700606 235224 700612
rect 300136 700534 300164 703520
rect 332520 700602 332548 703520
rect 332508 700596 332560 700602
rect 332508 700538 332560 700544
rect 300124 700528 300176 700534
rect 300124 700470 300176 700476
rect 364996 700466 365024 703520
rect 364984 700460 365036 700466
rect 364984 700402 365036 700408
rect 249064 52624 249116 52630
rect 249064 52566 249116 52572
rect 218058 51300 218114 51309
rect 218058 51235 218114 51244
rect 218072 51134 218100 51235
rect 176568 51128 176620 51134
rect 178132 51128 178184 51134
rect 176568 51070 176620 51076
rect 178130 51096 178132 51105
rect 216588 51128 216640 51134
rect 178184 51096 178186 51105
rect 176476 48340 176528 48346
rect 176476 48282 176528 48288
rect 176292 42832 176344 42838
rect 176292 42774 176344 42780
rect 171416 42016 171468 42022
rect 171414 41984 171416 41993
rect 175924 42016 175976 42022
rect 171468 41984 171470 41993
rect 175924 41958 175976 41964
rect 171414 41919 171470 41928
rect 175936 19854 175964 41958
rect 176304 36417 176332 42774
rect 176488 40905 176516 48282
rect 176580 42401 176608 51070
rect 216588 51070 216640 51076
rect 218060 51128 218112 51134
rect 218060 51070 218112 51076
rect 178130 51031 178186 51040
rect 178130 49056 178186 49065
rect 178130 48991 178186 49000
rect 178144 48346 178172 48991
rect 178132 48340 178184 48346
rect 178132 48282 178184 48288
rect 178038 47016 178094 47025
rect 178038 46951 178094 46960
rect 216496 46980 216548 46986
rect 177854 45248 177910 45257
rect 177854 45183 177910 45192
rect 176566 42392 176622 42401
rect 176566 42327 176622 42336
rect 176474 40896 176530 40905
rect 176474 40831 176530 40840
rect 176384 40112 176436 40118
rect 176384 40054 176436 40060
rect 176290 36408 176346 36417
rect 176290 36343 176346 36352
rect 176396 34921 176424 40054
rect 176568 39432 176620 39438
rect 176566 39400 176568 39409
rect 176620 39400 176622 39409
rect 176566 39335 176622 39344
rect 176476 38684 176528 38690
rect 176476 38626 176528 38632
rect 176382 34912 176438 34921
rect 176382 34847 176438 34856
rect 176488 33425 176516 38626
rect 177868 37942 177896 45183
rect 178052 39438 178080 46951
rect 216496 46922 216548 46928
rect 216404 43104 216456 43110
rect 216404 43046 216456 43052
rect 178130 42936 178186 42945
rect 178130 42871 178186 42880
rect 178144 42838 178172 42871
rect 178132 42832 178184 42838
rect 178132 42774 178184 42780
rect 209686 41440 209742 41449
rect 209686 41375 209742 41384
rect 178130 40896 178186 40905
rect 178130 40831 178186 40840
rect 178144 40118 178172 40831
rect 178132 40112 178184 40118
rect 178132 40054 178184 40060
rect 178040 39432 178092 39438
rect 178040 39374 178092 39380
rect 178130 38856 178186 38865
rect 178130 38791 178186 38800
rect 178144 38690 178172 38791
rect 178132 38684 178184 38690
rect 178132 38626 178184 38632
rect 209594 38448 209650 38457
rect 209594 38383 209650 38392
rect 176752 37936 176804 37942
rect 176750 37904 176752 37913
rect 177856 37936 177908 37942
rect 176804 37904 176806 37913
rect 177856 37878 177908 37884
rect 176750 37839 176806 37848
rect 178130 36816 178186 36825
rect 178130 36751 178186 36760
rect 177854 35048 177910 35057
rect 177854 34983 177910 34992
rect 177868 34542 177896 34983
rect 176752 34536 176804 34542
rect 176752 34478 176804 34484
rect 177856 34536 177908 34542
rect 177856 34478 177908 34484
rect 176474 33416 176530 33425
rect 176474 33351 176530 33360
rect 176568 31952 176620 31958
rect 176566 31920 176568 31929
rect 176620 31920 176622 31929
rect 176566 31855 176622 31864
rect 176764 30433 176792 34478
rect 178038 32736 178094 32745
rect 178038 32671 178094 32680
rect 176750 30424 176806 30433
rect 176750 30359 176806 30368
rect 178052 28966 178080 32671
rect 178144 31958 178172 36751
rect 209502 35456 209558 35465
rect 209502 35391 209558 35400
rect 209410 32464 209466 32473
rect 209410 32399 209466 32408
rect 178132 31952 178184 31958
rect 178132 31894 178184 31900
rect 178130 30696 178186 30705
rect 178130 30631 178186 30640
rect 176568 28960 176620 28966
rect 176566 28928 176568 28937
rect 178040 28960 178092 28966
rect 176620 28928 176622 28937
rect 176566 28863 176622 28872
rect 177854 28928 177910 28937
rect 178040 28902 178092 28908
rect 177854 28863 177910 28872
rect 177868 27674 177896 28863
rect 176752 27668 176804 27674
rect 176752 27610 176804 27616
rect 177856 27668 177908 27674
rect 177856 27610 177908 27616
rect 176568 27464 176620 27470
rect 176566 27432 176568 27441
rect 176620 27432 176622 27441
rect 176566 27367 176622 27376
rect 176764 25945 176792 27610
rect 178144 27470 178172 30631
rect 209042 29472 209098 29481
rect 209042 29407 209098 29416
rect 178132 27464 178184 27470
rect 178132 27406 178184 27412
rect 177854 26888 177910 26897
rect 177854 26823 177910 26832
rect 176750 25936 176806 25945
rect 176750 25871 176806 25880
rect 177868 24818 177896 26823
rect 208490 26480 208546 26489
rect 208490 26415 208546 26424
rect 176752 24812 176804 24818
rect 176752 24754 176804 24760
rect 177856 24812 177908 24818
rect 177856 24754 177908 24760
rect 176764 24449 176792 24754
rect 178130 24576 178186 24585
rect 178130 24511 178186 24520
rect 176750 24440 176806 24449
rect 176750 24375 176806 24384
rect 178144 22982 178172 24511
rect 176568 22976 176620 22982
rect 176566 22944 176568 22953
rect 178132 22976 178184 22982
rect 176620 22944 176622 22953
rect 178132 22918 178184 22924
rect 176566 22879 176622 22888
rect 178130 22536 178186 22545
rect 178130 22471 178186 22480
rect 178144 21486 178172 22471
rect 176568 21480 176620 21486
rect 176566 21448 176568 21457
rect 178132 21480 178184 21486
rect 176620 21448 176622 21457
rect 178132 21422 178184 21428
rect 176566 21383 176622 21392
rect 208398 20496 208454 20505
rect 208398 20431 208454 20440
rect 208412 19854 208440 20431
rect 208504 19990 208532 26415
rect 208582 23488 208638 23497
rect 208582 23423 208638 23432
rect 208492 19984 208544 19990
rect 208492 19926 208544 19932
rect 175924 19848 175976 19854
rect 175924 19790 175976 19796
rect 208400 19848 208452 19854
rect 208400 19790 208452 19796
rect 208596 19553 208624 23423
rect 209056 19922 209084 29407
rect 209044 19916 209096 19922
rect 209044 19858 209096 19864
rect 208582 19544 208638 19553
rect 208582 19479 208638 19488
rect 209424 19242 209452 32399
rect 209412 19236 209464 19242
rect 209412 19178 209464 19184
rect 209516 19038 209544 35391
rect 209608 19106 209636 38383
rect 209700 19174 209728 41375
rect 216416 36417 216444 43046
rect 216508 39409 216536 46922
rect 216600 42401 216628 51070
rect 218058 49260 218114 49269
rect 218058 49195 218114 49204
rect 218072 48346 218100 49195
rect 217324 48340 217376 48346
rect 217324 48282 217376 48288
rect 218060 48340 218112 48346
rect 218060 48282 218112 48288
rect 216586 42392 216642 42401
rect 216586 42327 216642 42336
rect 217336 40769 217364 48282
rect 218058 47220 218114 47229
rect 218058 47155 218114 47164
rect 218072 46986 218100 47155
rect 218060 46980 218112 46986
rect 218060 46922 218112 46928
rect 218058 45180 218114 45189
rect 218058 45115 218114 45124
rect 217966 43140 218022 43149
rect 217966 43075 217968 43084
rect 218020 43075 218022 43084
rect 217968 43046 218020 43052
rect 217506 41168 217562 41177
rect 217506 41103 217562 41112
rect 217322 40760 217378 40769
rect 217322 40695 217378 40704
rect 216494 39400 216550 39409
rect 216494 39335 216550 39344
rect 217414 39128 217470 39137
rect 217414 39063 217470 39072
rect 216588 37936 216640 37942
rect 216586 37904 216588 37913
rect 216640 37904 216642 37913
rect 216586 37839 216642 37848
rect 216402 36408 216458 36417
rect 216402 36343 216458 36352
rect 216864 34536 216916 34542
rect 216864 34478 216916 34484
rect 216496 32904 216548 32910
rect 216496 32846 216548 32852
rect 216508 28937 216536 32846
rect 216588 31952 216640 31958
rect 216586 31920 216588 31929
rect 216640 31920 216642 31929
rect 216586 31855 216642 31864
rect 216876 30433 216904 34478
rect 217428 33289 217456 39063
rect 217520 34785 217548 41103
rect 218072 37942 218100 45115
rect 249076 38457 249104 52566
rect 249156 52556 249208 52562
rect 249156 52498 249208 52504
rect 249168 41449 249196 52498
rect 287704 52488 287756 52494
rect 287704 52430 287756 52436
rect 258170 51368 258226 51377
rect 258170 51303 258226 51312
rect 257894 49192 257950 49201
rect 257894 49127 257950 49136
rect 257344 46980 257396 46986
rect 257344 46922 257396 46928
rect 257252 44192 257304 44198
rect 257252 44134 257304 44140
rect 257160 42696 257212 42702
rect 257160 42638 257212 42644
rect 257172 42401 257200 42638
rect 257158 42392 257214 42401
rect 257158 42327 257214 42336
rect 249154 41440 249210 41449
rect 249154 41375 249210 41384
rect 249062 38448 249118 38457
rect 249062 38383 249118 38392
rect 218060 37936 218112 37942
rect 257264 37913 257292 44134
rect 257356 39273 257384 46922
rect 257618 43072 257674 43081
rect 257618 43007 257674 43016
rect 257342 39264 257398 39273
rect 257342 39199 257398 39208
rect 218060 37878 218112 37884
rect 257250 37904 257306 37913
rect 257250 37839 257306 37848
rect 218058 37020 218114 37029
rect 218058 36955 218114 36964
rect 217966 34980 218022 34989
rect 217966 34915 218022 34924
rect 217506 34776 217562 34785
rect 217506 34711 217562 34720
rect 217980 34542 218008 34915
rect 217968 34536 218020 34542
rect 217968 34478 218020 34484
rect 217414 33280 217470 33289
rect 217414 33215 217470 33224
rect 217966 32940 218022 32949
rect 217966 32875 217968 32884
rect 218020 32875 218022 32884
rect 217968 32846 218020 32852
rect 218072 31958 218100 36955
rect 257632 36281 257660 43007
rect 257908 40769 257936 49127
rect 258184 42702 258212 51303
rect 258262 47220 258318 47229
rect 258262 47155 258318 47164
rect 258276 46986 258304 47155
rect 258264 46980 258316 46986
rect 258264 46922 258316 46928
rect 258262 45180 258318 45189
rect 258262 45115 258318 45124
rect 258276 44198 258304 45115
rect 258264 44192 258316 44198
rect 258264 44134 258316 44140
rect 258172 42696 258224 42702
rect 258172 42638 258224 42644
rect 257986 41032 258042 41041
rect 257986 40967 258042 40976
rect 257894 40760 257950 40769
rect 257894 40695 257950 40704
rect 258000 39114 258028 40967
rect 257908 39086 258028 39114
rect 257618 36272 257674 36281
rect 257618 36207 257674 36216
rect 257344 35964 257396 35970
rect 257344 35906 257396 35912
rect 257160 34536 257212 34542
rect 257160 34478 257212 34484
rect 218060 31952 218112 31958
rect 218060 31894 218112 31900
rect 218058 30900 218114 30909
rect 218058 30835 218114 30844
rect 216862 30424 216918 30433
rect 216862 30359 216918 30368
rect 216494 28928 216550 28937
rect 216494 28863 216550 28872
rect 217966 28860 218022 28869
rect 217966 28795 218022 28804
rect 216588 27464 216640 27470
rect 216586 27432 216588 27441
rect 216640 27432 216642 27441
rect 216586 27367 216642 27376
rect 216864 26580 216916 26586
rect 216864 26522 216916 26528
rect 216876 26058 216904 26522
rect 216784 26030 216904 26058
rect 216784 24449 216812 26030
rect 217980 25974 218008 28795
rect 218072 27470 218100 30835
rect 257172 30433 257200 34478
rect 257356 31793 257384 35906
rect 257908 34785 257936 39086
rect 257986 38992 258042 39001
rect 257986 38927 258042 38936
rect 257894 34776 257950 34785
rect 257894 34711 257950 34720
rect 258000 33289 258028 38927
rect 258262 37020 258318 37029
rect 258262 36955 258318 36964
rect 258276 35970 258304 36955
rect 258264 35964 258316 35970
rect 258264 35906 258316 35912
rect 258262 34980 258318 34989
rect 258262 34915 258318 34924
rect 258276 34542 258304 34915
rect 258264 34536 258316 34542
rect 258264 34478 258316 34484
rect 257986 33280 258042 33289
rect 257986 33215 258042 33224
rect 287716 33114 287744 52430
rect 366364 40724 366416 40730
rect 366364 40666 366416 40672
rect 287704 33108 287756 33114
rect 287704 33050 287756 33056
rect 257986 32872 258042 32881
rect 257986 32807 258042 32816
rect 257342 31784 257398 31793
rect 257342 31719 257398 31728
rect 257434 30832 257490 30841
rect 257434 30767 257490 30776
rect 257158 30424 257214 30433
rect 257158 30359 257214 30368
rect 249062 29472 249118 29481
rect 249062 29407 249118 29416
rect 218060 27464 218112 27470
rect 218060 27406 218112 27412
rect 218058 26820 218114 26829
rect 218058 26755 218114 26764
rect 218072 26586 218100 26755
rect 218060 26580 218112 26586
rect 218060 26522 218112 26528
rect 216864 25968 216916 25974
rect 216862 25936 216864 25945
rect 217968 25968 218020 25974
rect 216916 25936 216918 25945
rect 217968 25910 218020 25916
rect 216862 25871 216918 25880
rect 218058 24780 218114 24789
rect 218058 24715 218114 24724
rect 216770 24440 216826 24449
rect 216770 24375 216826 24384
rect 218072 22982 218100 24715
rect 248602 23488 248658 23497
rect 248602 23423 248658 23432
rect 216588 22976 216640 22982
rect 216586 22944 216588 22953
rect 218060 22976 218112 22982
rect 216640 22944 216642 22953
rect 218060 22918 218112 22924
rect 216586 22879 216642 22888
rect 218058 22740 218114 22749
rect 218058 22675 218114 22684
rect 218072 21486 218100 22675
rect 216588 21480 216640 21486
rect 216586 21448 216588 21457
rect 218060 21480 218112 21486
rect 216640 21448 216642 21457
rect 218060 21422 218112 21428
rect 216586 21383 216642 21392
rect 218058 20768 218114 20777
rect 216588 20732 216640 20738
rect 218058 20703 218060 20712
rect 216588 20674 216640 20680
rect 218112 20703 218114 20712
rect 218060 20674 218112 20680
rect 216600 20233 216628 20674
rect 216586 20224 216642 20233
rect 216586 20159 216642 20168
rect 209688 19168 209740 19174
rect 209688 19110 209740 19116
rect 248616 19106 248644 23423
rect 249076 19242 249104 29407
rect 257344 27668 257396 27674
rect 257344 27610 257396 27616
rect 249154 26480 249210 26489
rect 249154 26415 249210 26424
rect 249064 19236 249116 19242
rect 249064 19178 249116 19184
rect 209596 19100 209648 19106
rect 209596 19042 209648 19048
rect 248604 19100 248656 19106
rect 248604 19042 248656 19048
rect 249168 19038 249196 26415
rect 257160 26308 257212 26314
rect 257160 26250 257212 26256
rect 257172 24449 257200 26250
rect 257356 25809 257384 27610
rect 257448 27305 257476 30767
rect 258000 28801 258028 32807
rect 258262 28860 258318 28869
rect 257986 28792 258042 28801
rect 258262 28795 258318 28804
rect 257986 28727 258042 28736
rect 258276 27674 258304 28795
rect 258264 27668 258316 27674
rect 258264 27610 258316 27616
rect 257434 27296 257490 27305
rect 257434 27231 257490 27240
rect 258262 26820 258318 26829
rect 258262 26755 258318 26764
rect 258276 26314 258304 26755
rect 258264 26308 258316 26314
rect 258264 26250 258316 26256
rect 257342 25800 257398 25809
rect 257342 25735 257398 25744
rect 288348 25560 288400 25566
rect 288348 25502 288400 25508
rect 258262 24780 258318 24789
rect 258262 24715 258318 24724
rect 257158 24440 257214 24449
rect 257158 24375 257214 24384
rect 258276 23866 258304 24715
rect 257160 23860 257212 23866
rect 257160 23802 257212 23808
rect 258264 23860 258316 23866
rect 258264 23802 258316 23808
rect 257172 22953 257200 23802
rect 257158 22944 257214 22953
rect 257158 22879 257214 22888
rect 258262 22740 258318 22749
rect 258262 22675 258318 22684
rect 258276 22166 258304 22675
rect 257160 22160 257212 22166
rect 257160 22102 257212 22108
rect 258264 22160 258316 22166
rect 258264 22102 258316 22108
rect 257172 21457 257200 22102
rect 257158 21448 257214 21457
rect 257158 21383 257214 21392
rect 249706 20496 249762 20505
rect 249706 20431 249762 20440
rect 249720 19174 249748 20431
rect 288360 19310 288388 25502
rect 288348 19304 288400 19310
rect 288348 19246 288400 19252
rect 249708 19168 249760 19174
rect 249708 19110 249760 19116
rect 209504 19032 209556 19038
rect 209504 18974 209556 18980
rect 249156 19032 249208 19038
rect 249156 18974 249208 18980
rect 366376 17270 366404 40666
rect 397472 17338 397500 703520
rect 429856 17406 429884 703520
rect 462332 700398 462360 703520
rect 462320 700392 462372 700398
rect 462320 700334 462372 700340
rect 494808 700330 494836 703520
rect 494796 700324 494848 700330
rect 494796 700266 494848 700272
rect 527192 17542 527220 703520
rect 527180 17536 527232 17542
rect 527180 17478 527232 17484
rect 559668 17474 559696 703520
rect 580170 697232 580226 697241
rect 580170 697167 580226 697176
rect 580184 696998 580212 697167
rect 580172 696992 580224 696998
rect 580172 696934 580224 696940
rect 580262 670712 580318 670721
rect 580262 670647 580318 670656
rect 580170 591016 580226 591025
rect 580170 590951 580226 590960
rect 580184 590714 580212 590951
rect 580172 590708 580224 590714
rect 580172 590650 580224 590656
rect 580170 564360 580226 564369
rect 580170 564295 580226 564304
rect 580184 563106 580212 564295
rect 580172 563100 580224 563106
rect 580172 563042 580224 563048
rect 580170 537840 580226 537849
rect 580170 537775 580226 537784
rect 580184 536858 580212 537775
rect 580172 536852 580224 536858
rect 580172 536794 580224 536800
rect 580170 511320 580226 511329
rect 580170 511255 580226 511264
rect 580184 510678 580212 511255
rect 580172 510672 580224 510678
rect 580172 510614 580224 510620
rect 579986 471472 580042 471481
rect 579986 471407 580042 471416
rect 580000 470626 580028 471407
rect 579988 470620 580040 470626
rect 579988 470562 580040 470568
rect 579618 431624 579674 431633
rect 579618 431559 579674 431568
rect 579632 430642 579660 431559
rect 579620 430636 579672 430642
rect 579620 430578 579672 430584
rect 580170 404968 580226 404977
rect 580170 404903 580226 404912
rect 580184 404394 580212 404903
rect 580172 404388 580224 404394
rect 580172 404330 580224 404336
rect 580170 378448 580226 378457
rect 580170 378383 580226 378392
rect 580184 378214 580212 378383
rect 580172 378208 580224 378214
rect 580172 378150 580224 378156
rect 579802 232384 579858 232393
rect 579802 232319 579858 232328
rect 579816 231878 579844 232319
rect 579804 231872 579856 231878
rect 579804 231814 579856 231820
rect 580170 192536 580226 192545
rect 580170 192471 580226 192480
rect 580184 191894 580212 192471
rect 580172 191888 580224 191894
rect 580172 191830 580224 191836
rect 579986 152688 580042 152697
rect 579986 152623 580042 152632
rect 580000 151842 580028 152623
rect 579988 151836 580040 151842
rect 579988 151778 580040 151784
rect 580170 33144 580226 33153
rect 580170 33079 580172 33088
rect 580224 33079 580226 33088
rect 580172 33050 580224 33056
rect 580276 17610 580304 670647
rect 580354 644056 580410 644065
rect 580354 643991 580410 644000
rect 580368 17746 580396 643991
rect 580446 617536 580502 617545
rect 580446 617471 580502 617480
rect 580356 17740 580408 17746
rect 580356 17682 580408 17688
rect 580460 17678 580488 617471
rect 580538 484664 580594 484673
rect 580538 484599 580594 484608
rect 580552 17882 580580 484599
rect 580630 351928 580686 351937
rect 580630 351863 580686 351872
rect 580540 17876 580592 17882
rect 580540 17818 580592 17824
rect 580644 17814 580672 351863
rect 580722 272232 580778 272241
rect 580722 272167 580778 272176
rect 580632 17808 580684 17814
rect 580632 17750 580684 17756
rect 580448 17672 580500 17678
rect 580448 17614 580500 17620
rect 580264 17604 580316 17610
rect 580264 17546 580316 17552
rect 559656 17468 559708 17474
rect 559656 17410 559708 17416
rect 429844 17400 429896 17406
rect 429844 17342 429896 17348
rect 397460 17332 397512 17338
rect 397460 17274 397512 17280
rect 366364 17264 366416 17270
rect 366364 17206 366416 17212
rect 170312 17196 170364 17202
rect 170312 17138 170364 17144
rect 137744 17128 137796 17134
rect 137744 17070 137796 17076
rect 580736 17066 580764 272167
rect 580814 112840 580870 112849
rect 580814 112775 580870 112784
rect 580828 25566 580856 112775
rect 580906 72992 580962 73001
rect 580906 72927 580962 72936
rect 580920 40730 580948 72927
rect 580908 40724 580960 40730
rect 580908 40666 580960 40672
rect 580816 25560 580868 25566
rect 580816 25502 580868 25508
rect 580724 17060 580776 17066
rect 580724 17002 580776 17008
rect 68468 3596 68520 3602
rect 68468 3538 68520 3544
rect 125876 3596 125928 3602
rect 125876 3538 125928 3544
rect 52460 3460 52512 3466
rect 52460 3402 52512 3408
rect 68376 3460 68428 3466
rect 68376 3402 68428 3408
rect 125888 480 125916 3538
rect 129372 3528 129424 3534
rect 129372 3470 129424 3476
rect 132958 3496 133014 3505
rect 126980 3460 127032 3466
rect 126980 3402 127032 3408
rect 126992 480 127020 3402
rect 129384 480 129412 3470
rect 132958 3431 133014 3440
rect 132972 480 133000 3431
rect 136454 3360 136510 3369
rect 136454 3295 136510 3304
rect 136468 480 136496 3295
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9926 -960 10038 480
rect 11122 -960 11234 480
rect 12318 -960 12430 480
rect 13514 -960 13626 480
rect 14710 -960 14822 480
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 18206 -960 18318 480
rect 19402 -960 19514 480
rect 20598 -960 20710 480
rect 21794 -960 21906 480
rect 22990 -960 23102 480
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26486 -960 26598 480
rect 27682 -960 27794 480
rect 28878 -960 28990 480
rect 30074 -960 30186 480
rect 31270 -960 31382 480
rect 32374 -960 32486 480
rect 33570 -960 33682 480
rect 34766 -960 34878 480
rect 35962 -960 36074 480
rect 37158 -960 37270 480
rect 38354 -960 38466 480
rect 39550 -960 39662 480
rect 40654 -960 40766 480
rect 41850 -960 41962 480
rect 43046 -960 43158 480
rect 44242 -960 44354 480
rect 45438 -960 45550 480
rect 46634 -960 46746 480
rect 47830 -960 47942 480
rect 48934 -960 49046 480
rect 50130 -960 50242 480
rect 51326 -960 51438 480
rect 52522 -960 52634 480
rect 53718 -960 53830 480
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 57214 -960 57326 480
rect 58410 -960 58522 480
rect 59606 -960 59718 480
rect 60802 -960 60914 480
rect 61998 -960 62110 480
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65494 -960 65606 480
rect 66690 -960 66802 480
rect 67886 -960 67998 480
rect 69082 -960 69194 480
rect 70278 -960 70390 480
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73774 -960 73886 480
rect 74970 -960 75082 480
rect 76166 -960 76278 480
rect 77362 -960 77474 480
rect 78558 -960 78670 480
rect 79662 -960 79774 480
rect 80858 -960 80970 480
rect 82054 -960 82166 480
rect 83250 -960 83362 480
rect 84446 -960 84558 480
rect 85642 -960 85754 480
rect 86838 -960 86950 480
rect 87942 -960 88054 480
rect 89138 -960 89250 480
rect 90334 -960 90446 480
rect 91530 -960 91642 480
rect 92726 -960 92838 480
rect 93922 -960 94034 480
rect 95118 -960 95230 480
rect 96222 -960 96334 480
rect 97418 -960 97530 480
rect 98614 -960 98726 480
rect 99810 -960 99922 480
rect 101006 -960 101118 480
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104502 -960 104614 480
rect 105698 -960 105810 480
rect 106894 -960 107006 480
rect 108090 -960 108202 480
rect 109286 -960 109398 480
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112782 -960 112894 480
rect 113978 -960 114090 480
rect 115174 -960 115286 480
rect 116370 -960 116482 480
rect 117566 -960 117678 480
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 121062 -960 121174 480
rect 122258 -960 122370 480
rect 123454 -960 123566 480
rect 124650 -960 124762 480
rect 125846 -960 125958 480
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 129342 -960 129454 480
rect 130538 -960 130650 480
rect 131734 -960 131846 480
rect 132930 -960 133042 480
rect 134126 -960 134238 480
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137622 -960 137734 480
rect 138818 -960 138930 480
rect 140014 -960 140126 480
rect 141210 -960 141322 480
rect 142406 -960 142518 480
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145902 -960 146014 480
rect 147098 -960 147210 480
rect 148294 -960 148406 480
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 154182 -960 154294 480
rect 155378 -960 155490 480
rect 156574 -960 156686 480
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162462 -960 162574 480
rect 163658 -960 163770 480
rect 164854 -960 164966 480
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170742 -960 170854 480
rect 171938 -960 172050 480
rect 173134 -960 173246 480
rect 174238 -960 174350 480
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 179022 -960 179134 480
rect 180218 -960 180330 480
rect 181414 -960 181526 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 187302 -960 187414 480
rect 188498 -960 188610 480
rect 189694 -960 189806 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 199078 -960 199190 480
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207358 -960 207470 480
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 212142 -960 212254 480
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215638 -960 215750 480
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 220422 -960 220534 480
rect 221526 -960 221638 480
rect 222722 -960 222834 480
rect 223918 -960 224030 480
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228702 -960 228814 480
rect 229806 -960 229918 480
rect 231002 -960 231114 480
rect 232198 -960 232310 480
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236982 -960 237094 480
rect 238086 -960 238198 480
rect 239282 -960 239394 480
rect 240478 -960 240590 480
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 246366 -960 246478 480
rect 247562 -960 247674 480
rect 248758 -960 248870 480
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254646 -960 254758 480
rect 255842 -960 255954 480
rect 257038 -960 257150 480
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262926 -960 263038 480
rect 264122 -960 264234 480
rect 265318 -960 265430 480
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268814 -960 268926 480
rect 270010 -960 270122 480
rect 271206 -960 271318 480
rect 272402 -960 272514 480
rect 273598 -960 273710 480
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 277094 -960 277206 480
rect 278290 -960 278402 480
rect 279486 -960 279598 480
rect 280682 -960 280794 480
rect 281878 -960 281990 480
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 285374 -960 285486 480
rect 286570 -960 286682 480
rect 287766 -960 287878 480
rect 288962 -960 289074 480
rect 290158 -960 290270 480
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293654 -960 293766 480
rect 294850 -960 294962 480
rect 296046 -960 296158 480
rect 297242 -960 297354 480
rect 298438 -960 298550 480
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301934 -960 302046 480
rect 303130 -960 303242 480
rect 304326 -960 304438 480
rect 305522 -960 305634 480
rect 306718 -960 306830 480
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 310214 -960 310326 480
rect 311410 -960 311522 480
rect 312606 -960 312718 480
rect 313802 -960 313914 480
rect 314998 -960 315110 480
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318494 -960 318606 480
rect 319690 -960 319802 480
rect 320886 -960 320998 480
rect 322082 -960 322194 480
rect 323278 -960 323390 480
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326774 -960 326886 480
rect 327970 -960 328082 480
rect 329166 -960 329278 480
rect 330362 -960 330474 480
rect 331558 -960 331670 480
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 335054 -960 335166 480
rect 336250 -960 336362 480
rect 337446 -960 337558 480
rect 338642 -960 338754 480
rect 339838 -960 339950 480
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 343334 -960 343446 480
rect 344530 -960 344642 480
rect 345726 -960 345838 480
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351614 -960 351726 480
rect 352810 -960 352922 480
rect 354006 -960 354118 480
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 -960 358810 480
rect 359894 -960 360006 480
rect 361090 -960 361202 480
rect 362286 -960 362398 480
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 368174 -960 368286 480
rect 369370 -960 369482 480
rect 370566 -960 370678 480
rect 371670 -960 371782 480
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376454 -960 376566 480
rect 377650 -960 377762 480
rect 378846 -960 378958 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384734 -960 384846 480
rect 385930 -960 386042 480
rect 387126 -960 387238 480
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396510 -960 396622 480
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404790 -960 404902 480
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409574 -960 409686 480
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 413070 -960 413182 480
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 417854 -960 417966 480
rect 418958 -960 419070 480
rect 420154 -960 420266 480
rect 421350 -960 421462 480
rect 422546 -960 422658 480
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 426134 -960 426246 480
rect 427238 -960 427350 480
rect 428434 -960 428546 480
rect 429630 -960 429742 480
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 433218 -960 433330 480
rect 434414 -960 434526 480
rect 435518 -960 435630 480
rect 436714 -960 436826 480
rect 437910 -960 438022 480
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443798 -960 443910 480
rect 444994 -960 445106 480
rect 446190 -960 446302 480
rect 447386 -960 447498 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 452078 -960 452190 480
rect 453274 -960 453386 480
rect 454470 -960 454582 480
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 460358 -960 460470 480
rect 461554 -960 461666 480
rect 462750 -960 462862 480
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 466246 -960 466358 480
rect 467442 -960 467554 480
rect 468638 -960 468750 480
rect 469834 -960 469946 480
rect 471030 -960 471142 480
rect 472226 -960 472338 480
rect 473422 -960 473534 480
rect 474526 -960 474638 480
rect 475722 -960 475834 480
rect 476918 -960 477030 480
rect 478114 -960 478226 480
rect 479310 -960 479422 480
rect 480506 -960 480618 480
rect 481702 -960 481814 480
rect 482806 -960 482918 480
rect 484002 -960 484114 480
rect 485198 -960 485310 480
rect 486394 -960 486506 480
rect 487590 -960 487702 480
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 491086 -960 491198 480
rect 492282 -960 492394 480
rect 493478 -960 493590 480
rect 494674 -960 494786 480
rect 495870 -960 495982 480
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 499366 -960 499478 480
rect 500562 -960 500674 480
rect 501758 -960 501870 480
rect 502954 -960 503066 480
rect 504150 -960 504262 480
rect 505346 -960 505458 480
rect 506450 -960 506562 480
rect 507646 -960 507758 480
rect 508842 -960 508954 480
rect 510038 -960 510150 480
rect 511234 -960 511346 480
rect 512430 -960 512542 480
rect 513534 -960 513646 480
rect 514730 -960 514842 480
rect 515926 -960 516038 480
rect 517122 -960 517234 480
rect 518318 -960 518430 480
rect 519514 -960 519626 480
rect 520710 -960 520822 480
rect 521814 -960 521926 480
rect 523010 -960 523122 480
rect 524206 -960 524318 480
rect 525402 -960 525514 480
rect 526598 -960 526710 480
rect 527794 -960 527906 480
rect 528990 -960 529102 480
rect 530094 -960 530206 480
rect 531290 -960 531402 480
rect 532486 -960 532598 480
rect 533682 -960 533794 480
rect 534878 -960 534990 480
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538374 -960 538486 480
rect 539570 -960 539682 480
rect 540766 -960 540878 480
rect 541962 -960 542074 480
rect 543158 -960 543270 480
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546654 -960 546766 480
rect 547850 -960 547962 480
rect 549046 -960 549158 480
rect 550242 -960 550354 480
rect 551438 -960 551550 480
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554934 -960 555046 480
rect 556130 -960 556242 480
rect 557326 -960 557438 480
rect 558522 -960 558634 480
rect 559718 -960 559830 480
rect 560822 -960 560934 480
rect 562018 -960 562130 480
rect 563214 -960 563326 480
rect 564410 -960 564522 480
rect 565606 -960 565718 480
rect 566802 -960 566914 480
rect 567998 -960 568110 480
rect 569102 -960 569214 480
rect 570298 -960 570410 480
rect 571494 -960 571606 480
rect 572690 -960 572802 480
rect 573886 -960 573998 480
rect 575082 -960 575194 480
rect 576278 -960 576390 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 3422 684256 3478 684312
rect 3330 553832 3386 553888
rect 2778 527856 2834 527912
rect 3146 449520 3202 449576
rect 3330 358400 3386 358456
rect 3330 345344 3386 345400
rect 3330 293120 3386 293176
rect 3330 254088 3386 254144
rect 3330 201864 3386 201920
rect 3330 136720 3386 136776
rect 3330 84632 3386 84688
rect 3238 58520 3294 58576
rect 2962 45464 3018 45520
rect 3514 658144 3570 658200
rect 3514 632068 3516 632088
rect 3516 632068 3568 632088
rect 3568 632068 3570 632088
rect 3514 632032 3570 632068
rect 3514 410488 3570 410544
rect 3238 19352 3294 19408
rect 3606 397432 3662 397488
rect 3698 306176 3754 306232
rect 3790 241032 3846 241088
rect 3882 188808 3938 188864
rect 3974 149776 4030 149832
rect 4066 97552 4122 97608
rect 16486 37848 16542 37904
rect 43994 39344 44050 39400
rect 47306 39344 47362 39400
rect 54574 39344 54630 39400
rect 60554 39208 60610 39264
rect 17866 37032 17922 37088
rect 65338 38256 65394 38312
rect 17866 34992 17922 35048
rect 17774 33632 17830 33688
rect 17590 31592 17646 31648
rect 17774 30232 17830 30288
rect 17682 28192 17738 28248
rect 15842 24112 15898 24168
rect 17866 26832 17922 26888
rect 17866 24812 17922 24848
rect 17866 24792 17868 24812
rect 17868 24792 17920 24812
rect 17920 24792 17922 24812
rect 67730 30912 67786 30968
rect 68374 35672 68430 35728
rect 68374 34312 68430 34368
rect 68282 27512 68338 27568
rect 67638 25472 67694 25528
rect 65338 24656 65394 24712
rect 17774 21392 17830 21448
rect 21638 20576 21694 20632
rect 66166 20576 66222 20632
rect 32862 17448 32918 17504
rect 39302 17584 39358 17640
rect 50250 17720 50306 17776
rect 61842 17312 61898 17368
rect 68466 32272 68522 32328
rect 68466 28872 68522 28928
rect 68650 39072 68706 39128
rect 68558 22072 68614 22128
rect 96802 51312 96858 51368
rect 136546 51312 136602 51368
rect 91006 41964 91008 41984
rect 91008 41964 91060 41984
rect 91060 41964 91062 41984
rect 91006 41928 91062 41964
rect 88246 38392 88302 38448
rect 88154 35400 88210 35456
rect 88062 32408 88118 32464
rect 87602 29416 87658 29472
rect 87418 26424 87474 26480
rect 87234 23432 87290 23488
rect 96250 39344 96306 39400
rect 97446 49272 97502 49328
rect 97446 47232 97502 47288
rect 97446 45192 97502 45248
rect 97446 43152 97502 43208
rect 96802 42200 96858 42256
rect 96802 41112 96858 41168
rect 96526 40704 96582 40760
rect 96618 39072 96674 39128
rect 96342 37848 96398 37904
rect 96342 36352 96398 36408
rect 136730 48592 136786 48648
rect 136638 46960 136694 47016
rect 136546 42336 136602 42392
rect 131026 41964 131028 41984
rect 131028 41964 131080 41984
rect 131080 41964 131082 41984
rect 131026 41928 131082 41964
rect 128266 38392 128322 38448
rect 97446 37032 97502 37088
rect 96894 34992 96950 35048
rect 96802 34720 96858 34776
rect 96618 33224 96674 33280
rect 96342 31864 96398 31920
rect 128174 35400 128230 35456
rect 97538 32680 97594 32736
rect 97354 30912 97410 30968
rect 96894 30232 96950 30288
rect 96342 28908 96344 28928
rect 96344 28908 96396 28928
rect 96396 28908 96398 28928
rect 96342 28872 96398 28908
rect 96342 27412 96344 27432
rect 96344 27412 96396 27432
rect 96396 27412 96398 27432
rect 96342 27376 96398 27412
rect 127990 32408 128046 32464
rect 127622 29416 127678 29472
rect 97446 28872 97502 28928
rect 97446 26832 97502 26888
rect 127530 26424 127586 26480
rect 96526 25744 96582 25800
rect 97446 24792 97502 24848
rect 96342 24384 96398 24440
rect 127070 23432 127126 23488
rect 96342 22924 96344 22944
rect 96344 22924 96396 22944
rect 96396 22924 96398 22944
rect 96342 22888 96398 22924
rect 97446 22752 97502 22808
rect 96342 21428 96344 21448
rect 96344 21428 96396 21448
rect 96396 21428 96398 21448
rect 96342 21392 96398 21428
rect 126978 20440 127034 20496
rect 88246 19488 88302 19544
rect 127070 19488 127126 19544
rect 136362 40432 136418 40488
rect 136270 34992 136326 35048
rect 136822 44512 136878 44568
rect 136730 40704 136786 40760
rect 136638 39344 136694 39400
rect 136454 38664 136510 38720
rect 136362 34856 136418 34912
rect 136914 42880 136970 42936
rect 136822 37712 136878 37768
rect 136638 36488 136694 36544
rect 136454 33360 136510 33416
rect 136914 36216 136970 36272
rect 136638 32272 136694 32328
rect 136546 31864 136602 31920
rect 136270 30368 136326 30424
rect 136454 28192 136510 28248
rect 136270 26560 136326 26616
rect 136454 25880 136510 25936
rect 136270 24384 136326 24440
rect 136454 24384 136510 24440
rect 136454 22888 136510 22944
rect 136730 30368 136786 30424
rect 136638 28872 136694 28928
rect 136730 27240 136786 27296
rect 136546 19896 136602 19952
rect 169666 38392 169722 38448
rect 169574 35400 169630 35456
rect 169482 32408 169538 32464
rect 169022 29416 169078 29472
rect 168378 23432 168434 23488
rect 169114 26424 169170 26480
rect 169666 19488 169722 19544
rect 218058 51244 218114 51300
rect 178130 51076 178132 51096
rect 178132 51076 178184 51096
rect 178184 51076 178186 51096
rect 171414 41964 171416 41984
rect 171416 41964 171468 41984
rect 171468 41964 171470 41984
rect 171414 41928 171470 41964
rect 178130 51040 178186 51076
rect 178130 49000 178186 49056
rect 178038 46960 178094 47016
rect 177854 45192 177910 45248
rect 176566 42336 176622 42392
rect 176474 40840 176530 40896
rect 176290 36352 176346 36408
rect 176566 39380 176568 39400
rect 176568 39380 176620 39400
rect 176620 39380 176622 39400
rect 176566 39344 176622 39380
rect 176382 34856 176438 34912
rect 178130 42880 178186 42936
rect 209686 41384 209742 41440
rect 178130 40840 178186 40896
rect 178130 38800 178186 38856
rect 209594 38392 209650 38448
rect 176750 37884 176752 37904
rect 176752 37884 176804 37904
rect 176804 37884 176806 37904
rect 176750 37848 176806 37884
rect 178130 36760 178186 36816
rect 177854 34992 177910 35048
rect 176474 33360 176530 33416
rect 176566 31900 176568 31920
rect 176568 31900 176620 31920
rect 176620 31900 176622 31920
rect 176566 31864 176622 31900
rect 178038 32680 178094 32736
rect 176750 30368 176806 30424
rect 209502 35400 209558 35456
rect 209410 32408 209466 32464
rect 178130 30640 178186 30696
rect 176566 28908 176568 28928
rect 176568 28908 176620 28928
rect 176620 28908 176622 28928
rect 176566 28872 176622 28908
rect 177854 28872 177910 28928
rect 176566 27412 176568 27432
rect 176568 27412 176620 27432
rect 176620 27412 176622 27432
rect 176566 27376 176622 27412
rect 209042 29416 209098 29472
rect 177854 26832 177910 26888
rect 176750 25880 176806 25936
rect 208490 26424 208546 26480
rect 178130 24520 178186 24576
rect 176750 24384 176806 24440
rect 176566 22924 176568 22944
rect 176568 22924 176620 22944
rect 176620 22924 176622 22944
rect 176566 22888 176622 22924
rect 178130 22480 178186 22536
rect 176566 21428 176568 21448
rect 176568 21428 176620 21448
rect 176620 21428 176622 21448
rect 176566 21392 176622 21428
rect 208398 20440 208454 20496
rect 208582 23432 208638 23488
rect 208582 19488 208638 19544
rect 218058 49204 218114 49260
rect 216586 42336 216642 42392
rect 218058 47164 218114 47220
rect 218058 45124 218114 45180
rect 217966 43104 218022 43140
rect 217966 43084 217968 43104
rect 217968 43084 218020 43104
rect 218020 43084 218022 43104
rect 217506 41112 217562 41168
rect 217322 40704 217378 40760
rect 216494 39344 216550 39400
rect 217414 39072 217470 39128
rect 216586 37884 216588 37904
rect 216588 37884 216640 37904
rect 216640 37884 216642 37904
rect 216586 37848 216642 37884
rect 216402 36352 216458 36408
rect 216586 31900 216588 31920
rect 216588 31900 216640 31920
rect 216640 31900 216642 31920
rect 216586 31864 216642 31900
rect 258170 51312 258226 51368
rect 257894 49136 257950 49192
rect 257158 42336 257214 42392
rect 249154 41384 249210 41440
rect 249062 38392 249118 38448
rect 257618 43016 257674 43072
rect 257342 39208 257398 39264
rect 257250 37848 257306 37904
rect 218058 36964 218114 37020
rect 217966 34924 218022 34980
rect 217506 34720 217562 34776
rect 217414 33224 217470 33280
rect 217966 32904 218022 32940
rect 217966 32884 217968 32904
rect 217968 32884 218020 32904
rect 218020 32884 218022 32904
rect 258262 47164 258318 47220
rect 258262 45124 258318 45180
rect 257986 40976 258042 41032
rect 257894 40704 257950 40760
rect 257618 36216 257674 36272
rect 218058 30844 218114 30900
rect 216862 30368 216918 30424
rect 216494 28872 216550 28928
rect 217966 28804 218022 28860
rect 216586 27412 216588 27432
rect 216588 27412 216640 27432
rect 216640 27412 216642 27432
rect 216586 27376 216642 27412
rect 257986 38936 258042 38992
rect 257894 34720 257950 34776
rect 258262 36964 258318 37020
rect 258262 34924 258318 34980
rect 257986 33224 258042 33280
rect 257986 32816 258042 32872
rect 257342 31728 257398 31784
rect 257434 30776 257490 30832
rect 257158 30368 257214 30424
rect 249062 29416 249118 29472
rect 218058 26764 218114 26820
rect 216862 25916 216864 25936
rect 216864 25916 216916 25936
rect 216916 25916 216918 25936
rect 216862 25880 216918 25916
rect 218058 24724 218114 24780
rect 216770 24384 216826 24440
rect 248602 23432 248658 23488
rect 216586 22924 216588 22944
rect 216588 22924 216640 22944
rect 216640 22924 216642 22944
rect 216586 22888 216642 22924
rect 218058 22684 218114 22740
rect 216586 21428 216588 21448
rect 216588 21428 216640 21448
rect 216640 21428 216642 21448
rect 216586 21392 216642 21428
rect 218058 20732 218114 20768
rect 218058 20712 218060 20732
rect 218060 20712 218112 20732
rect 218112 20712 218114 20732
rect 216586 20168 216642 20224
rect 249154 26424 249210 26480
rect 258262 28804 258318 28860
rect 257986 28736 258042 28792
rect 257434 27240 257490 27296
rect 258262 26764 258318 26820
rect 257342 25744 257398 25800
rect 258262 24724 258318 24780
rect 257158 24384 257214 24440
rect 257158 22888 257214 22944
rect 258262 22684 258318 22740
rect 257158 21392 257214 21448
rect 249706 20440 249762 20496
rect 580170 697176 580226 697232
rect 580262 670656 580318 670712
rect 580170 590960 580226 591016
rect 580170 564304 580226 564360
rect 580170 537784 580226 537840
rect 580170 511264 580226 511320
rect 579986 471416 580042 471472
rect 579618 431568 579674 431624
rect 580170 404912 580226 404968
rect 580170 378392 580226 378448
rect 579802 232328 579858 232384
rect 580170 192480 580226 192536
rect 579986 152632 580042 152688
rect 580170 33108 580226 33144
rect 580170 33088 580172 33108
rect 580172 33088 580224 33108
rect 580224 33088 580226 33108
rect 580354 644000 580410 644056
rect 580446 617480 580502 617536
rect 580538 484608 580594 484664
rect 580630 351872 580686 351928
rect 580722 272176 580778 272232
rect 580814 112784 580870 112840
rect 580906 72936 580962 72992
rect 132958 3440 133014 3496
rect 136454 3304 136510 3360
<< metal3 >>
rect -960 697220 480 697460
rect 580165 697234 580231 697237
rect 583520 697234 584960 697324
rect 580165 697232 584960 697234
rect 580165 697176 580170 697232
rect 580226 697176 584960 697232
rect 580165 697174 584960 697176
rect 580165 697171 580231 697174
rect 583520 697084 584960 697174
rect -960 684314 480 684404
rect 3417 684314 3483 684317
rect -960 684312 3483 684314
rect -960 684256 3422 684312
rect 3478 684256 3483 684312
rect -960 684254 3483 684256
rect -960 684164 480 684254
rect 3417 684251 3483 684254
rect 583520 683756 584960 683996
rect -960 671108 480 671348
rect 580257 670714 580323 670717
rect 583520 670714 584960 670804
rect 580257 670712 584960 670714
rect 580257 670656 580262 670712
rect 580318 670656 584960 670712
rect 580257 670654 584960 670656
rect 580257 670651 580323 670654
rect 583520 670564 584960 670654
rect -960 658202 480 658292
rect 3509 658202 3575 658205
rect -960 658200 3575 658202
rect -960 658144 3514 658200
rect 3570 658144 3575 658200
rect -960 658142 3575 658144
rect -960 658052 480 658142
rect 3509 658139 3575 658142
rect 583520 657236 584960 657476
rect -960 644996 480 645236
rect 580349 644058 580415 644061
rect 583520 644058 584960 644148
rect 580349 644056 584960 644058
rect 580349 644000 580354 644056
rect 580410 644000 584960 644056
rect 580349 643998 584960 644000
rect 580349 643995 580415 643998
rect 583520 643908 584960 643998
rect -960 632090 480 632180
rect 3509 632090 3575 632093
rect -960 632088 3575 632090
rect -960 632032 3514 632088
rect 3570 632032 3575 632088
rect -960 632030 3575 632032
rect -960 631940 480 632030
rect 3509 632027 3575 632030
rect 583520 630716 584960 630956
rect -960 619020 480 619260
rect 580441 617538 580507 617541
rect 583520 617538 584960 617628
rect 580441 617536 584960 617538
rect 580441 617480 580446 617536
rect 580502 617480 584960 617536
rect 580441 617478 584960 617480
rect 580441 617475 580507 617478
rect 583520 617388 584960 617478
rect -960 606114 480 606204
rect 3366 606114 3372 606116
rect -960 606054 3372 606114
rect -960 605964 480 606054
rect 3366 606052 3372 606054
rect 3436 606052 3442 606116
rect 583520 604060 584960 604300
rect -960 592908 480 593148
rect 580165 591018 580231 591021
rect 583520 591018 584960 591108
rect 580165 591016 584960 591018
rect 580165 590960 580170 591016
rect 580226 590960 584960 591016
rect 580165 590958 584960 590960
rect 580165 590955 580231 590958
rect 583520 590868 584960 590958
rect -960 580002 480 580092
rect 3550 580002 3556 580004
rect -960 579942 3556 580002
rect -960 579852 480 579942
rect 3550 579940 3556 579942
rect 3620 579940 3626 580004
rect 583520 577540 584960 577780
rect -960 566796 480 567036
rect 580165 564362 580231 564365
rect 583520 564362 584960 564452
rect 580165 564360 584960 564362
rect 580165 564304 580170 564360
rect 580226 564304 584960 564360
rect 580165 564302 584960 564304
rect 580165 564299 580231 564302
rect 583520 564212 584960 564302
rect -960 553890 480 553980
rect 3325 553890 3391 553893
rect -960 553888 3391 553890
rect -960 553832 3330 553888
rect 3386 553832 3391 553888
rect -960 553830 3391 553832
rect -960 553740 480 553830
rect 3325 553827 3391 553830
rect 583520 551020 584960 551260
rect -960 540684 480 540924
rect 580165 537842 580231 537845
rect 583520 537842 584960 537932
rect 580165 537840 584960 537842
rect 580165 537784 580170 537840
rect 580226 537784 584960 537840
rect 580165 537782 584960 537784
rect 580165 537779 580231 537782
rect 583520 537692 584960 537782
rect -960 527914 480 528004
rect 2773 527914 2839 527917
rect -960 527912 2839 527914
rect -960 527856 2778 527912
rect 2834 527856 2839 527912
rect -960 527854 2839 527856
rect -960 527764 480 527854
rect 2773 527851 2839 527854
rect 583520 524364 584960 524604
rect -960 514708 480 514948
rect 580165 511322 580231 511325
rect 583520 511322 584960 511412
rect 580165 511320 584960 511322
rect 580165 511264 580170 511320
rect 580226 511264 584960 511320
rect 580165 511262 584960 511264
rect 580165 511259 580231 511262
rect 583520 511172 584960 511262
rect -960 501802 480 501892
rect 3734 501802 3740 501804
rect -960 501742 3740 501802
rect -960 501652 480 501742
rect 3734 501740 3740 501742
rect 3804 501740 3810 501804
rect 583520 497844 584960 498084
rect -960 488596 480 488836
rect 580533 484666 580599 484669
rect 583520 484666 584960 484756
rect 580533 484664 584960 484666
rect 580533 484608 580538 484664
rect 580594 484608 584960 484664
rect 580533 484606 584960 484608
rect 580533 484603 580599 484606
rect 583520 484516 584960 484606
rect -960 475690 480 475780
rect 3918 475690 3924 475692
rect -960 475630 3924 475690
rect -960 475540 480 475630
rect 3918 475628 3924 475630
rect 3988 475628 3994 475692
rect 579981 471474 580047 471477
rect 583520 471474 584960 471564
rect 579981 471472 584960 471474
rect 579981 471416 579986 471472
rect 580042 471416 584960 471472
rect 579981 471414 584960 471416
rect 579981 471411 580047 471414
rect 583520 471324 584960 471414
rect -960 462484 480 462724
rect 583520 457996 584960 458236
rect -960 449578 480 449668
rect 3141 449578 3207 449581
rect -960 449576 3207 449578
rect -960 449520 3146 449576
rect 3202 449520 3207 449576
rect -960 449518 3207 449520
rect -960 449428 480 449518
rect 3141 449515 3207 449518
rect 583520 444668 584960 444908
rect -960 436508 480 436748
rect 579613 431626 579679 431629
rect 583520 431626 584960 431716
rect 579613 431624 584960 431626
rect 579613 431568 579618 431624
rect 579674 431568 584960 431624
rect 579613 431566 584960 431568
rect 579613 431563 579679 431566
rect 583520 431476 584960 431566
rect -960 423452 480 423692
rect 583520 418148 584960 418388
rect -960 410546 480 410636
rect 3509 410546 3575 410549
rect -960 410544 3575 410546
rect -960 410488 3514 410544
rect 3570 410488 3575 410544
rect -960 410486 3575 410488
rect -960 410396 480 410486
rect 3509 410483 3575 410486
rect 580165 404970 580231 404973
rect 583520 404970 584960 405060
rect 580165 404968 584960 404970
rect 580165 404912 580170 404968
rect 580226 404912 584960 404968
rect 580165 404910 584960 404912
rect 580165 404907 580231 404910
rect 583520 404820 584960 404910
rect -960 397490 480 397580
rect 3601 397490 3667 397493
rect -960 397488 3667 397490
rect -960 397432 3606 397488
rect 3662 397432 3667 397488
rect -960 397430 3667 397432
rect -960 397340 480 397430
rect 3601 397427 3667 397430
rect 583520 391628 584960 391868
rect -960 384284 480 384524
rect 580165 378450 580231 378453
rect 583520 378450 584960 378540
rect 580165 378448 584960 378450
rect 580165 378392 580170 378448
rect 580226 378392 584960 378448
rect 580165 378390 584960 378392
rect 580165 378387 580231 378390
rect 583520 378300 584960 378390
rect -960 371228 480 371468
rect 583520 364972 584960 365212
rect -960 358458 480 358548
rect 3325 358458 3391 358461
rect -960 358456 3391 358458
rect -960 358400 3330 358456
rect 3386 358400 3391 358456
rect -960 358398 3391 358400
rect -960 358308 480 358398
rect 3325 358395 3391 358398
rect 580625 351930 580691 351933
rect 583520 351930 584960 352020
rect 580625 351928 584960 351930
rect 580625 351872 580630 351928
rect 580686 351872 584960 351928
rect 580625 351870 584960 351872
rect 580625 351867 580691 351870
rect 583520 351780 584960 351870
rect -960 345402 480 345492
rect 3325 345402 3391 345405
rect -960 345400 3391 345402
rect -960 345344 3330 345400
rect 3386 345344 3391 345400
rect -960 345342 3391 345344
rect -960 345252 480 345342
rect 3325 345339 3391 345342
rect 583520 338452 584960 338692
rect -960 332196 480 332436
rect 21950 325212 21956 325276
rect 22020 325274 22026 325276
rect 583520 325274 584960 325364
rect 22020 325214 584960 325274
rect 22020 325212 22026 325214
rect 583520 325124 584960 325214
rect -960 319140 480 319380
rect 583520 311932 584960 312172
rect -960 306234 480 306324
rect 3693 306234 3759 306237
rect -960 306232 3759 306234
rect -960 306176 3698 306232
rect 3754 306176 3759 306232
rect -960 306174 3759 306176
rect -960 306084 480 306174
rect 3693 306171 3759 306174
rect 583520 298604 584960 298844
rect -960 293178 480 293268
rect 3325 293178 3391 293181
rect -960 293176 3391 293178
rect -960 293120 3330 293176
rect 3386 293120 3391 293176
rect -960 293118 3391 293120
rect -960 293028 480 293118
rect 3325 293115 3391 293118
rect 583520 285276 584960 285516
rect -960 279972 480 280212
rect 580717 272234 580783 272237
rect 583520 272234 584960 272324
rect 580717 272232 584960 272234
rect 580717 272176 580722 272232
rect 580778 272176 584960 272232
rect 580717 272174 584960 272176
rect 580717 272171 580783 272174
rect 583520 272084 584960 272174
rect -960 267052 480 267292
rect 583520 258756 584960 258996
rect -960 254146 480 254236
rect 3325 254146 3391 254149
rect -960 254144 3391 254146
rect -960 254088 3330 254144
rect 3386 254088 3391 254144
rect -960 254086 3391 254088
rect -960 253996 480 254086
rect 3325 254083 3391 254086
rect 583520 245428 584960 245668
rect -960 241090 480 241180
rect 3785 241090 3851 241093
rect -960 241088 3851 241090
rect -960 241032 3790 241088
rect 3846 241032 3851 241088
rect -960 241030 3851 241032
rect -960 240940 480 241030
rect 3785 241027 3851 241030
rect 579797 232386 579863 232389
rect 583520 232386 584960 232476
rect 579797 232384 584960 232386
rect 579797 232328 579802 232384
rect 579858 232328 584960 232384
rect 579797 232326 584960 232328
rect 579797 232323 579863 232326
rect 583520 232236 584960 232326
rect -960 227884 480 228124
rect 583520 218908 584960 219148
rect -960 214828 480 215068
rect 583520 205580 584960 205820
rect -960 201922 480 202012
rect 3325 201922 3391 201925
rect -960 201920 3391 201922
rect -960 201864 3330 201920
rect 3386 201864 3391 201920
rect -960 201862 3391 201864
rect -960 201772 480 201862
rect 3325 201859 3391 201862
rect 580165 192538 580231 192541
rect 583520 192538 584960 192628
rect 580165 192536 584960 192538
rect 580165 192480 580170 192536
rect 580226 192480 584960 192536
rect 580165 192478 584960 192480
rect 580165 192475 580231 192478
rect 583520 192388 584960 192478
rect -960 188866 480 188956
rect 3877 188866 3943 188869
rect -960 188864 3943 188866
rect -960 188808 3882 188864
rect 3938 188808 3943 188864
rect -960 188806 3943 188808
rect -960 188716 480 188806
rect 3877 188803 3943 188806
rect 583520 179060 584960 179300
rect -960 175796 480 176036
rect 583520 165732 584960 165972
rect -960 162740 480 162980
rect 579981 152690 580047 152693
rect 583520 152690 584960 152780
rect 579981 152688 584960 152690
rect 579981 152632 579986 152688
rect 580042 152632 584960 152688
rect 579981 152630 584960 152632
rect 579981 152627 580047 152630
rect 583520 152540 584960 152630
rect -960 149834 480 149924
rect 3969 149834 4035 149837
rect -960 149832 4035 149834
rect -960 149776 3974 149832
rect 4030 149776 4035 149832
rect -960 149774 4035 149776
rect -960 149684 480 149774
rect 3969 149771 4035 149774
rect 583520 139212 584960 139452
rect -960 136778 480 136868
rect 3325 136778 3391 136781
rect -960 136776 3391 136778
rect -960 136720 3330 136776
rect 3386 136720 3391 136776
rect -960 136718 3391 136720
rect -960 136628 480 136718
rect 3325 136715 3391 136718
rect 583520 125884 584960 126124
rect -960 123572 480 123812
rect 580809 112842 580875 112845
rect 583520 112842 584960 112932
rect 580809 112840 584960 112842
rect 580809 112784 580814 112840
rect 580870 112784 584960 112840
rect 580809 112782 584960 112784
rect 580809 112779 580875 112782
rect 583520 112692 584960 112782
rect -960 110516 480 110756
rect 583520 99364 584960 99604
rect -960 97610 480 97700
rect 4061 97610 4127 97613
rect -960 97608 4127 97610
rect -960 97552 4066 97608
rect 4122 97552 4127 97608
rect -960 97550 4127 97552
rect -960 97460 480 97550
rect 4061 97547 4127 97550
rect 583520 86036 584960 86276
rect -960 84690 480 84780
rect 3325 84690 3391 84693
rect -960 84688 3391 84690
rect -960 84632 3330 84688
rect 3386 84632 3391 84688
rect -960 84630 3391 84632
rect -960 84540 480 84630
rect 3325 84627 3391 84630
rect 580901 72994 580967 72997
rect 583520 72994 584960 73084
rect 580901 72992 584960 72994
rect 580901 72936 580906 72992
rect 580962 72936 584960 72992
rect 580901 72934 584960 72936
rect 580901 72931 580967 72934
rect 583520 72844 584960 72934
rect -960 71484 480 71724
rect 583520 59516 584960 59756
rect -960 58578 480 58668
rect 3233 58578 3299 58581
rect -960 58576 3299 58578
rect -960 58520 3238 58576
rect 3294 58520 3299 58576
rect -960 58518 3299 58520
rect -960 58428 480 58518
rect 3233 58515 3299 58518
rect 96797 51370 96863 51373
rect 136541 51370 136607 51373
rect 258165 51370 258231 51373
rect 96797 51368 97704 51370
rect 96797 51312 96802 51368
rect 96858 51312 97704 51368
rect 96797 51310 97704 51312
rect 136541 51368 137908 51370
rect 136541 51312 136546 51368
rect 136602 51312 137908 51368
rect 136541 51310 137908 51312
rect 258165 51368 258520 51370
rect 258165 51312 258170 51368
rect 258226 51312 258520 51368
rect 258165 51310 258520 51312
rect 96797 51307 96863 51310
rect 136541 51307 136607 51310
rect 258165 51307 258231 51310
rect 218053 51302 218119 51305
rect 218053 51300 218316 51302
rect 178174 51101 178234 51272
rect 218053 51244 218058 51300
rect 218114 51244 218316 51300
rect 218053 51242 218316 51244
rect 218053 51239 218119 51242
rect 178125 51096 178234 51101
rect 178125 51040 178130 51096
rect 178186 51040 178234 51096
rect 178125 51038 178234 51040
rect 178125 51035 178191 51038
rect 97441 49330 97507 49333
rect 97441 49328 97704 49330
rect 97441 49272 97446 49328
rect 97502 49272 97704 49328
rect 97441 49270 97704 49272
rect 97441 49267 97507 49270
rect 218053 49262 218119 49265
rect 218053 49260 218316 49262
rect 136725 48650 136791 48653
rect 137878 48650 137938 49232
rect 178174 49061 178234 49232
rect 218053 49204 218058 49260
rect 218114 49204 218316 49260
rect 218053 49202 218316 49204
rect 258030 49202 258520 49262
rect 218053 49199 218119 49202
rect 257889 49194 257955 49197
rect 258030 49194 258090 49202
rect 257889 49192 258090 49194
rect 257889 49136 257894 49192
rect 257950 49136 258090 49192
rect 257889 49134 258090 49136
rect 257889 49131 257955 49134
rect 178125 49056 178234 49061
rect 178125 49000 178130 49056
rect 178186 49000 178234 49056
rect 178125 48998 178234 49000
rect 178125 48995 178191 48998
rect 136725 48648 137938 48650
rect 136725 48592 136730 48648
rect 136786 48592 137938 48648
rect 136725 48590 137938 48592
rect 136725 48587 136791 48590
rect 97441 47290 97507 47293
rect 97441 47288 97704 47290
rect 97441 47232 97446 47288
rect 97502 47232 97704 47288
rect 97441 47230 97704 47232
rect 97441 47227 97507 47230
rect 136633 47018 136699 47021
rect 137878 47018 137938 47192
rect 178082 47021 178142 47260
rect 218053 47222 218119 47225
rect 258257 47222 258323 47225
rect 218053 47220 218316 47222
rect 218053 47164 218058 47220
rect 218114 47164 218316 47220
rect 218053 47162 218316 47164
rect 258257 47220 258520 47222
rect 258257 47164 258262 47220
rect 258318 47164 258520 47220
rect 258257 47162 258520 47164
rect 218053 47159 218119 47162
rect 258257 47159 258323 47162
rect 136633 47016 137938 47018
rect 136633 46960 136638 47016
rect 136694 46960 137938 47016
rect 136633 46958 137938 46960
rect 178033 47016 178142 47021
rect 178033 46960 178038 47016
rect 178094 46960 178142 47016
rect 178033 46958 178142 46960
rect 136633 46955 136699 46958
rect 178033 46955 178099 46958
rect 583520 46188 584960 46428
rect -960 45522 480 45612
rect 2957 45522 3023 45525
rect -960 45520 3023 45522
rect -960 45464 2962 45520
rect 3018 45464 3023 45520
rect -960 45462 3023 45464
rect -960 45372 480 45462
rect 2957 45459 3023 45462
rect 97441 45250 97507 45253
rect 177849 45250 177915 45253
rect 97441 45248 97704 45250
rect 97441 45192 97446 45248
rect 97502 45192 97704 45248
rect 97441 45190 97704 45192
rect 177849 45248 178112 45250
rect 177849 45192 177854 45248
rect 177910 45192 178112 45248
rect 177849 45190 178112 45192
rect 97441 45187 97507 45190
rect 177849 45187 177915 45190
rect 218053 45182 218119 45185
rect 258257 45182 258323 45185
rect 218053 45180 218316 45182
rect 136817 44570 136883 44573
rect 137878 44570 137938 45152
rect 218053 45124 218058 45180
rect 218114 45124 218316 45180
rect 218053 45122 218316 45124
rect 258257 45180 258520 45182
rect 258257 45124 258262 45180
rect 258318 45124 258520 45180
rect 258257 45122 258520 45124
rect 218053 45119 218119 45122
rect 258257 45119 258323 45122
rect 136817 44568 137938 44570
rect 136817 44512 136822 44568
rect 136878 44512 137938 44568
rect 136817 44510 137938 44512
rect 136817 44507 136883 44510
rect 97441 43210 97507 43213
rect 97441 43208 97704 43210
rect 97441 43152 97446 43208
rect 97502 43152 97704 43208
rect 97441 43150 97704 43152
rect 97441 43147 97507 43150
rect 217961 43142 218027 43145
rect 217961 43140 218316 43142
rect 136909 42938 136975 42941
rect 137878 42938 137938 43112
rect 178174 42941 178234 43112
rect 217961 43084 217966 43140
rect 218022 43084 218316 43140
rect 217961 43082 218316 43084
rect 258030 43082 258520 43142
rect 217961 43079 218027 43082
rect 257613 43074 257679 43077
rect 258030 43074 258090 43082
rect 257613 43072 258090 43074
rect 257613 43016 257618 43072
rect 257674 43016 258090 43072
rect 257613 43014 258090 43016
rect 257613 43011 257679 43014
rect 136909 42936 137938 42938
rect 136909 42880 136914 42936
rect 136970 42880 137938 42936
rect 136909 42878 137938 42880
rect 178125 42936 178234 42941
rect 178125 42880 178130 42936
rect 178186 42880 178234 42936
rect 178125 42878 178234 42880
rect 136909 42875 136975 42878
rect 178125 42875 178191 42878
rect 136541 42394 136607 42397
rect 176561 42394 176627 42397
rect 136406 42392 136607 42394
rect 136406 42336 136546 42392
rect 136602 42336 136607 42392
rect 136406 42334 136607 42336
rect 96797 42258 96863 42261
rect 96324 42256 96863 42258
rect 96324 42200 96802 42256
rect 96858 42200 96863 42256
rect 136406 42228 136466 42334
rect 136541 42331 136607 42334
rect 176518 42392 176627 42394
rect 176518 42336 176566 42392
rect 176622 42336 176627 42392
rect 176518 42331 176627 42336
rect 216581 42394 216647 42397
rect 257153 42394 257219 42397
rect 216581 42392 216690 42394
rect 216581 42336 216586 42392
rect 216642 42336 216690 42392
rect 216581 42331 216690 42336
rect 176518 42228 176578 42331
rect 216630 42228 216690 42331
rect 257110 42392 257219 42394
rect 257110 42336 257158 42392
rect 257214 42336 257219 42392
rect 257110 42331 257219 42336
rect 257110 42228 257170 42331
rect 96324 42198 96863 42200
rect 96797 42195 96863 42198
rect 91001 41986 91067 41989
rect 90958 41984 91067 41986
rect 90958 41928 91006 41984
rect 91062 41928 91067 41984
rect 90958 41923 91067 41928
rect 131021 41986 131087 41989
rect 171409 41986 171475 41989
rect 131021 41984 131130 41986
rect 131021 41928 131026 41984
rect 131082 41928 131130 41984
rect 131021 41923 131130 41928
rect 90958 41412 91018 41923
rect 131070 41412 131130 41923
rect 171366 41984 171475 41986
rect 171366 41928 171414 41984
rect 171470 41928 171475 41984
rect 171366 41923 171475 41928
rect 171366 41412 171426 41923
rect 209681 41442 209747 41445
rect 249149 41442 249215 41445
rect 209681 41440 211140 41442
rect 209681 41384 209686 41440
rect 209742 41384 211140 41440
rect 209681 41382 211140 41384
rect 249149 41440 251252 41442
rect 249149 41384 249154 41440
rect 249210 41384 251252 41440
rect 249149 41382 251252 41384
rect 209681 41379 209747 41382
rect 249149 41379 249215 41382
rect 96797 41170 96863 41173
rect 217501 41170 217567 41173
rect 96797 41168 97704 41170
rect 96797 41112 96802 41168
rect 96858 41112 97704 41168
rect 96797 41110 97704 41112
rect 217501 41168 218316 41170
rect 217501 41112 217506 41168
rect 217562 41112 218316 41168
rect 217501 41110 218316 41112
rect 96797 41107 96863 41110
rect 217501 41107 217567 41110
rect 96521 40762 96587 40765
rect 136725 40762 136791 40765
rect 96324 40760 96587 40762
rect 96324 40704 96526 40760
rect 96582 40704 96587 40760
rect 96324 40702 96587 40704
rect 136436 40760 136791 40762
rect 136436 40704 136730 40760
rect 136786 40704 136791 40760
rect 136436 40702 136791 40704
rect 96521 40699 96587 40702
rect 136725 40699 136791 40702
rect 136357 40490 136423 40493
rect 137878 40490 137938 41072
rect 178174 40901 178234 41072
rect 258030 41042 258520 41102
rect 258030 41037 258090 41042
rect 257981 41032 258090 41037
rect 257981 40976 257986 41032
rect 258042 40976 258090 41032
rect 257981 40974 258090 40976
rect 257981 40971 258047 40974
rect 176469 40898 176535 40901
rect 176469 40896 176578 40898
rect 176469 40840 176474 40896
rect 176530 40840 176578 40896
rect 176469 40835 176578 40840
rect 178125 40896 178234 40901
rect 178125 40840 178130 40896
rect 178186 40840 178234 40896
rect 178125 40838 178234 40840
rect 178125 40835 178191 40838
rect 176518 40732 176578 40835
rect 217317 40762 217383 40765
rect 257889 40762 257955 40765
rect 216844 40760 217383 40762
rect 216844 40704 217322 40760
rect 217378 40704 217383 40760
rect 216844 40702 217383 40704
rect 257140 40760 257955 40762
rect 257140 40704 257894 40760
rect 257950 40704 257955 40760
rect 257140 40702 257955 40704
rect 217317 40699 217383 40702
rect 257889 40699 257955 40702
rect 136357 40488 137938 40490
rect 136357 40432 136362 40488
rect 136418 40432 137938 40488
rect 136357 40430 137938 40432
rect 136357 40427 136423 40430
rect 43989 39404 44055 39405
rect 43989 39400 44036 39404
rect 44100 39402 44106 39404
rect 43989 39344 43994 39400
rect 43989 39340 44036 39344
rect 44100 39342 44146 39402
rect 44100 39340 44106 39342
rect 46974 39340 46980 39404
rect 47044 39402 47050 39404
rect 47301 39402 47367 39405
rect 47044 39400 47367 39402
rect 47044 39344 47306 39400
rect 47362 39344 47367 39400
rect 47044 39342 47367 39344
rect 47044 39340 47050 39342
rect 43989 39339 44055 39340
rect 47301 39339 47367 39342
rect 54569 39402 54635 39405
rect 55070 39402 55076 39404
rect 54569 39400 55076 39402
rect 54569 39344 54574 39400
rect 54630 39344 55076 39400
rect 54569 39342 55076 39344
rect 54569 39339 54635 39342
rect 55070 39340 55076 39342
rect 55140 39340 55146 39404
rect 96245 39402 96311 39405
rect 136633 39402 136699 39405
rect 176561 39402 176627 39405
rect 216489 39402 216555 39405
rect 96245 39400 96354 39402
rect 96245 39344 96250 39400
rect 96306 39344 96354 39400
rect 96245 39339 96354 39344
rect 60549 39268 60615 39269
rect 60549 39264 60596 39268
rect 60660 39266 60666 39268
rect 60549 39208 60554 39264
rect 60549 39204 60596 39208
rect 60660 39206 60706 39266
rect 96294 39236 96354 39339
rect 136406 39400 136699 39402
rect 136406 39344 136638 39400
rect 136694 39344 136699 39400
rect 136406 39342 136699 39344
rect 136406 39236 136466 39342
rect 136633 39339 136699 39342
rect 176518 39400 176627 39402
rect 176518 39344 176566 39400
rect 176622 39344 176627 39400
rect 176518 39339 176627 39344
rect 216446 39400 216555 39402
rect 216446 39344 216494 39400
rect 216550 39344 216555 39400
rect 216446 39339 216555 39344
rect 176518 39236 176578 39339
rect 216446 39236 216506 39339
rect 257337 39266 257403 39269
rect 257140 39264 257403 39266
rect 257140 39208 257342 39264
rect 257398 39208 257403 39264
rect 257140 39206 257403 39208
rect 60660 39204 60666 39206
rect 60549 39203 60615 39204
rect 257337 39203 257403 39206
rect 68645 39130 68711 39133
rect 65964 39128 68711 39130
rect 65964 39072 68650 39128
rect 68706 39072 68711 39128
rect 65964 39070 68711 39072
rect 68645 39067 68711 39070
rect 96613 39130 96679 39133
rect 217409 39130 217475 39133
rect 96613 39128 97704 39130
rect 96613 39072 96618 39128
rect 96674 39072 97704 39128
rect 96613 39070 97704 39072
rect 217409 39128 218316 39130
rect 217409 39072 217414 39128
rect 217470 39072 218316 39128
rect 217409 39070 218316 39072
rect 96613 39067 96679 39070
rect 217409 39067 217475 39070
rect 136449 38722 136515 38725
rect 137878 38722 137938 39032
rect 178174 38861 178234 39032
rect 258030 39002 258520 39062
rect 258030 38997 258090 39002
rect 257981 38992 258090 38997
rect 257981 38936 257986 38992
rect 258042 38936 258090 38992
rect 257981 38934 258090 38936
rect 257981 38931 258047 38934
rect 178125 38856 178234 38861
rect 178125 38800 178130 38856
rect 178186 38800 178234 38856
rect 178125 38798 178234 38800
rect 178125 38795 178191 38798
rect 136449 38720 137938 38722
rect 136449 38664 136454 38720
rect 136510 38664 137938 38720
rect 136449 38662 137938 38664
rect 136449 38659 136515 38662
rect 88241 38450 88307 38453
rect 128261 38450 128327 38453
rect 169661 38450 169727 38453
rect 209589 38450 209655 38453
rect 249057 38450 249123 38453
rect 88241 38448 90436 38450
rect 16481 37906 16547 37909
rect 20118 37906 20178 38420
rect 88241 38392 88246 38448
rect 88302 38392 90436 38448
rect 88241 38390 90436 38392
rect 128261 38448 130732 38450
rect 128261 38392 128266 38448
rect 128322 38392 130732 38448
rect 128261 38390 130732 38392
rect 169661 38448 170844 38450
rect 169661 38392 169666 38448
rect 169722 38392 170844 38448
rect 169661 38390 170844 38392
rect 209589 38448 211140 38450
rect 209589 38392 209594 38448
rect 209650 38392 211140 38448
rect 209589 38390 211140 38392
rect 249057 38448 251252 38450
rect 249057 38392 249062 38448
rect 249118 38392 251252 38448
rect 249057 38390 251252 38392
rect 88241 38387 88307 38390
rect 128261 38387 128327 38390
rect 169661 38387 169727 38390
rect 209589 38387 209655 38390
rect 249057 38387 249123 38390
rect 65333 38314 65399 38317
rect 65333 38312 65442 38314
rect 65333 38256 65338 38312
rect 65394 38256 65442 38312
rect 65333 38251 65442 38256
rect 16481 37904 20178 37906
rect 16481 37848 16486 37904
rect 16542 37848 20178 37904
rect 16481 37846 20178 37848
rect 16481 37843 16547 37846
rect 65382 37740 65442 38251
rect 96337 37906 96403 37909
rect 176745 37906 176811 37909
rect 96294 37904 96403 37906
rect 96294 37848 96342 37904
rect 96398 37848 96403 37904
rect 96294 37843 96403 37848
rect 176702 37904 176811 37906
rect 176702 37848 176750 37904
rect 176806 37848 176811 37904
rect 176702 37843 176811 37848
rect 216581 37906 216647 37909
rect 257245 37906 257311 37909
rect 216581 37904 216690 37906
rect 216581 37848 216586 37904
rect 216642 37848 216690 37904
rect 216581 37843 216690 37848
rect 96294 37740 96354 37843
rect 136817 37770 136883 37773
rect 136436 37768 136883 37770
rect 136436 37712 136822 37768
rect 136878 37712 136883 37768
rect 176702 37740 176762 37843
rect 216630 37740 216690 37843
rect 257110 37904 257311 37906
rect 257110 37848 257250 37904
rect 257306 37848 257311 37904
rect 257110 37846 257311 37848
rect 257110 37740 257170 37846
rect 257245 37843 257311 37846
rect 136436 37710 136883 37712
rect 136817 37707 136883 37710
rect 17861 37090 17927 37093
rect 97441 37090 97507 37093
rect 17861 37088 20148 37090
rect 17861 37032 17866 37088
rect 17922 37032 20148 37088
rect 17861 37030 20148 37032
rect 97441 37088 97704 37090
rect 97441 37032 97446 37088
rect 97502 37032 97704 37088
rect 97441 37030 97704 37032
rect 17861 37027 17927 37030
rect 97441 37027 97507 37030
rect 218053 37022 218119 37025
rect 258257 37022 258323 37025
rect 218053 37020 218316 37022
rect 136633 36546 136699 36549
rect 137878 36546 137938 36992
rect 178174 36821 178234 36992
rect 218053 36964 218058 37020
rect 218114 36964 218316 37020
rect 218053 36962 218316 36964
rect 258257 37020 258520 37022
rect 258257 36964 258262 37020
rect 258318 36964 258520 37020
rect 258257 36962 258520 36964
rect 218053 36959 218119 36962
rect 258257 36959 258323 36962
rect 178125 36816 178234 36821
rect 178125 36760 178130 36816
rect 178186 36760 178234 36816
rect 178125 36758 178234 36760
rect 178125 36755 178191 36758
rect 136633 36544 137938 36546
rect 136633 36488 136638 36544
rect 136694 36488 137938 36544
rect 136633 36486 137938 36488
rect 136633 36483 136699 36486
rect 96337 36410 96403 36413
rect 96294 36408 96403 36410
rect 96294 36352 96342 36408
rect 96398 36352 96403 36408
rect 96294 36347 96403 36352
rect 176285 36410 176351 36413
rect 216397 36410 216463 36413
rect 176285 36408 176394 36410
rect 176285 36352 176290 36408
rect 176346 36352 176394 36408
rect 176285 36347 176394 36352
rect 216397 36408 216506 36410
rect 216397 36352 216402 36408
rect 216458 36352 216506 36408
rect 216397 36347 216506 36352
rect 96294 36244 96354 36347
rect 136909 36274 136975 36277
rect 136436 36272 136975 36274
rect 136436 36216 136914 36272
rect 136970 36216 136975 36272
rect 176334 36244 176394 36347
rect 216446 36244 216506 36347
rect 257613 36274 257679 36277
rect 257140 36272 257679 36274
rect 136436 36214 136975 36216
rect 257140 36216 257618 36272
rect 257674 36216 257679 36272
rect 257140 36214 257679 36216
rect 136909 36211 136975 36214
rect 257613 36211 257679 36214
rect 68369 35730 68435 35733
rect 65964 35728 68435 35730
rect 65964 35672 68374 35728
rect 68430 35672 68435 35728
rect 65964 35670 68435 35672
rect 68369 35667 68435 35670
rect 88149 35458 88215 35461
rect 128169 35458 128235 35461
rect 169569 35458 169635 35461
rect 209497 35458 209563 35461
rect 88149 35456 90436 35458
rect 88149 35400 88154 35456
rect 88210 35400 90436 35456
rect 88149 35398 90436 35400
rect 128169 35456 130732 35458
rect 128169 35400 128174 35456
rect 128230 35400 130732 35456
rect 128169 35398 130732 35400
rect 169569 35456 170844 35458
rect 169569 35400 169574 35456
rect 169630 35400 170844 35456
rect 169569 35398 170844 35400
rect 209497 35456 211140 35458
rect 209497 35400 209502 35456
rect 209558 35400 211140 35456
rect 209497 35398 211140 35400
rect 88149 35395 88215 35398
rect 128169 35395 128235 35398
rect 169569 35395 169635 35398
rect 209497 35395 209563 35398
rect 17861 35050 17927 35053
rect 96889 35050 96955 35053
rect 136265 35050 136331 35053
rect 177849 35050 177915 35053
rect 17861 35048 20148 35050
rect 17861 34992 17866 35048
rect 17922 34992 20148 35048
rect 17861 34990 20148 34992
rect 96889 35048 97704 35050
rect 96889 34992 96894 35048
rect 96950 34992 97704 35048
rect 96889 34990 97704 34992
rect 136265 35048 137908 35050
rect 136265 34992 136270 35048
rect 136326 34992 137908 35048
rect 136265 34990 137908 34992
rect 177849 35048 178112 35050
rect 177849 34992 177854 35048
rect 177910 34992 178112 35048
rect 177849 34990 178112 34992
rect 17861 34987 17927 34990
rect 96889 34987 96955 34990
rect 136265 34987 136331 34990
rect 177849 34987 177915 34990
rect 217961 34982 218027 34985
rect 258257 34982 258323 34985
rect 217961 34980 218316 34982
rect 217961 34924 217966 34980
rect 218022 34924 218316 34980
rect 217961 34922 218316 34924
rect 258257 34980 258520 34982
rect 258257 34924 258262 34980
rect 258318 34924 258520 34980
rect 258257 34922 258520 34924
rect 217961 34919 218027 34922
rect 258257 34919 258323 34922
rect 136357 34914 136423 34917
rect 176377 34914 176443 34917
rect 136357 34912 136466 34914
rect 136357 34856 136362 34912
rect 136418 34856 136466 34912
rect 136357 34851 136466 34856
rect 96797 34778 96863 34781
rect 96324 34776 96863 34778
rect 96324 34720 96802 34776
rect 96858 34720 96863 34776
rect 136406 34748 136466 34851
rect 176334 34912 176443 34914
rect 176334 34856 176382 34912
rect 176438 34856 176443 34912
rect 176334 34851 176443 34856
rect 176334 34748 176394 34851
rect 217501 34778 217567 34781
rect 257889 34778 257955 34781
rect 216844 34776 217567 34778
rect 96324 34718 96863 34720
rect 216844 34720 217506 34776
rect 217562 34720 217567 34776
rect 216844 34718 217567 34720
rect 257140 34776 257955 34778
rect 257140 34720 257894 34776
rect 257950 34720 257955 34776
rect 257140 34718 257955 34720
rect 96797 34715 96863 34718
rect 217501 34715 217567 34718
rect 257889 34715 257955 34718
rect 68369 34370 68435 34373
rect 65964 34368 68435 34370
rect 65964 34312 68374 34368
rect 68430 34312 68435 34368
rect 65964 34310 68435 34312
rect 68369 34307 68435 34310
rect 17769 33690 17835 33693
rect 17769 33688 20148 33690
rect 17769 33632 17774 33688
rect 17830 33632 20148 33688
rect 17769 33630 20148 33632
rect 17769 33627 17835 33630
rect 136449 33418 136515 33421
rect 136406 33416 136515 33418
rect 136406 33360 136454 33416
rect 136510 33360 136515 33416
rect 136406 33355 136515 33360
rect 176469 33418 176535 33421
rect 176469 33416 176578 33418
rect 176469 33360 176474 33416
rect 176530 33360 176578 33416
rect 176469 33355 176578 33360
rect 96613 33282 96679 33285
rect 96324 33280 96679 33282
rect 96324 33224 96618 33280
rect 96674 33224 96679 33280
rect 136406 33252 136466 33355
rect 176518 33252 176578 33355
rect 217409 33282 217475 33285
rect 257981 33282 258047 33285
rect 216844 33280 217475 33282
rect 96324 33222 96679 33224
rect 216844 33224 217414 33280
rect 217470 33224 217475 33280
rect 216844 33222 217475 33224
rect 257140 33280 258047 33282
rect 257140 33224 257986 33280
rect 258042 33224 258047 33280
rect 257140 33222 258047 33224
rect 96613 33219 96679 33222
rect 217409 33219 217475 33222
rect 257981 33219 258047 33222
rect 580165 33146 580231 33149
rect 583520 33146 584960 33236
rect 580165 33144 584960 33146
rect 580165 33088 580170 33144
rect 580226 33088 584960 33144
rect 580165 33086 584960 33088
rect 580165 33083 580231 33086
rect 583520 32996 584960 33086
rect 97533 32738 97599 32741
rect 97674 32738 97734 32980
rect 97533 32736 97734 32738
rect 97533 32680 97538 32736
rect 97594 32680 97734 32736
rect 97533 32678 97734 32680
rect 97533 32675 97599 32678
rect -960 32316 480 32556
rect 88057 32466 88123 32469
rect 127985 32466 128051 32469
rect 88057 32464 90436 32466
rect 88057 32408 88062 32464
rect 88118 32408 90436 32464
rect 88057 32406 90436 32408
rect 127985 32464 130732 32466
rect 127985 32408 127990 32464
rect 128046 32408 130732 32464
rect 127985 32406 130732 32408
rect 88057 32403 88123 32406
rect 127985 32403 128051 32406
rect 68461 32330 68527 32333
rect 65964 32328 68527 32330
rect 65964 32272 68466 32328
rect 68522 32272 68527 32328
rect 65964 32270 68527 32272
rect 68461 32267 68527 32270
rect 136633 32330 136699 32333
rect 137878 32330 137938 32912
rect 178082 32741 178142 32980
rect 217961 32942 218027 32945
rect 217961 32940 218316 32942
rect 217961 32884 217966 32940
rect 218022 32884 218316 32940
rect 217961 32882 218316 32884
rect 258030 32882 258520 32942
rect 217961 32879 218027 32882
rect 258030 32877 258090 32882
rect 257981 32872 258090 32877
rect 257981 32816 257986 32872
rect 258042 32816 258090 32872
rect 257981 32814 258090 32816
rect 257981 32811 258047 32814
rect 178033 32736 178142 32741
rect 178033 32680 178038 32736
rect 178094 32680 178142 32736
rect 178033 32678 178142 32680
rect 178033 32675 178099 32678
rect 169477 32466 169543 32469
rect 209405 32466 209471 32469
rect 169477 32464 170844 32466
rect 169477 32408 169482 32464
rect 169538 32408 170844 32464
rect 169477 32406 170844 32408
rect 209405 32464 211140 32466
rect 209405 32408 209410 32464
rect 209466 32408 211140 32464
rect 209405 32406 211140 32408
rect 169477 32403 169543 32406
rect 209405 32403 209471 32406
rect 136633 32328 137938 32330
rect 136633 32272 136638 32328
rect 136694 32272 137938 32328
rect 136633 32270 137938 32272
rect 136633 32267 136699 32270
rect 96337 31922 96403 31925
rect 136541 31922 136607 31925
rect 176561 31922 176627 31925
rect 96294 31920 96403 31922
rect 96294 31864 96342 31920
rect 96398 31864 96403 31920
rect 96294 31859 96403 31864
rect 136406 31920 136607 31922
rect 136406 31864 136546 31920
rect 136602 31864 136607 31920
rect 136406 31862 136607 31864
rect 96294 31756 96354 31859
rect 136406 31756 136466 31862
rect 136541 31859 136607 31862
rect 176518 31920 176627 31922
rect 176518 31864 176566 31920
rect 176622 31864 176627 31920
rect 176518 31859 176627 31864
rect 216581 31922 216647 31925
rect 216581 31920 216690 31922
rect 216581 31864 216586 31920
rect 216642 31864 216690 31920
rect 216581 31859 216690 31864
rect 176518 31756 176578 31859
rect 216630 31756 216690 31859
rect 257337 31786 257403 31789
rect 257140 31784 257403 31786
rect 257140 31728 257342 31784
rect 257398 31728 257403 31784
rect 257140 31726 257403 31728
rect 257337 31723 257403 31726
rect 17585 31650 17651 31653
rect 17585 31648 20148 31650
rect 17585 31592 17590 31648
rect 17646 31592 20148 31648
rect 17585 31590 20148 31592
rect 17585 31587 17651 31590
rect 67725 30970 67791 30973
rect 65964 30968 67791 30970
rect 65964 30912 67730 30968
rect 67786 30912 67791 30968
rect 65964 30910 67791 30912
rect 67725 30907 67791 30910
rect 97349 30970 97415 30973
rect 97349 30968 97704 30970
rect 97349 30912 97354 30968
rect 97410 30912 97704 30968
rect 97349 30910 97704 30912
rect 97349 30907 97415 30910
rect 218053 30902 218119 30905
rect 218053 30900 218316 30902
rect 136265 30426 136331 30429
rect 136222 30424 136331 30426
rect 136222 30368 136270 30424
rect 136326 30368 136331 30424
rect 136222 30363 136331 30368
rect 136725 30426 136791 30429
rect 137878 30426 137938 30872
rect 178174 30701 178234 30872
rect 218053 30844 218058 30900
rect 218114 30844 218316 30900
rect 218053 30842 218316 30844
rect 258030 30842 258520 30902
rect 218053 30839 218119 30842
rect 257429 30834 257495 30837
rect 258030 30834 258090 30842
rect 257429 30832 258090 30834
rect 257429 30776 257434 30832
rect 257490 30776 258090 30832
rect 257429 30774 258090 30776
rect 257429 30771 257495 30774
rect 178125 30696 178234 30701
rect 178125 30640 178130 30696
rect 178186 30640 178234 30696
rect 178125 30638 178234 30640
rect 178125 30635 178191 30638
rect 176745 30426 176811 30429
rect 216857 30426 216923 30429
rect 257153 30426 257219 30429
rect 136725 30424 137938 30426
rect 136725 30368 136730 30424
rect 136786 30368 137938 30424
rect 136725 30366 137938 30368
rect 176702 30424 176811 30426
rect 176702 30368 176750 30424
rect 176806 30368 176811 30424
rect 136725 30363 136791 30366
rect 176702 30363 176811 30368
rect 216814 30424 216923 30426
rect 216814 30368 216862 30424
rect 216918 30368 216923 30424
rect 216814 30363 216923 30368
rect 257110 30424 257219 30426
rect 257110 30368 257158 30424
rect 257214 30368 257219 30424
rect 257110 30363 257219 30368
rect 17769 30290 17835 30293
rect 96889 30290 96955 30293
rect 17769 30288 20148 30290
rect 17769 30232 17774 30288
rect 17830 30232 20148 30288
rect 17769 30230 20148 30232
rect 96324 30288 96955 30290
rect 96324 30232 96894 30288
rect 96950 30232 96955 30288
rect 136222 30260 136282 30363
rect 176702 30260 176762 30363
rect 216814 30260 216874 30363
rect 257110 30260 257170 30363
rect 96324 30230 96955 30232
rect 17769 30227 17835 30230
rect 96889 30227 96955 30230
rect 87597 29474 87663 29477
rect 127617 29474 127683 29477
rect 169017 29474 169083 29477
rect 209037 29474 209103 29477
rect 249057 29474 249123 29477
rect 87597 29472 90436 29474
rect 87597 29416 87602 29472
rect 87658 29416 90436 29472
rect 87597 29414 90436 29416
rect 127617 29472 130732 29474
rect 127617 29416 127622 29472
rect 127678 29416 130732 29472
rect 127617 29414 130732 29416
rect 169017 29472 170844 29474
rect 169017 29416 169022 29472
rect 169078 29416 170844 29472
rect 169017 29414 170844 29416
rect 209037 29472 211140 29474
rect 209037 29416 209042 29472
rect 209098 29416 211140 29472
rect 209037 29414 211140 29416
rect 249057 29472 251252 29474
rect 249057 29416 249062 29472
rect 249118 29416 251252 29472
rect 249057 29414 251252 29416
rect 87597 29411 87663 29414
rect 127617 29411 127683 29414
rect 169017 29411 169083 29414
rect 209037 29411 209103 29414
rect 249057 29411 249123 29414
rect 68461 28930 68527 28933
rect 96337 28930 96403 28933
rect 65964 28928 68527 28930
rect 65964 28872 68466 28928
rect 68522 28872 68527 28928
rect 65964 28870 68527 28872
rect 68461 28867 68527 28870
rect 96294 28928 96403 28930
rect 96294 28872 96342 28928
rect 96398 28872 96403 28928
rect 96294 28867 96403 28872
rect 97441 28930 97507 28933
rect 136633 28930 136699 28933
rect 176561 28930 176627 28933
rect 97441 28928 97704 28930
rect 97441 28872 97446 28928
rect 97502 28872 97704 28928
rect 97441 28870 97704 28872
rect 136406 28928 136699 28930
rect 136406 28872 136638 28928
rect 136694 28872 136699 28928
rect 136406 28870 136699 28872
rect 97441 28867 97507 28870
rect 96294 28764 96354 28867
rect 136406 28764 136466 28870
rect 136633 28867 136699 28870
rect 176518 28928 176627 28930
rect 176518 28872 176566 28928
rect 176622 28872 176627 28928
rect 176518 28867 176627 28872
rect 177849 28930 177915 28933
rect 216489 28930 216555 28933
rect 177849 28928 178112 28930
rect 177849 28872 177854 28928
rect 177910 28872 178112 28928
rect 177849 28870 178112 28872
rect 216446 28928 216555 28930
rect 216446 28872 216494 28928
rect 216550 28872 216555 28928
rect 177849 28867 177915 28870
rect 216446 28867 216555 28872
rect 17677 28250 17743 28253
rect 136449 28250 136515 28253
rect 137878 28250 137938 28832
rect 176518 28764 176578 28867
rect 216446 28764 216506 28867
rect 217961 28862 218027 28865
rect 258257 28862 258323 28865
rect 217961 28860 218316 28862
rect 217961 28804 217966 28860
rect 218022 28804 218316 28860
rect 217961 28802 218316 28804
rect 258257 28860 258520 28862
rect 258257 28804 258262 28860
rect 258318 28804 258520 28860
rect 258257 28802 258520 28804
rect 217961 28799 218027 28802
rect 258257 28799 258323 28802
rect 257981 28794 258047 28797
rect 257140 28792 258047 28794
rect 257140 28736 257986 28792
rect 258042 28736 258047 28792
rect 257140 28734 258047 28736
rect 257981 28731 258047 28734
rect 17677 28248 20148 28250
rect 17677 28192 17682 28248
rect 17738 28192 20148 28248
rect 17677 28190 20148 28192
rect 136449 28248 137938 28250
rect 136449 28192 136454 28248
rect 136510 28192 137938 28248
rect 136449 28190 137938 28192
rect 17677 28187 17743 28190
rect 136449 28187 136515 28190
rect 68277 27570 68343 27573
rect 65964 27568 68343 27570
rect 65964 27512 68282 27568
rect 68338 27512 68343 27568
rect 65964 27510 68343 27512
rect 68277 27507 68343 27510
rect 96337 27434 96403 27437
rect 176561 27434 176627 27437
rect 96294 27432 96403 27434
rect 96294 27376 96342 27432
rect 96398 27376 96403 27432
rect 96294 27371 96403 27376
rect 176518 27432 176627 27434
rect 176518 27376 176566 27432
rect 176622 27376 176627 27432
rect 176518 27371 176627 27376
rect 216581 27434 216647 27437
rect 216581 27432 216690 27434
rect 216581 27376 216586 27432
rect 216642 27376 216690 27432
rect 216581 27371 216690 27376
rect 96294 27268 96354 27371
rect 136725 27298 136791 27301
rect 136436 27296 136791 27298
rect 136436 27240 136730 27296
rect 136786 27240 136791 27296
rect 176518 27268 176578 27371
rect 216630 27268 216690 27371
rect 257429 27298 257495 27301
rect 257140 27296 257495 27298
rect 136436 27238 136791 27240
rect 257140 27240 257434 27296
rect 257490 27240 257495 27296
rect 257140 27238 257495 27240
rect 136725 27235 136791 27238
rect 257429 27235 257495 27238
rect 17861 26890 17927 26893
rect 97441 26890 97507 26893
rect 177849 26890 177915 26893
rect 17861 26888 20148 26890
rect 17861 26832 17866 26888
rect 17922 26832 20148 26888
rect 17861 26830 20148 26832
rect 97441 26888 97704 26890
rect 97441 26832 97446 26888
rect 97502 26832 97704 26888
rect 97441 26830 97704 26832
rect 177849 26888 178112 26890
rect 177849 26832 177854 26888
rect 177910 26832 178112 26888
rect 177849 26830 178112 26832
rect 17861 26827 17927 26830
rect 97441 26827 97507 26830
rect 177849 26827 177915 26830
rect 218053 26822 218119 26825
rect 258257 26822 258323 26825
rect 218053 26820 218316 26822
rect 136265 26618 136331 26621
rect 137878 26618 137938 26792
rect 218053 26764 218058 26820
rect 218114 26764 218316 26820
rect 218053 26762 218316 26764
rect 258257 26820 258520 26822
rect 258257 26764 258262 26820
rect 258318 26764 258520 26820
rect 258257 26762 258520 26764
rect 218053 26759 218119 26762
rect 258257 26759 258323 26762
rect 136265 26616 137938 26618
rect 136265 26560 136270 26616
rect 136326 26560 137938 26616
rect 136265 26558 137938 26560
rect 136265 26555 136331 26558
rect 87413 26482 87479 26485
rect 127525 26482 127591 26485
rect 169109 26482 169175 26485
rect 208485 26482 208551 26485
rect 249149 26482 249215 26485
rect 87413 26480 90436 26482
rect 87413 26424 87418 26480
rect 87474 26424 90436 26480
rect 87413 26422 90436 26424
rect 127525 26480 130732 26482
rect 127525 26424 127530 26480
rect 127586 26424 130732 26480
rect 127525 26422 130732 26424
rect 169109 26480 170844 26482
rect 169109 26424 169114 26480
rect 169170 26424 170844 26480
rect 169109 26422 170844 26424
rect 208485 26480 211140 26482
rect 208485 26424 208490 26480
rect 208546 26424 211140 26480
rect 208485 26422 211140 26424
rect 249149 26480 251252 26482
rect 249149 26424 249154 26480
rect 249210 26424 251252 26480
rect 249149 26422 251252 26424
rect 87413 26419 87479 26422
rect 127525 26419 127591 26422
rect 169109 26419 169175 26422
rect 208485 26419 208551 26422
rect 249149 26419 249215 26422
rect 136449 25938 136515 25941
rect 176745 25938 176811 25941
rect 216857 25938 216923 25941
rect 136406 25936 136515 25938
rect 136406 25880 136454 25936
rect 136510 25880 136515 25936
rect 136406 25875 136515 25880
rect 176702 25936 176811 25938
rect 176702 25880 176750 25936
rect 176806 25880 176811 25936
rect 176702 25875 176811 25880
rect 216814 25936 216923 25938
rect 216814 25880 216862 25936
rect 216918 25880 216923 25936
rect 216814 25875 216923 25880
rect 96521 25802 96587 25805
rect 96324 25800 96587 25802
rect 96324 25744 96526 25800
rect 96582 25744 96587 25800
rect 136406 25772 136466 25875
rect 176702 25772 176762 25875
rect 216814 25772 216874 25875
rect 257337 25802 257403 25805
rect 257140 25800 257403 25802
rect 96324 25742 96587 25744
rect 257140 25744 257342 25800
rect 257398 25744 257403 25800
rect 257140 25742 257403 25744
rect 96521 25739 96587 25742
rect 257337 25739 257403 25742
rect 67633 25530 67699 25533
rect 65964 25528 67699 25530
rect 65964 25472 67638 25528
rect 67694 25472 67699 25528
rect 65964 25470 67699 25472
rect 67633 25467 67699 25470
rect 17861 24850 17927 24853
rect 97441 24850 97507 24853
rect 17861 24848 20148 24850
rect 17861 24792 17866 24848
rect 17922 24792 20148 24848
rect 17861 24790 20148 24792
rect 97441 24848 97704 24850
rect 97441 24792 97446 24848
rect 97502 24792 97704 24848
rect 97441 24790 97704 24792
rect 17861 24787 17927 24790
rect 97441 24787 97507 24790
rect 218053 24782 218119 24785
rect 258257 24782 258323 24785
rect 218053 24780 218316 24782
rect 65333 24714 65399 24717
rect 65333 24712 65442 24714
rect 65333 24656 65338 24712
rect 65394 24656 65442 24712
rect 65333 24651 65442 24656
rect 15837 24170 15903 24173
rect 15837 24168 20178 24170
rect 15837 24112 15842 24168
rect 15898 24112 20178 24168
rect 65382 24140 65442 24651
rect 96337 24442 96403 24445
rect 136265 24442 136331 24445
rect 96294 24440 96403 24442
rect 96294 24384 96342 24440
rect 96398 24384 96403 24440
rect 96294 24379 96403 24384
rect 136222 24440 136331 24442
rect 136222 24384 136270 24440
rect 136326 24384 136331 24440
rect 136222 24379 136331 24384
rect 136449 24442 136515 24445
rect 137878 24442 137938 24752
rect 178174 24581 178234 24752
rect 218053 24724 218058 24780
rect 218114 24724 218316 24780
rect 218053 24722 218316 24724
rect 258257 24780 258520 24782
rect 258257 24724 258262 24780
rect 258318 24724 258520 24780
rect 258257 24722 258520 24724
rect 218053 24719 218119 24722
rect 258257 24719 258323 24722
rect 178125 24576 178234 24581
rect 178125 24520 178130 24576
rect 178186 24520 178234 24576
rect 178125 24518 178234 24520
rect 178125 24515 178191 24518
rect 176745 24442 176811 24445
rect 136449 24440 137938 24442
rect 136449 24384 136454 24440
rect 136510 24384 137938 24440
rect 136449 24382 137938 24384
rect 176702 24440 176811 24442
rect 176702 24384 176750 24440
rect 176806 24384 176811 24440
rect 136449 24379 136515 24382
rect 176702 24379 176811 24384
rect 216765 24442 216831 24445
rect 257153 24442 257219 24445
rect 216765 24440 216874 24442
rect 216765 24384 216770 24440
rect 216826 24384 216874 24440
rect 216765 24379 216874 24384
rect 96294 24276 96354 24379
rect 136222 24276 136282 24379
rect 176702 24276 176762 24379
rect 216814 24276 216874 24379
rect 257110 24440 257219 24442
rect 257110 24384 257158 24440
rect 257214 24384 257219 24440
rect 257110 24379 257219 24384
rect 257110 24276 257170 24379
rect 15837 24110 20178 24112
rect 15837 24107 15903 24110
rect 20118 23460 20178 24110
rect 87229 23490 87295 23493
rect 127065 23490 127131 23493
rect 168373 23490 168439 23493
rect 208577 23490 208643 23493
rect 248597 23490 248663 23493
rect 87229 23488 90436 23490
rect 87229 23432 87234 23488
rect 87290 23432 90436 23488
rect 87229 23430 90436 23432
rect 127065 23488 130732 23490
rect 127065 23432 127070 23488
rect 127126 23432 130732 23488
rect 127065 23430 130732 23432
rect 168373 23488 170844 23490
rect 168373 23432 168378 23488
rect 168434 23432 170844 23488
rect 168373 23430 170844 23432
rect 208577 23488 211140 23490
rect 208577 23432 208582 23488
rect 208638 23432 211140 23488
rect 208577 23430 211140 23432
rect 248597 23488 251252 23490
rect 248597 23432 248602 23488
rect 248658 23432 251252 23488
rect 248597 23430 251252 23432
rect 87229 23427 87295 23430
rect 127065 23427 127131 23430
rect 168373 23427 168439 23430
rect 208577 23427 208643 23430
rect 248597 23427 248663 23430
rect 96337 22946 96403 22949
rect 136449 22946 136515 22949
rect 176561 22946 176627 22949
rect 96294 22944 96403 22946
rect 96294 22888 96342 22944
rect 96398 22888 96403 22944
rect 96294 22883 96403 22888
rect 136406 22944 136515 22946
rect 136406 22888 136454 22944
rect 136510 22888 136515 22944
rect 136406 22883 136515 22888
rect 176518 22944 176627 22946
rect 176518 22888 176566 22944
rect 176622 22888 176627 22944
rect 176518 22883 176627 22888
rect 216581 22946 216647 22949
rect 257153 22946 257219 22949
rect 216581 22944 216690 22946
rect 216581 22888 216586 22944
rect 216642 22888 216690 22944
rect 216581 22883 216690 22888
rect 96294 22780 96354 22883
rect 97441 22810 97507 22813
rect 97441 22808 97704 22810
rect 97441 22752 97446 22808
rect 97502 22752 97704 22808
rect 136406 22780 136466 22883
rect 176518 22780 176578 22883
rect 216630 22780 216690 22883
rect 257110 22944 257219 22946
rect 257110 22888 257158 22944
rect 257214 22888 257219 22944
rect 257110 22883 257219 22888
rect 257110 22780 257170 22883
rect 97441 22750 97704 22752
rect 97441 22747 97507 22750
rect 218053 22742 218119 22745
rect 258257 22742 258323 22745
rect 218053 22740 218316 22742
rect 68553 22130 68619 22133
rect 137878 22130 137938 22712
rect 178174 22541 178234 22712
rect 218053 22684 218058 22740
rect 218114 22684 218316 22740
rect 218053 22682 218316 22684
rect 258257 22740 258520 22742
rect 258257 22684 258262 22740
rect 258318 22684 258520 22740
rect 258257 22682 258520 22684
rect 218053 22679 218119 22682
rect 258257 22679 258323 22682
rect 178125 22536 178234 22541
rect 178125 22480 178130 22536
rect 178186 22480 178234 22536
rect 178125 22478 178234 22480
rect 178125 22475 178191 22478
rect 65964 22128 68619 22130
rect 65964 22072 68558 22128
rect 68614 22072 68619 22128
rect 65964 22070 68619 22072
rect 68553 22067 68619 22070
rect 136406 22070 137938 22130
rect 17769 21450 17835 21453
rect 96337 21450 96403 21453
rect 17769 21448 20148 21450
rect 17769 21392 17774 21448
rect 17830 21392 20148 21448
rect 17769 21390 20148 21392
rect 96294 21448 96403 21450
rect 96294 21392 96342 21448
rect 96398 21392 96403 21448
rect 17769 21387 17835 21390
rect 96294 21387 96403 21392
rect 96294 21284 96354 21387
rect 136406 21284 136466 22070
rect 176561 21450 176627 21453
rect 176518 21448 176627 21450
rect 176518 21392 176566 21448
rect 176622 21392 176627 21448
rect 176518 21387 176627 21392
rect 216581 21450 216647 21453
rect 257153 21450 257219 21453
rect 216581 21448 216690 21450
rect 216581 21392 216586 21448
rect 216642 21392 216690 21448
rect 216581 21387 216690 21392
rect 176518 21284 176578 21387
rect 216630 21284 216690 21387
rect 257110 21448 257219 21450
rect 257110 21392 257158 21448
rect 257214 21392 257219 21448
rect 257110 21387 257219 21392
rect 257110 21284 257170 21387
rect 218053 20770 218119 20773
rect 21633 20634 21699 20637
rect 21950 20634 21956 20636
rect 21633 20632 21956 20634
rect 21633 20576 21638 20632
rect 21694 20576 21956 20632
rect 21633 20574 21956 20576
rect 21633 20571 21699 20574
rect 21950 20572 21956 20574
rect 22020 20572 22026 20636
rect 65934 20634 65994 20740
rect 66161 20634 66227 20637
rect 65934 20632 66227 20634
rect 65934 20576 66166 20632
rect 66222 20576 66227 20632
rect 65934 20574 66227 20576
rect 66161 20571 66227 20574
rect 60590 20436 60596 20500
rect 60660 20498 60666 20500
rect 60660 20438 90436 20498
rect 60660 20436 60666 20438
rect 97674 20362 97734 20740
rect 136406 20710 137908 20770
rect 218053 20768 218316 20770
rect 126973 20498 127039 20501
rect 126973 20496 130732 20498
rect 126973 20440 126978 20496
rect 127034 20440 130732 20496
rect 126973 20438 130732 20440
rect 126973 20435 127039 20438
rect 96294 20302 97734 20362
rect 96294 19788 96354 20302
rect 136406 19788 136466 20710
rect 136541 19954 136607 19957
rect 170814 19954 170874 20468
rect 178082 20362 178142 20740
rect 218053 20712 218058 20768
rect 218114 20712 218316 20768
rect 218053 20710 218316 20712
rect 218053 20707 218119 20710
rect 258030 20642 258520 20702
rect 208393 20498 208459 20501
rect 249701 20498 249767 20501
rect 258030 20498 258090 20642
rect 208393 20496 211140 20498
rect 208393 20440 208398 20496
rect 208454 20440 211140 20496
rect 208393 20438 211140 20440
rect 249701 20496 251252 20498
rect 249701 20440 249706 20496
rect 249762 20440 251252 20496
rect 249701 20438 251252 20440
rect 257110 20438 258090 20498
rect 208393 20435 208459 20438
rect 249701 20435 249767 20438
rect 136541 19952 170874 19954
rect 136541 19896 136546 19952
rect 136602 19896 170874 19952
rect 136541 19894 170874 19896
rect 176518 20302 178142 20362
rect 136541 19891 136607 19894
rect 176518 19788 176578 20302
rect 216581 20226 216647 20229
rect 216581 20224 216690 20226
rect 216581 20168 216586 20224
rect 216642 20168 216690 20224
rect 216581 20163 216690 20168
rect 216630 19788 216690 20163
rect 257110 19788 257170 20438
rect 583520 19668 584960 19908
rect 88241 19546 88307 19549
rect 127065 19546 127131 19549
rect 88241 19544 127131 19546
rect -960 19410 480 19500
rect 88241 19488 88246 19544
rect 88302 19488 127070 19544
rect 127126 19488 127131 19544
rect 88241 19486 127131 19488
rect 88241 19483 88307 19486
rect 127065 19483 127131 19486
rect 169661 19546 169727 19549
rect 208577 19546 208643 19549
rect 169661 19544 208643 19546
rect 169661 19488 169666 19544
rect 169722 19488 208582 19544
rect 208638 19488 208643 19544
rect 169661 19486 208643 19488
rect 169661 19483 169727 19486
rect 208577 19483 208643 19486
rect 3233 19410 3299 19413
rect -960 19408 3299 19410
rect -960 19352 3238 19408
rect 3294 19352 3299 19408
rect -960 19350 3299 19352
rect -960 19260 480 19350
rect 3233 19347 3299 19350
rect 3734 17716 3740 17780
rect 3804 17778 3810 17780
rect 50245 17778 50311 17781
rect 3804 17776 50311 17778
rect 3804 17720 50250 17776
rect 50306 17720 50311 17776
rect 3804 17718 50311 17720
rect 3804 17716 3810 17718
rect 50245 17715 50311 17718
rect 3366 17580 3372 17644
rect 3436 17642 3442 17644
rect 39297 17642 39363 17645
rect 3436 17640 39363 17642
rect 3436 17584 39302 17640
rect 39358 17584 39363 17640
rect 3436 17582 39363 17584
rect 3436 17580 3442 17582
rect 39297 17579 39363 17582
rect 3550 17444 3556 17508
rect 3620 17506 3626 17508
rect 32857 17506 32923 17509
rect 3620 17504 32923 17506
rect 3620 17448 32862 17504
rect 32918 17448 32923 17504
rect 3620 17446 32923 17448
rect 3620 17444 3626 17446
rect 32857 17443 32923 17446
rect 3918 17308 3924 17372
rect 3988 17370 3994 17372
rect 61837 17370 61903 17373
rect 3988 17368 61903 17370
rect 3988 17312 61842 17368
rect 61898 17312 61903 17368
rect 3988 17310 61903 17312
rect 3988 17308 3994 17310
rect 61837 17307 61903 17310
rect -960 6490 480 6580
rect 46974 6490 46980 6492
rect -960 6430 46980 6490
rect -960 6340 480 6430
rect 46974 6428 46980 6430
rect 47044 6428 47050 6492
rect 583520 6476 584960 6716
rect 55070 3436 55076 3500
rect 55140 3498 55146 3500
rect 132953 3498 133019 3501
rect 55140 3496 133019 3498
rect 55140 3440 132958 3496
rect 133014 3440 133019 3496
rect 55140 3438 133019 3440
rect 55140 3436 55146 3438
rect 132953 3435 133019 3438
rect 44030 3300 44036 3364
rect 44100 3362 44106 3364
rect 136449 3362 136515 3365
rect 44100 3360 136515 3362
rect 44100 3304 136454 3360
rect 136510 3304 136515 3360
rect 44100 3302 136515 3304
rect 44100 3300 44106 3302
rect 136449 3299 136515 3302
<< via3 >>
rect 3372 606052 3436 606116
rect 3556 579940 3620 580004
rect 3740 501740 3804 501804
rect 3924 475628 3988 475692
rect 21956 325212 22020 325276
rect 44036 39400 44100 39404
rect 44036 39344 44050 39400
rect 44050 39344 44100 39400
rect 44036 39340 44100 39344
rect 46980 39340 47044 39404
rect 55076 39340 55140 39404
rect 60596 39264 60660 39268
rect 60596 39208 60610 39264
rect 60610 39208 60660 39264
rect 60596 39204 60660 39208
rect 21956 20572 22020 20636
rect 60596 20436 60660 20500
rect 3740 17716 3804 17780
rect 3372 17580 3436 17644
rect 3556 17444 3620 17508
rect 3924 17308 3988 17372
rect 46980 6428 47044 6492
rect 55076 3436 55140 3500
rect 44036 3300 44100 3364
<< metal4 >>
rect -8726 711558 -8106 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 -8106 711558
rect -8726 711238 -8106 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 -8106 711238
rect -8726 -7066 -8106 711002
rect -7766 710598 -7146 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 -7146 710598
rect -7766 710278 -7146 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 -7146 710278
rect -7766 -6106 -7146 710042
rect -6806 709638 -6186 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 -6186 709638
rect -6806 709318 -6186 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 -6186 709318
rect -6806 -5146 -6186 709082
rect -5846 708678 -5226 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 -5226 708678
rect -5846 708358 -5226 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 -5226 708358
rect -5846 -4186 -5226 708122
rect -4886 707718 -4266 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 -4266 707718
rect -4886 707398 -4266 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 -4266 707398
rect -4886 -3226 -4266 707162
rect -3926 706758 -3306 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 -3306 706758
rect -3926 706438 -3306 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 -3306 706438
rect -3926 -2266 -3306 706202
rect -2966 705798 -2346 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 -2346 705798
rect -2966 705478 -2346 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 -2346 705478
rect -2966 694454 -2346 705242
rect 37994 705798 38614 711590
rect 37994 705562 38026 705798
rect 38262 705562 38346 705798
rect 38582 705562 38614 705798
rect 37994 705478 38614 705562
rect 37994 705242 38026 705478
rect 38262 705242 38346 705478
rect 38582 705242 38614 705478
rect -2966 694218 -2934 694454
rect -2698 694218 -2614 694454
rect -2378 694218 -2346 694454
rect -2966 694134 -2346 694218
rect -2966 693898 -2934 694134
rect -2698 693898 -2614 694134
rect -2378 693898 -2346 694134
rect -2966 657454 -2346 693898
rect -2966 657218 -2934 657454
rect -2698 657218 -2614 657454
rect -2378 657218 -2346 657454
rect -2966 657134 -2346 657218
rect -2966 656898 -2934 657134
rect -2698 656898 -2614 657134
rect -2378 656898 -2346 657134
rect -2966 620454 -2346 656898
rect -2966 620218 -2934 620454
rect -2698 620218 -2614 620454
rect -2378 620218 -2346 620454
rect -2966 620134 -2346 620218
rect -2966 619898 -2934 620134
rect -2698 619898 -2614 620134
rect -2378 619898 -2346 620134
rect -2966 583454 -2346 619898
rect -2966 583218 -2934 583454
rect -2698 583218 -2614 583454
rect -2378 583218 -2346 583454
rect -2966 583134 -2346 583218
rect -2966 582898 -2934 583134
rect -2698 582898 -2614 583134
rect -2378 582898 -2346 583134
rect -2966 546454 -2346 582898
rect -2966 546218 -2934 546454
rect -2698 546218 -2614 546454
rect -2378 546218 -2346 546454
rect -2966 546134 -2346 546218
rect -2966 545898 -2934 546134
rect -2698 545898 -2614 546134
rect -2378 545898 -2346 546134
rect -2966 509454 -2346 545898
rect -2966 509218 -2934 509454
rect -2698 509218 -2614 509454
rect -2378 509218 -2346 509454
rect -2966 509134 -2346 509218
rect -2966 508898 -2934 509134
rect -2698 508898 -2614 509134
rect -2378 508898 -2346 509134
rect -2966 472454 -2346 508898
rect -2966 472218 -2934 472454
rect -2698 472218 -2614 472454
rect -2378 472218 -2346 472454
rect -2966 472134 -2346 472218
rect -2966 471898 -2934 472134
rect -2698 471898 -2614 472134
rect -2378 471898 -2346 472134
rect -2966 435454 -2346 471898
rect -2966 435218 -2934 435454
rect -2698 435218 -2614 435454
rect -2378 435218 -2346 435454
rect -2966 435134 -2346 435218
rect -2966 434898 -2934 435134
rect -2698 434898 -2614 435134
rect -2378 434898 -2346 435134
rect -2966 398454 -2346 434898
rect -2966 398218 -2934 398454
rect -2698 398218 -2614 398454
rect -2378 398218 -2346 398454
rect -2966 398134 -2346 398218
rect -2966 397898 -2934 398134
rect -2698 397898 -2614 398134
rect -2378 397898 -2346 398134
rect -2966 361454 -2346 397898
rect -2966 361218 -2934 361454
rect -2698 361218 -2614 361454
rect -2378 361218 -2346 361454
rect -2966 361134 -2346 361218
rect -2966 360898 -2934 361134
rect -2698 360898 -2614 361134
rect -2378 360898 -2346 361134
rect -2966 324454 -2346 360898
rect -2966 324218 -2934 324454
rect -2698 324218 -2614 324454
rect -2378 324218 -2346 324454
rect -2966 324134 -2346 324218
rect -2966 323898 -2934 324134
rect -2698 323898 -2614 324134
rect -2378 323898 -2346 324134
rect -2966 287454 -2346 323898
rect -2966 287218 -2934 287454
rect -2698 287218 -2614 287454
rect -2378 287218 -2346 287454
rect -2966 287134 -2346 287218
rect -2966 286898 -2934 287134
rect -2698 286898 -2614 287134
rect -2378 286898 -2346 287134
rect -2966 250454 -2346 286898
rect -2966 250218 -2934 250454
rect -2698 250218 -2614 250454
rect -2378 250218 -2346 250454
rect -2966 250134 -2346 250218
rect -2966 249898 -2934 250134
rect -2698 249898 -2614 250134
rect -2378 249898 -2346 250134
rect -2966 213454 -2346 249898
rect -2966 213218 -2934 213454
rect -2698 213218 -2614 213454
rect -2378 213218 -2346 213454
rect -2966 213134 -2346 213218
rect -2966 212898 -2934 213134
rect -2698 212898 -2614 213134
rect -2378 212898 -2346 213134
rect -2966 176454 -2346 212898
rect -2966 176218 -2934 176454
rect -2698 176218 -2614 176454
rect -2378 176218 -2346 176454
rect -2966 176134 -2346 176218
rect -2966 175898 -2934 176134
rect -2698 175898 -2614 176134
rect -2378 175898 -2346 176134
rect -2966 139454 -2346 175898
rect -2966 139218 -2934 139454
rect -2698 139218 -2614 139454
rect -2378 139218 -2346 139454
rect -2966 139134 -2346 139218
rect -2966 138898 -2934 139134
rect -2698 138898 -2614 139134
rect -2378 138898 -2346 139134
rect -2966 102454 -2346 138898
rect -2966 102218 -2934 102454
rect -2698 102218 -2614 102454
rect -2378 102218 -2346 102454
rect -2966 102134 -2346 102218
rect -2966 101898 -2934 102134
rect -2698 101898 -2614 102134
rect -2378 101898 -2346 102134
rect -2966 65454 -2346 101898
rect -2966 65218 -2934 65454
rect -2698 65218 -2614 65454
rect -2378 65218 -2346 65454
rect -2966 65134 -2346 65218
rect -2966 64898 -2934 65134
rect -2698 64898 -2614 65134
rect -2378 64898 -2346 65134
rect -2966 28454 -2346 64898
rect -2966 28218 -2934 28454
rect -2698 28218 -2614 28454
rect -2378 28218 -2346 28454
rect -2966 28134 -2346 28218
rect -2966 27898 -2934 28134
rect -2698 27898 -2614 28134
rect -2378 27898 -2346 28134
rect -2966 -1306 -2346 27898
rect -2006 704838 -1386 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 -1386 704838
rect -2006 704518 -1386 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 -1386 704518
rect -2006 698174 -1386 704282
rect -2006 697938 -1974 698174
rect -1738 697938 -1654 698174
rect -1418 697938 -1386 698174
rect -2006 697854 -1386 697938
rect -2006 697618 -1974 697854
rect -1738 697618 -1654 697854
rect -1418 697618 -1386 697854
rect -2006 661174 -1386 697618
rect -2006 660938 -1974 661174
rect -1738 660938 -1654 661174
rect -1418 660938 -1386 661174
rect -2006 660854 -1386 660938
rect -2006 660618 -1974 660854
rect -1738 660618 -1654 660854
rect -1418 660618 -1386 660854
rect -2006 624174 -1386 660618
rect -2006 623938 -1974 624174
rect -1738 623938 -1654 624174
rect -1418 623938 -1386 624174
rect -2006 623854 -1386 623938
rect -2006 623618 -1974 623854
rect -1738 623618 -1654 623854
rect -1418 623618 -1386 623854
rect -2006 587174 -1386 623618
rect 37994 694454 38614 705242
rect 37994 694218 38026 694454
rect 38262 694218 38346 694454
rect 38582 694218 38614 694454
rect 37994 694134 38614 694218
rect 37994 693898 38026 694134
rect 38262 693898 38346 694134
rect 38582 693898 38614 694134
rect 37994 657454 38614 693898
rect 37994 657218 38026 657454
rect 38262 657218 38346 657454
rect 38582 657218 38614 657454
rect 37994 657134 38614 657218
rect 37994 656898 38026 657134
rect 38262 656898 38346 657134
rect 38582 656898 38614 657134
rect 37994 620454 38614 656898
rect 37994 620218 38026 620454
rect 38262 620218 38346 620454
rect 38582 620218 38614 620454
rect 37994 620134 38614 620218
rect 37994 619898 38026 620134
rect 38262 619898 38346 620134
rect 38582 619898 38614 620134
rect 3371 606116 3437 606117
rect 3371 606052 3372 606116
rect 3436 606052 3437 606116
rect 3371 606051 3437 606052
rect -2006 586938 -1974 587174
rect -1738 586938 -1654 587174
rect -1418 586938 -1386 587174
rect -2006 586854 -1386 586938
rect -2006 586618 -1974 586854
rect -1738 586618 -1654 586854
rect -1418 586618 -1386 586854
rect -2006 550174 -1386 586618
rect -2006 549938 -1974 550174
rect -1738 549938 -1654 550174
rect -1418 549938 -1386 550174
rect -2006 549854 -1386 549938
rect -2006 549618 -1974 549854
rect -1738 549618 -1654 549854
rect -1418 549618 -1386 549854
rect -2006 513174 -1386 549618
rect -2006 512938 -1974 513174
rect -1738 512938 -1654 513174
rect -1418 512938 -1386 513174
rect -2006 512854 -1386 512938
rect -2006 512618 -1974 512854
rect -1738 512618 -1654 512854
rect -1418 512618 -1386 512854
rect -2006 476174 -1386 512618
rect -2006 475938 -1974 476174
rect -1738 475938 -1654 476174
rect -1418 475938 -1386 476174
rect -2006 475854 -1386 475938
rect -2006 475618 -1974 475854
rect -1738 475618 -1654 475854
rect -1418 475618 -1386 475854
rect -2006 439174 -1386 475618
rect -2006 438938 -1974 439174
rect -1738 438938 -1654 439174
rect -1418 438938 -1386 439174
rect -2006 438854 -1386 438938
rect -2006 438618 -1974 438854
rect -1738 438618 -1654 438854
rect -1418 438618 -1386 438854
rect -2006 402174 -1386 438618
rect -2006 401938 -1974 402174
rect -1738 401938 -1654 402174
rect -1418 401938 -1386 402174
rect -2006 401854 -1386 401938
rect -2006 401618 -1974 401854
rect -1738 401618 -1654 401854
rect -1418 401618 -1386 401854
rect -2006 365174 -1386 401618
rect -2006 364938 -1974 365174
rect -1738 364938 -1654 365174
rect -1418 364938 -1386 365174
rect -2006 364854 -1386 364938
rect -2006 364618 -1974 364854
rect -1738 364618 -1654 364854
rect -1418 364618 -1386 364854
rect -2006 328174 -1386 364618
rect -2006 327938 -1974 328174
rect -1738 327938 -1654 328174
rect -1418 327938 -1386 328174
rect -2006 327854 -1386 327938
rect -2006 327618 -1974 327854
rect -1738 327618 -1654 327854
rect -1418 327618 -1386 327854
rect -2006 291174 -1386 327618
rect -2006 290938 -1974 291174
rect -1738 290938 -1654 291174
rect -1418 290938 -1386 291174
rect -2006 290854 -1386 290938
rect -2006 290618 -1974 290854
rect -1738 290618 -1654 290854
rect -1418 290618 -1386 290854
rect -2006 254174 -1386 290618
rect -2006 253938 -1974 254174
rect -1738 253938 -1654 254174
rect -1418 253938 -1386 254174
rect -2006 253854 -1386 253938
rect -2006 253618 -1974 253854
rect -1738 253618 -1654 253854
rect -1418 253618 -1386 253854
rect -2006 217174 -1386 253618
rect -2006 216938 -1974 217174
rect -1738 216938 -1654 217174
rect -1418 216938 -1386 217174
rect -2006 216854 -1386 216938
rect -2006 216618 -1974 216854
rect -1738 216618 -1654 216854
rect -1418 216618 -1386 216854
rect -2006 180174 -1386 216618
rect -2006 179938 -1974 180174
rect -1738 179938 -1654 180174
rect -1418 179938 -1386 180174
rect -2006 179854 -1386 179938
rect -2006 179618 -1974 179854
rect -1738 179618 -1654 179854
rect -1418 179618 -1386 179854
rect -2006 143174 -1386 179618
rect -2006 142938 -1974 143174
rect -1738 142938 -1654 143174
rect -1418 142938 -1386 143174
rect -2006 142854 -1386 142938
rect -2006 142618 -1974 142854
rect -1738 142618 -1654 142854
rect -1418 142618 -1386 142854
rect -2006 106174 -1386 142618
rect -2006 105938 -1974 106174
rect -1738 105938 -1654 106174
rect -1418 105938 -1386 106174
rect -2006 105854 -1386 105938
rect -2006 105618 -1974 105854
rect -1738 105618 -1654 105854
rect -1418 105618 -1386 105854
rect -2006 69174 -1386 105618
rect -2006 68938 -1974 69174
rect -1738 68938 -1654 69174
rect -1418 68938 -1386 69174
rect -2006 68854 -1386 68938
rect -2006 68618 -1974 68854
rect -1738 68618 -1654 68854
rect -1418 68618 -1386 68854
rect -2006 32174 -1386 68618
rect -2006 31938 -1974 32174
rect -1738 31938 -1654 32174
rect -1418 31938 -1386 32174
rect -2006 31854 -1386 31938
rect -2006 31618 -1974 31854
rect -1738 31618 -1654 31854
rect -1418 31618 -1386 31854
rect -2006 -346 -1386 31618
rect 3374 17645 3434 606051
rect 37994 583454 38614 619898
rect 37994 583218 38026 583454
rect 38262 583218 38346 583454
rect 38582 583218 38614 583454
rect 37994 583134 38614 583218
rect 37994 582898 38026 583134
rect 38262 582898 38346 583134
rect 38582 582898 38614 583134
rect 3555 580004 3621 580005
rect 3555 579940 3556 580004
rect 3620 579940 3621 580004
rect 3555 579939 3621 579940
rect 3371 17644 3437 17645
rect 3371 17580 3372 17644
rect 3436 17580 3437 17644
rect 3371 17579 3437 17580
rect 3558 17509 3618 579939
rect 37994 546454 38614 582898
rect 37994 546218 38026 546454
rect 38262 546218 38346 546454
rect 38582 546218 38614 546454
rect 37994 546134 38614 546218
rect 37994 545898 38026 546134
rect 38262 545898 38346 546134
rect 38582 545898 38614 546134
rect 37994 509454 38614 545898
rect 37994 509218 38026 509454
rect 38262 509218 38346 509454
rect 38582 509218 38614 509454
rect 37994 509134 38614 509218
rect 37994 508898 38026 509134
rect 38262 508898 38346 509134
rect 38582 508898 38614 509134
rect 3739 501804 3805 501805
rect 3739 501740 3740 501804
rect 3804 501740 3805 501804
rect 3739 501739 3805 501740
rect 3742 17781 3802 501739
rect 3923 475692 3989 475693
rect 3923 475628 3924 475692
rect 3988 475628 3989 475692
rect 3923 475627 3989 475628
rect 3739 17780 3805 17781
rect 3739 17716 3740 17780
rect 3804 17716 3805 17780
rect 3739 17715 3805 17716
rect 3555 17508 3621 17509
rect 3555 17444 3556 17508
rect 3620 17444 3621 17508
rect 3555 17443 3621 17444
rect 3926 17373 3986 475627
rect 37994 472454 38614 508898
rect 37994 472218 38026 472454
rect 38262 472218 38346 472454
rect 38582 472218 38614 472454
rect 37994 472134 38614 472218
rect 37994 471898 38026 472134
rect 38262 471898 38346 472134
rect 38582 471898 38614 472134
rect 37994 435454 38614 471898
rect 37994 435218 38026 435454
rect 38262 435218 38346 435454
rect 38582 435218 38614 435454
rect 37994 435134 38614 435218
rect 37994 434898 38026 435134
rect 38262 434898 38346 435134
rect 38582 434898 38614 435134
rect 37994 398454 38614 434898
rect 37994 398218 38026 398454
rect 38262 398218 38346 398454
rect 38582 398218 38614 398454
rect 37994 398134 38614 398218
rect 37994 397898 38026 398134
rect 38262 397898 38346 398134
rect 38582 397898 38614 398134
rect 37994 361454 38614 397898
rect 37994 361218 38026 361454
rect 38262 361218 38346 361454
rect 38582 361218 38614 361454
rect 37994 361134 38614 361218
rect 37994 360898 38026 361134
rect 38262 360898 38346 361134
rect 38582 360898 38614 361134
rect 21955 325276 22021 325277
rect 21955 325212 21956 325276
rect 22020 325212 22021 325276
rect 21955 325211 22021 325212
rect 21958 20637 22018 325211
rect 37994 324454 38614 360898
rect 37994 324218 38026 324454
rect 38262 324218 38346 324454
rect 38582 324218 38614 324454
rect 37994 324134 38614 324218
rect 37994 323898 38026 324134
rect 38262 323898 38346 324134
rect 38582 323898 38614 324134
rect 37994 287454 38614 323898
rect 37994 287218 38026 287454
rect 38262 287218 38346 287454
rect 38582 287218 38614 287454
rect 37994 287134 38614 287218
rect 37994 286898 38026 287134
rect 38262 286898 38346 287134
rect 38582 286898 38614 287134
rect 37994 250454 38614 286898
rect 37994 250218 38026 250454
rect 38262 250218 38346 250454
rect 38582 250218 38614 250454
rect 37994 250134 38614 250218
rect 37994 249898 38026 250134
rect 38262 249898 38346 250134
rect 38582 249898 38614 250134
rect 37994 213454 38614 249898
rect 37994 213218 38026 213454
rect 38262 213218 38346 213454
rect 38582 213218 38614 213454
rect 37994 213134 38614 213218
rect 37994 212898 38026 213134
rect 38262 212898 38346 213134
rect 38582 212898 38614 213134
rect 37994 176454 38614 212898
rect 37994 176218 38026 176454
rect 38262 176218 38346 176454
rect 38582 176218 38614 176454
rect 37994 176134 38614 176218
rect 37994 175898 38026 176134
rect 38262 175898 38346 176134
rect 38582 175898 38614 176134
rect 37994 139454 38614 175898
rect 37994 139218 38026 139454
rect 38262 139218 38346 139454
rect 38582 139218 38614 139454
rect 37994 139134 38614 139218
rect 37994 138898 38026 139134
rect 38262 138898 38346 139134
rect 38582 138898 38614 139134
rect 37994 102454 38614 138898
rect 37994 102218 38026 102454
rect 38262 102218 38346 102454
rect 38582 102218 38614 102454
rect 37994 102134 38614 102218
rect 37994 101898 38026 102134
rect 38262 101898 38346 102134
rect 38582 101898 38614 102134
rect 37994 65454 38614 101898
rect 37994 65218 38026 65454
rect 38262 65218 38346 65454
rect 38582 65218 38614 65454
rect 37994 65134 38614 65218
rect 37994 64898 38026 65134
rect 38262 64898 38346 65134
rect 38582 64898 38614 65134
rect 26418 32174 26738 32206
rect 26418 31938 26460 32174
rect 26696 31938 26738 32174
rect 26418 31854 26738 31938
rect 26418 31618 26460 31854
rect 26696 31618 26738 31854
rect 26418 31586 26738 31618
rect 37366 32174 37686 32206
rect 37366 31938 37408 32174
rect 37644 31938 37686 32174
rect 37366 31854 37686 31938
rect 37366 31618 37408 31854
rect 37644 31618 37686 31854
rect 37366 31586 37686 31618
rect 31892 28454 32212 28486
rect 31892 28218 31934 28454
rect 32170 28218 32212 28454
rect 31892 28134 32212 28218
rect 31892 27898 31934 28134
rect 32170 27898 32212 28134
rect 31892 27866 32212 27898
rect 37994 28454 38614 64898
rect 37994 28218 38026 28454
rect 38262 28218 38346 28454
rect 38582 28218 38614 28454
rect 37994 28134 38614 28218
rect 37994 27898 38026 28134
rect 38262 27898 38346 28134
rect 38582 27898 38614 28134
rect 21955 20636 22021 20637
rect 21955 20572 21956 20636
rect 22020 20572 22021 20636
rect 21955 20571 22021 20572
rect 3923 17372 3989 17373
rect 3923 17308 3924 17372
rect 3988 17308 3989 17372
rect 3923 17307 3989 17308
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 -1386 -346
rect -2006 -666 -1386 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 -1386 -666
rect -2006 -934 -1386 -902
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 -2346 -1306
rect -2966 -1626 -2346 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 -2346 -1626
rect -2966 -1894 -2346 -1862
rect 37994 -1306 38614 27898
rect 37994 -1542 38026 -1306
rect 38262 -1542 38346 -1306
rect 38582 -1542 38614 -1306
rect 37994 -1626 38614 -1542
rect 37994 -1862 38026 -1626
rect 38262 -1862 38346 -1626
rect 38582 -1862 38614 -1626
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 -3306 -2266
rect -3926 -2586 -3306 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 -3306 -2586
rect -3926 -2854 -3306 -2822
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 -4266 -3226
rect -4886 -3546 -4266 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 -4266 -3546
rect -4886 -3814 -4266 -3782
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 -5226 -4186
rect -5846 -4506 -5226 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 -5226 -4506
rect -5846 -4774 -5226 -4742
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 -6186 -5146
rect -6806 -5466 -6186 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 -6186 -5466
rect -6806 -5734 -6186 -5702
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 -7146 -6106
rect -7766 -6426 -7146 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 -7146 -6426
rect -7766 -6694 -7146 -6662
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 -8106 -7066
rect -8726 -7386 -8106 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 -8106 -7386
rect -8726 -7654 -8106 -7622
rect 37994 -7654 38614 -1862
rect 41714 704838 42334 711590
rect 41714 704602 41746 704838
rect 41982 704602 42066 704838
rect 42302 704602 42334 704838
rect 41714 704518 42334 704602
rect 41714 704282 41746 704518
rect 41982 704282 42066 704518
rect 42302 704282 42334 704518
rect 41714 698174 42334 704282
rect 41714 697938 41746 698174
rect 41982 697938 42066 698174
rect 42302 697938 42334 698174
rect 41714 697854 42334 697938
rect 41714 697618 41746 697854
rect 41982 697618 42066 697854
rect 42302 697618 42334 697854
rect 41714 661174 42334 697618
rect 41714 660938 41746 661174
rect 41982 660938 42066 661174
rect 42302 660938 42334 661174
rect 41714 660854 42334 660938
rect 41714 660618 41746 660854
rect 41982 660618 42066 660854
rect 42302 660618 42334 660854
rect 41714 624174 42334 660618
rect 41714 623938 41746 624174
rect 41982 623938 42066 624174
rect 42302 623938 42334 624174
rect 41714 623854 42334 623938
rect 41714 623618 41746 623854
rect 41982 623618 42066 623854
rect 42302 623618 42334 623854
rect 41714 587174 42334 623618
rect 41714 586938 41746 587174
rect 41982 586938 42066 587174
rect 42302 586938 42334 587174
rect 41714 586854 42334 586938
rect 41714 586618 41746 586854
rect 41982 586618 42066 586854
rect 42302 586618 42334 586854
rect 41714 550174 42334 586618
rect 41714 549938 41746 550174
rect 41982 549938 42066 550174
rect 42302 549938 42334 550174
rect 41714 549854 42334 549938
rect 41714 549618 41746 549854
rect 41982 549618 42066 549854
rect 42302 549618 42334 549854
rect 41714 513174 42334 549618
rect 41714 512938 41746 513174
rect 41982 512938 42066 513174
rect 42302 512938 42334 513174
rect 41714 512854 42334 512938
rect 41714 512618 41746 512854
rect 41982 512618 42066 512854
rect 42302 512618 42334 512854
rect 41714 476174 42334 512618
rect 41714 475938 41746 476174
rect 41982 475938 42066 476174
rect 42302 475938 42334 476174
rect 41714 475854 42334 475938
rect 41714 475618 41746 475854
rect 41982 475618 42066 475854
rect 42302 475618 42334 475854
rect 41714 439174 42334 475618
rect 41714 438938 41746 439174
rect 41982 438938 42066 439174
rect 42302 438938 42334 439174
rect 41714 438854 42334 438938
rect 41714 438618 41746 438854
rect 41982 438618 42066 438854
rect 42302 438618 42334 438854
rect 41714 402174 42334 438618
rect 41714 401938 41746 402174
rect 41982 401938 42066 402174
rect 42302 401938 42334 402174
rect 41714 401854 42334 401938
rect 41714 401618 41746 401854
rect 41982 401618 42066 401854
rect 42302 401618 42334 401854
rect 41714 365174 42334 401618
rect 41714 364938 41746 365174
rect 41982 364938 42066 365174
rect 42302 364938 42334 365174
rect 41714 364854 42334 364938
rect 41714 364618 41746 364854
rect 41982 364618 42066 364854
rect 42302 364618 42334 364854
rect 41714 328174 42334 364618
rect 41714 327938 41746 328174
rect 41982 327938 42066 328174
rect 42302 327938 42334 328174
rect 41714 327854 42334 327938
rect 41714 327618 41746 327854
rect 41982 327618 42066 327854
rect 42302 327618 42334 327854
rect 41714 291174 42334 327618
rect 41714 290938 41746 291174
rect 41982 290938 42066 291174
rect 42302 290938 42334 291174
rect 41714 290854 42334 290938
rect 41714 290618 41746 290854
rect 41982 290618 42066 290854
rect 42302 290618 42334 290854
rect 41714 254174 42334 290618
rect 41714 253938 41746 254174
rect 41982 253938 42066 254174
rect 42302 253938 42334 254174
rect 41714 253854 42334 253938
rect 41714 253618 41746 253854
rect 41982 253618 42066 253854
rect 42302 253618 42334 253854
rect 41714 217174 42334 253618
rect 41714 216938 41746 217174
rect 41982 216938 42066 217174
rect 42302 216938 42334 217174
rect 41714 216854 42334 216938
rect 41714 216618 41746 216854
rect 41982 216618 42066 216854
rect 42302 216618 42334 216854
rect 41714 180174 42334 216618
rect 41714 179938 41746 180174
rect 41982 179938 42066 180174
rect 42302 179938 42334 180174
rect 41714 179854 42334 179938
rect 41714 179618 41746 179854
rect 41982 179618 42066 179854
rect 42302 179618 42334 179854
rect 41714 143174 42334 179618
rect 41714 142938 41746 143174
rect 41982 142938 42066 143174
rect 42302 142938 42334 143174
rect 41714 142854 42334 142938
rect 41714 142618 41746 142854
rect 41982 142618 42066 142854
rect 42302 142618 42334 142854
rect 41714 106174 42334 142618
rect 41714 105938 41746 106174
rect 41982 105938 42066 106174
rect 42302 105938 42334 106174
rect 41714 105854 42334 105938
rect 41714 105618 41746 105854
rect 41982 105618 42066 105854
rect 42302 105618 42334 105854
rect 41714 69174 42334 105618
rect 41714 68938 41746 69174
rect 41982 68938 42066 69174
rect 42302 68938 42334 69174
rect 41714 68854 42334 68938
rect 41714 68618 41746 68854
rect 41982 68618 42066 68854
rect 42302 68618 42334 68854
rect 41714 32174 42334 68618
rect 65994 705798 66614 711590
rect 65994 705562 66026 705798
rect 66262 705562 66346 705798
rect 66582 705562 66614 705798
rect 65994 705478 66614 705562
rect 65994 705242 66026 705478
rect 66262 705242 66346 705478
rect 66582 705242 66614 705478
rect 65994 694454 66614 705242
rect 65994 694218 66026 694454
rect 66262 694218 66346 694454
rect 66582 694218 66614 694454
rect 65994 694134 66614 694218
rect 65994 693898 66026 694134
rect 66262 693898 66346 694134
rect 66582 693898 66614 694134
rect 65994 657454 66614 693898
rect 65994 657218 66026 657454
rect 66262 657218 66346 657454
rect 66582 657218 66614 657454
rect 65994 657134 66614 657218
rect 65994 656898 66026 657134
rect 66262 656898 66346 657134
rect 66582 656898 66614 657134
rect 65994 620454 66614 656898
rect 65994 620218 66026 620454
rect 66262 620218 66346 620454
rect 66582 620218 66614 620454
rect 65994 620134 66614 620218
rect 65994 619898 66026 620134
rect 66262 619898 66346 620134
rect 66582 619898 66614 620134
rect 65994 583454 66614 619898
rect 65994 583218 66026 583454
rect 66262 583218 66346 583454
rect 66582 583218 66614 583454
rect 65994 583134 66614 583218
rect 65994 582898 66026 583134
rect 66262 582898 66346 583134
rect 66582 582898 66614 583134
rect 65994 546454 66614 582898
rect 65994 546218 66026 546454
rect 66262 546218 66346 546454
rect 66582 546218 66614 546454
rect 65994 546134 66614 546218
rect 65994 545898 66026 546134
rect 66262 545898 66346 546134
rect 66582 545898 66614 546134
rect 65994 509454 66614 545898
rect 65994 509218 66026 509454
rect 66262 509218 66346 509454
rect 66582 509218 66614 509454
rect 65994 509134 66614 509218
rect 65994 508898 66026 509134
rect 66262 508898 66346 509134
rect 66582 508898 66614 509134
rect 65994 472454 66614 508898
rect 65994 472218 66026 472454
rect 66262 472218 66346 472454
rect 66582 472218 66614 472454
rect 65994 472134 66614 472218
rect 65994 471898 66026 472134
rect 66262 471898 66346 472134
rect 66582 471898 66614 472134
rect 65994 435454 66614 471898
rect 65994 435218 66026 435454
rect 66262 435218 66346 435454
rect 66582 435218 66614 435454
rect 65994 435134 66614 435218
rect 65994 434898 66026 435134
rect 66262 434898 66346 435134
rect 66582 434898 66614 435134
rect 65994 398454 66614 434898
rect 65994 398218 66026 398454
rect 66262 398218 66346 398454
rect 66582 398218 66614 398454
rect 65994 398134 66614 398218
rect 65994 397898 66026 398134
rect 66262 397898 66346 398134
rect 66582 397898 66614 398134
rect 65994 361454 66614 397898
rect 65994 361218 66026 361454
rect 66262 361218 66346 361454
rect 66582 361218 66614 361454
rect 65994 361134 66614 361218
rect 65994 360898 66026 361134
rect 66262 360898 66346 361134
rect 66582 360898 66614 361134
rect 65994 324454 66614 360898
rect 65994 324218 66026 324454
rect 66262 324218 66346 324454
rect 66582 324218 66614 324454
rect 65994 324134 66614 324218
rect 65994 323898 66026 324134
rect 66262 323898 66346 324134
rect 66582 323898 66614 324134
rect 65994 287454 66614 323898
rect 65994 287218 66026 287454
rect 66262 287218 66346 287454
rect 66582 287218 66614 287454
rect 65994 287134 66614 287218
rect 65994 286898 66026 287134
rect 66262 286898 66346 287134
rect 66582 286898 66614 287134
rect 65994 250454 66614 286898
rect 65994 250218 66026 250454
rect 66262 250218 66346 250454
rect 66582 250218 66614 250454
rect 65994 250134 66614 250218
rect 65994 249898 66026 250134
rect 66262 249898 66346 250134
rect 66582 249898 66614 250134
rect 65994 213454 66614 249898
rect 65994 213218 66026 213454
rect 66262 213218 66346 213454
rect 66582 213218 66614 213454
rect 65994 213134 66614 213218
rect 65994 212898 66026 213134
rect 66262 212898 66346 213134
rect 66582 212898 66614 213134
rect 65994 176454 66614 212898
rect 65994 176218 66026 176454
rect 66262 176218 66346 176454
rect 66582 176218 66614 176454
rect 65994 176134 66614 176218
rect 65994 175898 66026 176134
rect 66262 175898 66346 176134
rect 66582 175898 66614 176134
rect 65994 139454 66614 175898
rect 65994 139218 66026 139454
rect 66262 139218 66346 139454
rect 66582 139218 66614 139454
rect 65994 139134 66614 139218
rect 65994 138898 66026 139134
rect 66262 138898 66346 139134
rect 66582 138898 66614 139134
rect 65994 102454 66614 138898
rect 65994 102218 66026 102454
rect 66262 102218 66346 102454
rect 66582 102218 66614 102454
rect 65994 102134 66614 102218
rect 65994 101898 66026 102134
rect 66262 101898 66346 102134
rect 66582 101898 66614 102134
rect 65994 65454 66614 101898
rect 65994 65218 66026 65454
rect 66262 65218 66346 65454
rect 66582 65218 66614 65454
rect 65994 65134 66614 65218
rect 65994 64898 66026 65134
rect 66262 64898 66346 65134
rect 66582 64898 66614 65134
rect 44035 39404 44101 39405
rect 44035 39340 44036 39404
rect 44100 39340 44101 39404
rect 44035 39339 44101 39340
rect 46979 39404 47045 39405
rect 46979 39340 46980 39404
rect 47044 39340 47045 39404
rect 46979 39339 47045 39340
rect 55075 39404 55141 39405
rect 55075 39340 55076 39404
rect 55140 39340 55141 39404
rect 55075 39339 55141 39340
rect 41714 31938 41746 32174
rect 41982 31938 42066 32174
rect 42302 31938 42334 32174
rect 41714 31854 42334 31938
rect 41714 31618 41746 31854
rect 41982 31618 42066 31854
rect 42302 31618 42334 31854
rect 41714 -346 42334 31618
rect 42840 28454 43160 28486
rect 42840 28218 42882 28454
rect 43118 28218 43160 28454
rect 42840 28134 43160 28218
rect 42840 27898 42882 28134
rect 43118 27898 43160 28134
rect 42840 27866 43160 27898
rect 44038 3365 44098 39339
rect 46982 6493 47042 39339
rect 48314 32174 48634 32206
rect 48314 31938 48356 32174
rect 48592 31938 48634 32174
rect 48314 31854 48634 31938
rect 48314 31618 48356 31854
rect 48592 31618 48634 31854
rect 48314 31586 48634 31618
rect 53788 28454 54108 28486
rect 53788 28218 53830 28454
rect 54066 28218 54108 28454
rect 53788 28134 54108 28218
rect 53788 27898 53830 28134
rect 54066 27898 54108 28134
rect 53788 27866 54108 27898
rect 46979 6492 47045 6493
rect 46979 6428 46980 6492
rect 47044 6428 47045 6492
rect 46979 6427 47045 6428
rect 55078 3501 55138 39339
rect 60595 39268 60661 39269
rect 60595 39204 60596 39268
rect 60660 39204 60661 39268
rect 60595 39203 60661 39204
rect 59262 32174 59582 32206
rect 59262 31938 59304 32174
rect 59540 31938 59582 32174
rect 59262 31854 59582 31938
rect 59262 31618 59304 31854
rect 59540 31618 59582 31854
rect 59262 31586 59582 31618
rect 60598 20501 60658 39203
rect 64736 28454 65056 28486
rect 64736 28218 64778 28454
rect 65014 28218 65056 28454
rect 64736 28134 65056 28218
rect 64736 27898 64778 28134
rect 65014 27898 65056 28134
rect 64736 27866 65056 27898
rect 65994 28454 66614 64898
rect 65994 28218 66026 28454
rect 66262 28218 66346 28454
rect 66582 28218 66614 28454
rect 65994 28134 66614 28218
rect 65994 27898 66026 28134
rect 66262 27898 66346 28134
rect 66582 27898 66614 28134
rect 60595 20500 60661 20501
rect 60595 20436 60596 20500
rect 60660 20436 60661 20500
rect 60595 20435 60661 20436
rect 55075 3500 55141 3501
rect 55075 3436 55076 3500
rect 55140 3436 55141 3500
rect 55075 3435 55141 3436
rect 44035 3364 44101 3365
rect 44035 3300 44036 3364
rect 44100 3300 44101 3364
rect 44035 3299 44101 3300
rect 41714 -582 41746 -346
rect 41982 -582 42066 -346
rect 42302 -582 42334 -346
rect 41714 -666 42334 -582
rect 41714 -902 41746 -666
rect 41982 -902 42066 -666
rect 42302 -902 42334 -666
rect 41714 -7654 42334 -902
rect 65994 -1306 66614 27898
rect 65994 -1542 66026 -1306
rect 66262 -1542 66346 -1306
rect 66582 -1542 66614 -1306
rect 65994 -1626 66614 -1542
rect 65994 -1862 66026 -1626
rect 66262 -1862 66346 -1626
rect 66582 -1862 66614 -1626
rect 65994 -7654 66614 -1862
rect 69714 704838 70334 711590
rect 69714 704602 69746 704838
rect 69982 704602 70066 704838
rect 70302 704602 70334 704838
rect 69714 704518 70334 704602
rect 69714 704282 69746 704518
rect 69982 704282 70066 704518
rect 70302 704282 70334 704518
rect 69714 698174 70334 704282
rect 69714 697938 69746 698174
rect 69982 697938 70066 698174
rect 70302 697938 70334 698174
rect 69714 697854 70334 697938
rect 69714 697618 69746 697854
rect 69982 697618 70066 697854
rect 70302 697618 70334 697854
rect 69714 661174 70334 697618
rect 69714 660938 69746 661174
rect 69982 660938 70066 661174
rect 70302 660938 70334 661174
rect 69714 660854 70334 660938
rect 69714 660618 69746 660854
rect 69982 660618 70066 660854
rect 70302 660618 70334 660854
rect 69714 624174 70334 660618
rect 69714 623938 69746 624174
rect 69982 623938 70066 624174
rect 70302 623938 70334 624174
rect 69714 623854 70334 623938
rect 69714 623618 69746 623854
rect 69982 623618 70066 623854
rect 70302 623618 70334 623854
rect 69714 587174 70334 623618
rect 69714 586938 69746 587174
rect 69982 586938 70066 587174
rect 70302 586938 70334 587174
rect 69714 586854 70334 586938
rect 69714 586618 69746 586854
rect 69982 586618 70066 586854
rect 70302 586618 70334 586854
rect 69714 550174 70334 586618
rect 69714 549938 69746 550174
rect 69982 549938 70066 550174
rect 70302 549938 70334 550174
rect 69714 549854 70334 549938
rect 69714 549618 69746 549854
rect 69982 549618 70066 549854
rect 70302 549618 70334 549854
rect 69714 513174 70334 549618
rect 69714 512938 69746 513174
rect 69982 512938 70066 513174
rect 70302 512938 70334 513174
rect 69714 512854 70334 512938
rect 69714 512618 69746 512854
rect 69982 512618 70066 512854
rect 70302 512618 70334 512854
rect 69714 476174 70334 512618
rect 69714 475938 69746 476174
rect 69982 475938 70066 476174
rect 70302 475938 70334 476174
rect 69714 475854 70334 475938
rect 69714 475618 69746 475854
rect 69982 475618 70066 475854
rect 70302 475618 70334 475854
rect 69714 439174 70334 475618
rect 69714 438938 69746 439174
rect 69982 438938 70066 439174
rect 70302 438938 70334 439174
rect 69714 438854 70334 438938
rect 69714 438618 69746 438854
rect 69982 438618 70066 438854
rect 70302 438618 70334 438854
rect 69714 402174 70334 438618
rect 69714 401938 69746 402174
rect 69982 401938 70066 402174
rect 70302 401938 70334 402174
rect 69714 401854 70334 401938
rect 69714 401618 69746 401854
rect 69982 401618 70066 401854
rect 70302 401618 70334 401854
rect 69714 365174 70334 401618
rect 69714 364938 69746 365174
rect 69982 364938 70066 365174
rect 70302 364938 70334 365174
rect 69714 364854 70334 364938
rect 69714 364618 69746 364854
rect 69982 364618 70066 364854
rect 70302 364618 70334 364854
rect 69714 328174 70334 364618
rect 69714 327938 69746 328174
rect 69982 327938 70066 328174
rect 70302 327938 70334 328174
rect 69714 327854 70334 327938
rect 69714 327618 69746 327854
rect 69982 327618 70066 327854
rect 70302 327618 70334 327854
rect 69714 291174 70334 327618
rect 69714 290938 69746 291174
rect 69982 290938 70066 291174
rect 70302 290938 70334 291174
rect 69714 290854 70334 290938
rect 69714 290618 69746 290854
rect 69982 290618 70066 290854
rect 70302 290618 70334 290854
rect 69714 254174 70334 290618
rect 69714 253938 69746 254174
rect 69982 253938 70066 254174
rect 70302 253938 70334 254174
rect 69714 253854 70334 253938
rect 69714 253618 69746 253854
rect 69982 253618 70066 253854
rect 70302 253618 70334 253854
rect 69714 217174 70334 253618
rect 69714 216938 69746 217174
rect 69982 216938 70066 217174
rect 70302 216938 70334 217174
rect 69714 216854 70334 216938
rect 69714 216618 69746 216854
rect 69982 216618 70066 216854
rect 70302 216618 70334 216854
rect 69714 180174 70334 216618
rect 69714 179938 69746 180174
rect 69982 179938 70066 180174
rect 70302 179938 70334 180174
rect 69714 179854 70334 179938
rect 69714 179618 69746 179854
rect 69982 179618 70066 179854
rect 70302 179618 70334 179854
rect 69714 143174 70334 179618
rect 69714 142938 69746 143174
rect 69982 142938 70066 143174
rect 70302 142938 70334 143174
rect 69714 142854 70334 142938
rect 69714 142618 69746 142854
rect 69982 142618 70066 142854
rect 70302 142618 70334 142854
rect 69714 106174 70334 142618
rect 69714 105938 69746 106174
rect 69982 105938 70066 106174
rect 70302 105938 70334 106174
rect 69714 105854 70334 105938
rect 69714 105618 69746 105854
rect 69982 105618 70066 105854
rect 70302 105618 70334 105854
rect 69714 69174 70334 105618
rect 69714 68938 69746 69174
rect 69982 68938 70066 69174
rect 70302 68938 70334 69174
rect 69714 68854 70334 68938
rect 69714 68618 69746 68854
rect 69982 68618 70066 68854
rect 70302 68618 70334 68854
rect 69714 32174 70334 68618
rect 93994 705798 94614 711590
rect 93994 705562 94026 705798
rect 94262 705562 94346 705798
rect 94582 705562 94614 705798
rect 93994 705478 94614 705562
rect 93994 705242 94026 705478
rect 94262 705242 94346 705478
rect 94582 705242 94614 705478
rect 93994 694454 94614 705242
rect 93994 694218 94026 694454
rect 94262 694218 94346 694454
rect 94582 694218 94614 694454
rect 93994 694134 94614 694218
rect 93994 693898 94026 694134
rect 94262 693898 94346 694134
rect 94582 693898 94614 694134
rect 93994 657454 94614 693898
rect 93994 657218 94026 657454
rect 94262 657218 94346 657454
rect 94582 657218 94614 657454
rect 93994 657134 94614 657218
rect 93994 656898 94026 657134
rect 94262 656898 94346 657134
rect 94582 656898 94614 657134
rect 93994 620454 94614 656898
rect 93994 620218 94026 620454
rect 94262 620218 94346 620454
rect 94582 620218 94614 620454
rect 93994 620134 94614 620218
rect 93994 619898 94026 620134
rect 94262 619898 94346 620134
rect 94582 619898 94614 620134
rect 93994 583454 94614 619898
rect 93994 583218 94026 583454
rect 94262 583218 94346 583454
rect 94582 583218 94614 583454
rect 93994 583134 94614 583218
rect 93994 582898 94026 583134
rect 94262 582898 94346 583134
rect 94582 582898 94614 583134
rect 93994 546454 94614 582898
rect 93994 546218 94026 546454
rect 94262 546218 94346 546454
rect 94582 546218 94614 546454
rect 93994 546134 94614 546218
rect 93994 545898 94026 546134
rect 94262 545898 94346 546134
rect 94582 545898 94614 546134
rect 93994 509454 94614 545898
rect 93994 509218 94026 509454
rect 94262 509218 94346 509454
rect 94582 509218 94614 509454
rect 93994 509134 94614 509218
rect 93994 508898 94026 509134
rect 94262 508898 94346 509134
rect 94582 508898 94614 509134
rect 93994 472454 94614 508898
rect 93994 472218 94026 472454
rect 94262 472218 94346 472454
rect 94582 472218 94614 472454
rect 93994 472134 94614 472218
rect 93994 471898 94026 472134
rect 94262 471898 94346 472134
rect 94582 471898 94614 472134
rect 93994 435454 94614 471898
rect 93994 435218 94026 435454
rect 94262 435218 94346 435454
rect 94582 435218 94614 435454
rect 93994 435134 94614 435218
rect 93994 434898 94026 435134
rect 94262 434898 94346 435134
rect 94582 434898 94614 435134
rect 93994 398454 94614 434898
rect 93994 398218 94026 398454
rect 94262 398218 94346 398454
rect 94582 398218 94614 398454
rect 93994 398134 94614 398218
rect 93994 397898 94026 398134
rect 94262 397898 94346 398134
rect 94582 397898 94614 398134
rect 93994 361454 94614 397898
rect 93994 361218 94026 361454
rect 94262 361218 94346 361454
rect 94582 361218 94614 361454
rect 93994 361134 94614 361218
rect 93994 360898 94026 361134
rect 94262 360898 94346 361134
rect 94582 360898 94614 361134
rect 93994 324454 94614 360898
rect 93994 324218 94026 324454
rect 94262 324218 94346 324454
rect 94582 324218 94614 324454
rect 93994 324134 94614 324218
rect 93994 323898 94026 324134
rect 94262 323898 94346 324134
rect 94582 323898 94614 324134
rect 93994 287454 94614 323898
rect 93994 287218 94026 287454
rect 94262 287218 94346 287454
rect 94582 287218 94614 287454
rect 93994 287134 94614 287218
rect 93994 286898 94026 287134
rect 94262 286898 94346 287134
rect 94582 286898 94614 287134
rect 93994 250454 94614 286898
rect 93994 250218 94026 250454
rect 94262 250218 94346 250454
rect 94582 250218 94614 250454
rect 93994 250134 94614 250218
rect 93994 249898 94026 250134
rect 94262 249898 94346 250134
rect 94582 249898 94614 250134
rect 93994 213454 94614 249898
rect 93994 213218 94026 213454
rect 94262 213218 94346 213454
rect 94582 213218 94614 213454
rect 93994 213134 94614 213218
rect 93994 212898 94026 213134
rect 94262 212898 94346 213134
rect 94582 212898 94614 213134
rect 93994 176454 94614 212898
rect 93994 176218 94026 176454
rect 94262 176218 94346 176454
rect 94582 176218 94614 176454
rect 93994 176134 94614 176218
rect 93994 175898 94026 176134
rect 94262 175898 94346 176134
rect 94582 175898 94614 176134
rect 93994 139454 94614 175898
rect 93994 139218 94026 139454
rect 94262 139218 94346 139454
rect 94582 139218 94614 139454
rect 93994 139134 94614 139218
rect 93994 138898 94026 139134
rect 94262 138898 94346 139134
rect 94582 138898 94614 139134
rect 93994 102454 94614 138898
rect 93994 102218 94026 102454
rect 94262 102218 94346 102454
rect 94582 102218 94614 102454
rect 93994 102134 94614 102218
rect 93994 101898 94026 102134
rect 94262 101898 94346 102134
rect 94582 101898 94614 102134
rect 93994 65454 94614 101898
rect 93994 65218 94026 65454
rect 94262 65218 94346 65454
rect 94582 65218 94614 65454
rect 93994 65134 94614 65218
rect 93994 64898 94026 65134
rect 94262 64898 94346 65134
rect 94582 64898 94614 65134
rect 93994 43956 94614 64898
rect 97714 704838 98334 711590
rect 97714 704602 97746 704838
rect 97982 704602 98066 704838
rect 98302 704602 98334 704838
rect 97714 704518 98334 704602
rect 97714 704282 97746 704518
rect 97982 704282 98066 704518
rect 98302 704282 98334 704518
rect 97714 698174 98334 704282
rect 97714 697938 97746 698174
rect 97982 697938 98066 698174
rect 98302 697938 98334 698174
rect 97714 697854 98334 697938
rect 97714 697618 97746 697854
rect 97982 697618 98066 697854
rect 98302 697618 98334 697854
rect 97714 661174 98334 697618
rect 97714 660938 97746 661174
rect 97982 660938 98066 661174
rect 98302 660938 98334 661174
rect 97714 660854 98334 660938
rect 97714 660618 97746 660854
rect 97982 660618 98066 660854
rect 98302 660618 98334 660854
rect 97714 624174 98334 660618
rect 97714 623938 97746 624174
rect 97982 623938 98066 624174
rect 98302 623938 98334 624174
rect 97714 623854 98334 623938
rect 97714 623618 97746 623854
rect 97982 623618 98066 623854
rect 98302 623618 98334 623854
rect 97714 587174 98334 623618
rect 97714 586938 97746 587174
rect 97982 586938 98066 587174
rect 98302 586938 98334 587174
rect 97714 586854 98334 586938
rect 97714 586618 97746 586854
rect 97982 586618 98066 586854
rect 98302 586618 98334 586854
rect 97714 550174 98334 586618
rect 97714 549938 97746 550174
rect 97982 549938 98066 550174
rect 98302 549938 98334 550174
rect 97714 549854 98334 549938
rect 97714 549618 97746 549854
rect 97982 549618 98066 549854
rect 98302 549618 98334 549854
rect 97714 513174 98334 549618
rect 97714 512938 97746 513174
rect 97982 512938 98066 513174
rect 98302 512938 98334 513174
rect 97714 512854 98334 512938
rect 97714 512618 97746 512854
rect 97982 512618 98066 512854
rect 98302 512618 98334 512854
rect 97714 476174 98334 512618
rect 97714 475938 97746 476174
rect 97982 475938 98066 476174
rect 98302 475938 98334 476174
rect 97714 475854 98334 475938
rect 97714 475618 97746 475854
rect 97982 475618 98066 475854
rect 98302 475618 98334 475854
rect 97714 439174 98334 475618
rect 97714 438938 97746 439174
rect 97982 438938 98066 439174
rect 98302 438938 98334 439174
rect 97714 438854 98334 438938
rect 97714 438618 97746 438854
rect 97982 438618 98066 438854
rect 98302 438618 98334 438854
rect 97714 402174 98334 438618
rect 97714 401938 97746 402174
rect 97982 401938 98066 402174
rect 98302 401938 98334 402174
rect 97714 401854 98334 401938
rect 97714 401618 97746 401854
rect 97982 401618 98066 401854
rect 98302 401618 98334 401854
rect 97714 365174 98334 401618
rect 97714 364938 97746 365174
rect 97982 364938 98066 365174
rect 98302 364938 98334 365174
rect 97714 364854 98334 364938
rect 97714 364618 97746 364854
rect 97982 364618 98066 364854
rect 98302 364618 98334 364854
rect 97714 328174 98334 364618
rect 97714 327938 97746 328174
rect 97982 327938 98066 328174
rect 98302 327938 98334 328174
rect 97714 327854 98334 327938
rect 97714 327618 97746 327854
rect 97982 327618 98066 327854
rect 98302 327618 98334 327854
rect 97714 291174 98334 327618
rect 97714 290938 97746 291174
rect 97982 290938 98066 291174
rect 98302 290938 98334 291174
rect 97714 290854 98334 290938
rect 97714 290618 97746 290854
rect 97982 290618 98066 290854
rect 98302 290618 98334 290854
rect 97714 254174 98334 290618
rect 97714 253938 97746 254174
rect 97982 253938 98066 254174
rect 98302 253938 98334 254174
rect 97714 253854 98334 253938
rect 97714 253618 97746 253854
rect 97982 253618 98066 253854
rect 98302 253618 98334 253854
rect 97714 217174 98334 253618
rect 97714 216938 97746 217174
rect 97982 216938 98066 217174
rect 98302 216938 98334 217174
rect 97714 216854 98334 216938
rect 97714 216618 97746 216854
rect 97982 216618 98066 216854
rect 98302 216618 98334 216854
rect 97714 180174 98334 216618
rect 97714 179938 97746 180174
rect 97982 179938 98066 180174
rect 98302 179938 98334 180174
rect 97714 179854 98334 179938
rect 97714 179618 97746 179854
rect 97982 179618 98066 179854
rect 98302 179618 98334 179854
rect 97714 143174 98334 179618
rect 97714 142938 97746 143174
rect 97982 142938 98066 143174
rect 98302 142938 98334 143174
rect 97714 142854 98334 142938
rect 97714 142618 97746 142854
rect 97982 142618 98066 142854
rect 98302 142618 98334 142854
rect 97714 106174 98334 142618
rect 97714 105938 97746 106174
rect 97982 105938 98066 106174
rect 98302 105938 98334 106174
rect 97714 105854 98334 105938
rect 97714 105618 97746 105854
rect 97982 105618 98066 105854
rect 98302 105618 98334 105854
rect 97714 69174 98334 105618
rect 97714 68938 97746 69174
rect 97982 68938 98066 69174
rect 98302 68938 98334 69174
rect 97714 68854 98334 68938
rect 97714 68618 97746 68854
rect 97982 68618 98066 68854
rect 98302 68618 98334 68854
rect 69714 31938 69746 32174
rect 69982 31938 70066 32174
rect 70302 31938 70334 32174
rect 69714 31854 70334 31938
rect 69714 31618 69746 31854
rect 69982 31618 70066 31854
rect 70302 31618 70334 31854
rect 69714 -346 70334 31618
rect 91818 32174 92138 32206
rect 91818 31938 91860 32174
rect 92096 31938 92138 32174
rect 91818 31854 92138 31938
rect 91818 31618 91860 31854
rect 92096 31618 92138 31854
rect 91818 31586 92138 31618
rect 92766 32174 93086 32206
rect 92766 31938 92808 32174
rect 93044 31938 93086 32174
rect 92766 31854 93086 31938
rect 92766 31618 92808 31854
rect 93044 31618 93086 31854
rect 92766 31586 93086 31618
rect 93714 32174 94034 32206
rect 93714 31938 93756 32174
rect 93992 31938 94034 32174
rect 93714 31854 94034 31938
rect 93714 31618 93756 31854
rect 93992 31618 94034 31854
rect 93714 31586 94034 31618
rect 94662 32174 94982 32206
rect 94662 31938 94704 32174
rect 94940 31938 94982 32174
rect 94662 31854 94982 31938
rect 94662 31618 94704 31854
rect 94940 31618 94982 31854
rect 94662 31586 94982 31618
rect 97714 32174 98334 68618
rect 121994 705798 122614 711590
rect 121994 705562 122026 705798
rect 122262 705562 122346 705798
rect 122582 705562 122614 705798
rect 121994 705478 122614 705562
rect 121994 705242 122026 705478
rect 122262 705242 122346 705478
rect 122582 705242 122614 705478
rect 121994 694454 122614 705242
rect 121994 694218 122026 694454
rect 122262 694218 122346 694454
rect 122582 694218 122614 694454
rect 121994 694134 122614 694218
rect 121994 693898 122026 694134
rect 122262 693898 122346 694134
rect 122582 693898 122614 694134
rect 121994 657454 122614 693898
rect 121994 657218 122026 657454
rect 122262 657218 122346 657454
rect 122582 657218 122614 657454
rect 121994 657134 122614 657218
rect 121994 656898 122026 657134
rect 122262 656898 122346 657134
rect 122582 656898 122614 657134
rect 121994 620454 122614 656898
rect 121994 620218 122026 620454
rect 122262 620218 122346 620454
rect 122582 620218 122614 620454
rect 121994 620134 122614 620218
rect 121994 619898 122026 620134
rect 122262 619898 122346 620134
rect 122582 619898 122614 620134
rect 121994 583454 122614 619898
rect 121994 583218 122026 583454
rect 122262 583218 122346 583454
rect 122582 583218 122614 583454
rect 121994 583134 122614 583218
rect 121994 582898 122026 583134
rect 122262 582898 122346 583134
rect 122582 582898 122614 583134
rect 121994 546454 122614 582898
rect 121994 546218 122026 546454
rect 122262 546218 122346 546454
rect 122582 546218 122614 546454
rect 121994 546134 122614 546218
rect 121994 545898 122026 546134
rect 122262 545898 122346 546134
rect 122582 545898 122614 546134
rect 121994 509454 122614 545898
rect 121994 509218 122026 509454
rect 122262 509218 122346 509454
rect 122582 509218 122614 509454
rect 121994 509134 122614 509218
rect 121994 508898 122026 509134
rect 122262 508898 122346 509134
rect 122582 508898 122614 509134
rect 121994 472454 122614 508898
rect 121994 472218 122026 472454
rect 122262 472218 122346 472454
rect 122582 472218 122614 472454
rect 121994 472134 122614 472218
rect 121994 471898 122026 472134
rect 122262 471898 122346 472134
rect 122582 471898 122614 472134
rect 121994 435454 122614 471898
rect 121994 435218 122026 435454
rect 122262 435218 122346 435454
rect 122582 435218 122614 435454
rect 121994 435134 122614 435218
rect 121994 434898 122026 435134
rect 122262 434898 122346 435134
rect 122582 434898 122614 435134
rect 121994 398454 122614 434898
rect 121994 398218 122026 398454
rect 122262 398218 122346 398454
rect 122582 398218 122614 398454
rect 121994 398134 122614 398218
rect 121994 397898 122026 398134
rect 122262 397898 122346 398134
rect 122582 397898 122614 398134
rect 121994 361454 122614 397898
rect 121994 361218 122026 361454
rect 122262 361218 122346 361454
rect 122582 361218 122614 361454
rect 121994 361134 122614 361218
rect 121994 360898 122026 361134
rect 122262 360898 122346 361134
rect 122582 360898 122614 361134
rect 121994 324454 122614 360898
rect 121994 324218 122026 324454
rect 122262 324218 122346 324454
rect 122582 324218 122614 324454
rect 121994 324134 122614 324218
rect 121994 323898 122026 324134
rect 122262 323898 122346 324134
rect 122582 323898 122614 324134
rect 121994 287454 122614 323898
rect 121994 287218 122026 287454
rect 122262 287218 122346 287454
rect 122582 287218 122614 287454
rect 121994 287134 122614 287218
rect 121994 286898 122026 287134
rect 122262 286898 122346 287134
rect 122582 286898 122614 287134
rect 121994 250454 122614 286898
rect 121994 250218 122026 250454
rect 122262 250218 122346 250454
rect 122582 250218 122614 250454
rect 121994 250134 122614 250218
rect 121994 249898 122026 250134
rect 122262 249898 122346 250134
rect 122582 249898 122614 250134
rect 121994 213454 122614 249898
rect 121994 213218 122026 213454
rect 122262 213218 122346 213454
rect 122582 213218 122614 213454
rect 121994 213134 122614 213218
rect 121994 212898 122026 213134
rect 122262 212898 122346 213134
rect 122582 212898 122614 213134
rect 121994 176454 122614 212898
rect 121994 176218 122026 176454
rect 122262 176218 122346 176454
rect 122582 176218 122614 176454
rect 121994 176134 122614 176218
rect 121994 175898 122026 176134
rect 122262 175898 122346 176134
rect 122582 175898 122614 176134
rect 121994 139454 122614 175898
rect 121994 139218 122026 139454
rect 122262 139218 122346 139454
rect 122582 139218 122614 139454
rect 121994 139134 122614 139218
rect 121994 138898 122026 139134
rect 122262 138898 122346 139134
rect 122582 138898 122614 139134
rect 121994 102454 122614 138898
rect 121994 102218 122026 102454
rect 122262 102218 122346 102454
rect 122582 102218 122614 102454
rect 121994 102134 122614 102218
rect 121994 101898 122026 102134
rect 122262 101898 122346 102134
rect 122582 101898 122614 102134
rect 121994 65454 122614 101898
rect 121994 65218 122026 65454
rect 122262 65218 122346 65454
rect 122582 65218 122614 65454
rect 121994 65134 122614 65218
rect 121994 64898 122026 65134
rect 122262 64898 122346 65134
rect 122582 64898 122614 65134
rect 97714 31938 97746 32174
rect 97982 31938 98066 32174
rect 98302 31938 98334 32174
rect 97714 31854 98334 31938
rect 97714 31618 97746 31854
rect 97982 31618 98066 31854
rect 98302 31618 98334 31854
rect 92292 28454 92612 28486
rect 92292 28218 92334 28454
rect 92570 28218 92612 28454
rect 92292 28134 92612 28218
rect 92292 27898 92334 28134
rect 92570 27898 92612 28134
rect 92292 27866 92612 27898
rect 93240 28454 93560 28486
rect 93240 28218 93282 28454
rect 93518 28218 93560 28454
rect 93240 28134 93560 28218
rect 93240 27898 93282 28134
rect 93518 27898 93560 28134
rect 93240 27866 93560 27898
rect 94188 28454 94508 28486
rect 94188 28218 94230 28454
rect 94466 28218 94508 28454
rect 94188 28134 94508 28218
rect 94188 27898 94230 28134
rect 94466 27898 94508 28134
rect 94188 27866 94508 27898
rect 69714 -582 69746 -346
rect 69982 -582 70066 -346
rect 70302 -582 70334 -346
rect 69714 -666 70334 -582
rect 69714 -902 69746 -666
rect 69982 -902 70066 -666
rect 70302 -902 70334 -666
rect 69714 -7654 70334 -902
rect 97714 -346 98334 31618
rect 102017 32174 102337 32206
rect 102017 31938 102059 32174
rect 102295 31938 102337 32174
rect 102017 31854 102337 31938
rect 102017 31618 102059 31854
rect 102295 31618 102337 31854
rect 102017 31586 102337 31618
rect 108963 32174 109283 32206
rect 108963 31938 109005 32174
rect 109241 31938 109283 32174
rect 108963 31854 109283 31938
rect 108963 31618 109005 31854
rect 109241 31618 109283 31854
rect 108963 31586 109283 31618
rect 115909 32174 116229 32206
rect 115909 31938 115951 32174
rect 116187 31938 116229 32174
rect 115909 31854 116229 31938
rect 115909 31618 115951 31854
rect 116187 31618 116229 31854
rect 115909 31586 116229 31618
rect 105490 28454 105810 28486
rect 105490 28218 105532 28454
rect 105768 28218 105810 28454
rect 105490 28134 105810 28218
rect 105490 27898 105532 28134
rect 105768 27898 105810 28134
rect 105490 27866 105810 27898
rect 112436 28454 112756 28486
rect 112436 28218 112478 28454
rect 112714 28218 112756 28454
rect 112436 28134 112756 28218
rect 112436 27898 112478 28134
rect 112714 27898 112756 28134
rect 112436 27866 112756 27898
rect 119382 28454 119702 28486
rect 119382 28218 119424 28454
rect 119660 28218 119702 28454
rect 119382 28134 119702 28218
rect 119382 27898 119424 28134
rect 119660 27898 119702 28134
rect 119382 27866 119702 27898
rect 121994 28454 122614 64898
rect 125714 704838 126334 711590
rect 125714 704602 125746 704838
rect 125982 704602 126066 704838
rect 126302 704602 126334 704838
rect 125714 704518 126334 704602
rect 125714 704282 125746 704518
rect 125982 704282 126066 704518
rect 126302 704282 126334 704518
rect 125714 698174 126334 704282
rect 125714 697938 125746 698174
rect 125982 697938 126066 698174
rect 126302 697938 126334 698174
rect 125714 697854 126334 697938
rect 125714 697618 125746 697854
rect 125982 697618 126066 697854
rect 126302 697618 126334 697854
rect 125714 661174 126334 697618
rect 125714 660938 125746 661174
rect 125982 660938 126066 661174
rect 126302 660938 126334 661174
rect 125714 660854 126334 660938
rect 125714 660618 125746 660854
rect 125982 660618 126066 660854
rect 126302 660618 126334 660854
rect 125714 624174 126334 660618
rect 125714 623938 125746 624174
rect 125982 623938 126066 624174
rect 126302 623938 126334 624174
rect 125714 623854 126334 623938
rect 125714 623618 125746 623854
rect 125982 623618 126066 623854
rect 126302 623618 126334 623854
rect 125714 587174 126334 623618
rect 125714 586938 125746 587174
rect 125982 586938 126066 587174
rect 126302 586938 126334 587174
rect 125714 586854 126334 586938
rect 125714 586618 125746 586854
rect 125982 586618 126066 586854
rect 126302 586618 126334 586854
rect 125714 550174 126334 586618
rect 125714 549938 125746 550174
rect 125982 549938 126066 550174
rect 126302 549938 126334 550174
rect 125714 549854 126334 549938
rect 125714 549618 125746 549854
rect 125982 549618 126066 549854
rect 126302 549618 126334 549854
rect 125714 513174 126334 549618
rect 125714 512938 125746 513174
rect 125982 512938 126066 513174
rect 126302 512938 126334 513174
rect 125714 512854 126334 512938
rect 125714 512618 125746 512854
rect 125982 512618 126066 512854
rect 126302 512618 126334 512854
rect 125714 476174 126334 512618
rect 125714 475938 125746 476174
rect 125982 475938 126066 476174
rect 126302 475938 126334 476174
rect 125714 475854 126334 475938
rect 125714 475618 125746 475854
rect 125982 475618 126066 475854
rect 126302 475618 126334 475854
rect 125714 439174 126334 475618
rect 125714 438938 125746 439174
rect 125982 438938 126066 439174
rect 126302 438938 126334 439174
rect 125714 438854 126334 438938
rect 125714 438618 125746 438854
rect 125982 438618 126066 438854
rect 126302 438618 126334 438854
rect 125714 402174 126334 438618
rect 125714 401938 125746 402174
rect 125982 401938 126066 402174
rect 126302 401938 126334 402174
rect 125714 401854 126334 401938
rect 125714 401618 125746 401854
rect 125982 401618 126066 401854
rect 126302 401618 126334 401854
rect 125714 365174 126334 401618
rect 125714 364938 125746 365174
rect 125982 364938 126066 365174
rect 126302 364938 126334 365174
rect 125714 364854 126334 364938
rect 125714 364618 125746 364854
rect 125982 364618 126066 364854
rect 126302 364618 126334 364854
rect 125714 328174 126334 364618
rect 125714 327938 125746 328174
rect 125982 327938 126066 328174
rect 126302 327938 126334 328174
rect 125714 327854 126334 327938
rect 125714 327618 125746 327854
rect 125982 327618 126066 327854
rect 126302 327618 126334 327854
rect 125714 291174 126334 327618
rect 125714 290938 125746 291174
rect 125982 290938 126066 291174
rect 126302 290938 126334 291174
rect 125714 290854 126334 290938
rect 125714 290618 125746 290854
rect 125982 290618 126066 290854
rect 126302 290618 126334 290854
rect 125714 254174 126334 290618
rect 125714 253938 125746 254174
rect 125982 253938 126066 254174
rect 126302 253938 126334 254174
rect 125714 253854 126334 253938
rect 125714 253618 125746 253854
rect 125982 253618 126066 253854
rect 126302 253618 126334 253854
rect 125714 217174 126334 253618
rect 125714 216938 125746 217174
rect 125982 216938 126066 217174
rect 126302 216938 126334 217174
rect 125714 216854 126334 216938
rect 125714 216618 125746 216854
rect 125982 216618 126066 216854
rect 126302 216618 126334 216854
rect 125714 180174 126334 216618
rect 125714 179938 125746 180174
rect 125982 179938 126066 180174
rect 126302 179938 126334 180174
rect 125714 179854 126334 179938
rect 125714 179618 125746 179854
rect 125982 179618 126066 179854
rect 126302 179618 126334 179854
rect 125714 143174 126334 179618
rect 125714 142938 125746 143174
rect 125982 142938 126066 143174
rect 126302 142938 126334 143174
rect 125714 142854 126334 142938
rect 125714 142618 125746 142854
rect 125982 142618 126066 142854
rect 126302 142618 126334 142854
rect 125714 106174 126334 142618
rect 125714 105938 125746 106174
rect 125982 105938 126066 106174
rect 126302 105938 126334 106174
rect 125714 105854 126334 105938
rect 125714 105618 125746 105854
rect 125982 105618 126066 105854
rect 126302 105618 126334 105854
rect 125714 69174 126334 105618
rect 125714 68938 125746 69174
rect 125982 68938 126066 69174
rect 126302 68938 126334 69174
rect 125714 68854 126334 68938
rect 125714 68618 125746 68854
rect 125982 68618 126066 68854
rect 126302 68618 126334 68854
rect 125714 53748 126334 68618
rect 149994 705798 150614 711590
rect 149994 705562 150026 705798
rect 150262 705562 150346 705798
rect 150582 705562 150614 705798
rect 149994 705478 150614 705562
rect 149994 705242 150026 705478
rect 150262 705242 150346 705478
rect 150582 705242 150614 705478
rect 149994 694454 150614 705242
rect 149994 694218 150026 694454
rect 150262 694218 150346 694454
rect 150582 694218 150614 694454
rect 149994 694134 150614 694218
rect 149994 693898 150026 694134
rect 150262 693898 150346 694134
rect 150582 693898 150614 694134
rect 149994 657454 150614 693898
rect 149994 657218 150026 657454
rect 150262 657218 150346 657454
rect 150582 657218 150614 657454
rect 149994 657134 150614 657218
rect 149994 656898 150026 657134
rect 150262 656898 150346 657134
rect 150582 656898 150614 657134
rect 149994 620454 150614 656898
rect 149994 620218 150026 620454
rect 150262 620218 150346 620454
rect 150582 620218 150614 620454
rect 149994 620134 150614 620218
rect 149994 619898 150026 620134
rect 150262 619898 150346 620134
rect 150582 619898 150614 620134
rect 149994 583454 150614 619898
rect 149994 583218 150026 583454
rect 150262 583218 150346 583454
rect 150582 583218 150614 583454
rect 149994 583134 150614 583218
rect 149994 582898 150026 583134
rect 150262 582898 150346 583134
rect 150582 582898 150614 583134
rect 149994 546454 150614 582898
rect 149994 546218 150026 546454
rect 150262 546218 150346 546454
rect 150582 546218 150614 546454
rect 149994 546134 150614 546218
rect 149994 545898 150026 546134
rect 150262 545898 150346 546134
rect 150582 545898 150614 546134
rect 149994 509454 150614 545898
rect 149994 509218 150026 509454
rect 150262 509218 150346 509454
rect 150582 509218 150614 509454
rect 149994 509134 150614 509218
rect 149994 508898 150026 509134
rect 150262 508898 150346 509134
rect 150582 508898 150614 509134
rect 149994 472454 150614 508898
rect 149994 472218 150026 472454
rect 150262 472218 150346 472454
rect 150582 472218 150614 472454
rect 149994 472134 150614 472218
rect 149994 471898 150026 472134
rect 150262 471898 150346 472134
rect 150582 471898 150614 472134
rect 149994 435454 150614 471898
rect 149994 435218 150026 435454
rect 150262 435218 150346 435454
rect 150582 435218 150614 435454
rect 149994 435134 150614 435218
rect 149994 434898 150026 435134
rect 150262 434898 150346 435134
rect 150582 434898 150614 435134
rect 149994 398454 150614 434898
rect 149994 398218 150026 398454
rect 150262 398218 150346 398454
rect 150582 398218 150614 398454
rect 149994 398134 150614 398218
rect 149994 397898 150026 398134
rect 150262 397898 150346 398134
rect 150582 397898 150614 398134
rect 149994 361454 150614 397898
rect 149994 361218 150026 361454
rect 150262 361218 150346 361454
rect 150582 361218 150614 361454
rect 149994 361134 150614 361218
rect 149994 360898 150026 361134
rect 150262 360898 150346 361134
rect 150582 360898 150614 361134
rect 149994 324454 150614 360898
rect 149994 324218 150026 324454
rect 150262 324218 150346 324454
rect 150582 324218 150614 324454
rect 149994 324134 150614 324218
rect 149994 323898 150026 324134
rect 150262 323898 150346 324134
rect 150582 323898 150614 324134
rect 149994 287454 150614 323898
rect 149994 287218 150026 287454
rect 150262 287218 150346 287454
rect 150582 287218 150614 287454
rect 149994 287134 150614 287218
rect 149994 286898 150026 287134
rect 150262 286898 150346 287134
rect 150582 286898 150614 287134
rect 149994 250454 150614 286898
rect 149994 250218 150026 250454
rect 150262 250218 150346 250454
rect 150582 250218 150614 250454
rect 149994 250134 150614 250218
rect 149994 249898 150026 250134
rect 150262 249898 150346 250134
rect 150582 249898 150614 250134
rect 149994 213454 150614 249898
rect 149994 213218 150026 213454
rect 150262 213218 150346 213454
rect 150582 213218 150614 213454
rect 149994 213134 150614 213218
rect 149994 212898 150026 213134
rect 150262 212898 150346 213134
rect 150582 212898 150614 213134
rect 149994 176454 150614 212898
rect 149994 176218 150026 176454
rect 150262 176218 150346 176454
rect 150582 176218 150614 176454
rect 149994 176134 150614 176218
rect 149994 175898 150026 176134
rect 150262 175898 150346 176134
rect 150582 175898 150614 176134
rect 149994 139454 150614 175898
rect 149994 139218 150026 139454
rect 150262 139218 150346 139454
rect 150582 139218 150614 139454
rect 149994 139134 150614 139218
rect 149994 138898 150026 139134
rect 150262 138898 150346 139134
rect 150582 138898 150614 139134
rect 149994 102454 150614 138898
rect 149994 102218 150026 102454
rect 150262 102218 150346 102454
rect 150582 102218 150614 102454
rect 149994 102134 150614 102218
rect 149994 101898 150026 102134
rect 150262 101898 150346 102134
rect 150582 101898 150614 102134
rect 149994 65454 150614 101898
rect 149994 65218 150026 65454
rect 150262 65218 150346 65454
rect 150582 65218 150614 65454
rect 149994 65134 150614 65218
rect 149994 64898 150026 65134
rect 150262 64898 150346 65134
rect 150582 64898 150614 65134
rect 122855 32174 123175 32206
rect 122855 31938 122897 32174
rect 123133 31938 123175 32174
rect 122855 31854 123175 31938
rect 122855 31618 122897 31854
rect 123133 31618 123175 31854
rect 122855 31586 123175 31618
rect 132018 32174 132338 32206
rect 132018 31938 132060 32174
rect 132296 31938 132338 32174
rect 132018 31854 132338 31938
rect 132018 31618 132060 31854
rect 132296 31618 132338 31854
rect 132018 31586 132338 31618
rect 132966 32174 133286 32206
rect 132966 31938 133008 32174
rect 133244 31938 133286 32174
rect 132966 31854 133286 31938
rect 132966 31618 133008 31854
rect 133244 31618 133286 31854
rect 132966 31586 133286 31618
rect 133914 32174 134234 32206
rect 133914 31938 133956 32174
rect 134192 31938 134234 32174
rect 133914 31854 134234 31938
rect 133914 31618 133956 31854
rect 134192 31618 134234 31854
rect 133914 31586 134234 31618
rect 134862 32174 135182 32206
rect 134862 31938 134904 32174
rect 135140 31938 135182 32174
rect 134862 31854 135182 31938
rect 134862 31618 134904 31854
rect 135140 31618 135182 31854
rect 134862 31586 135182 31618
rect 142217 32174 142537 32206
rect 142217 31938 142259 32174
rect 142495 31938 142537 32174
rect 142217 31854 142537 31938
rect 142217 31618 142259 31854
rect 142495 31618 142537 31854
rect 142217 31586 142537 31618
rect 149163 32174 149483 32206
rect 149163 31938 149205 32174
rect 149441 31938 149483 32174
rect 149163 31854 149483 31938
rect 149163 31618 149205 31854
rect 149441 31618 149483 31854
rect 149163 31586 149483 31618
rect 121994 28218 122026 28454
rect 122262 28218 122346 28454
rect 122582 28218 122614 28454
rect 121994 28134 122614 28218
rect 121994 27898 122026 28134
rect 122262 27898 122346 28134
rect 122582 27898 122614 28134
rect 97714 -582 97746 -346
rect 97982 -582 98066 -346
rect 98302 -582 98334 -346
rect 97714 -666 98334 -582
rect 97714 -902 97746 -666
rect 97982 -902 98066 -666
rect 98302 -902 98334 -666
rect 97714 -7654 98334 -902
rect 121994 -1306 122614 27898
rect 126328 28454 126648 28486
rect 126328 28218 126370 28454
rect 126606 28218 126648 28454
rect 126328 28134 126648 28218
rect 126328 27898 126370 28134
rect 126606 27898 126648 28134
rect 126328 27866 126648 27898
rect 132492 28454 132812 28486
rect 132492 28218 132534 28454
rect 132770 28218 132812 28454
rect 132492 28134 132812 28218
rect 132492 27898 132534 28134
rect 132770 27898 132812 28134
rect 132492 27866 132812 27898
rect 133440 28454 133760 28486
rect 133440 28218 133482 28454
rect 133718 28218 133760 28454
rect 133440 28134 133760 28218
rect 133440 27898 133482 28134
rect 133718 27898 133760 28134
rect 133440 27866 133760 27898
rect 134388 28454 134708 28486
rect 134388 28218 134430 28454
rect 134666 28218 134708 28454
rect 134388 28134 134708 28218
rect 134388 27898 134430 28134
rect 134666 27898 134708 28134
rect 134388 27866 134708 27898
rect 145690 28454 146010 28486
rect 145690 28218 145732 28454
rect 145968 28218 146010 28454
rect 145690 28134 146010 28218
rect 145690 27898 145732 28134
rect 145968 27898 146010 28134
rect 145690 27866 146010 27898
rect 149994 28454 150614 64898
rect 153714 704838 154334 711590
rect 153714 704602 153746 704838
rect 153982 704602 154066 704838
rect 154302 704602 154334 704838
rect 153714 704518 154334 704602
rect 153714 704282 153746 704518
rect 153982 704282 154066 704518
rect 154302 704282 154334 704518
rect 153714 698174 154334 704282
rect 153714 697938 153746 698174
rect 153982 697938 154066 698174
rect 154302 697938 154334 698174
rect 153714 697854 154334 697938
rect 153714 697618 153746 697854
rect 153982 697618 154066 697854
rect 154302 697618 154334 697854
rect 153714 661174 154334 697618
rect 153714 660938 153746 661174
rect 153982 660938 154066 661174
rect 154302 660938 154334 661174
rect 153714 660854 154334 660938
rect 153714 660618 153746 660854
rect 153982 660618 154066 660854
rect 154302 660618 154334 660854
rect 153714 624174 154334 660618
rect 153714 623938 153746 624174
rect 153982 623938 154066 624174
rect 154302 623938 154334 624174
rect 153714 623854 154334 623938
rect 153714 623618 153746 623854
rect 153982 623618 154066 623854
rect 154302 623618 154334 623854
rect 153714 587174 154334 623618
rect 153714 586938 153746 587174
rect 153982 586938 154066 587174
rect 154302 586938 154334 587174
rect 153714 586854 154334 586938
rect 153714 586618 153746 586854
rect 153982 586618 154066 586854
rect 154302 586618 154334 586854
rect 153714 550174 154334 586618
rect 153714 549938 153746 550174
rect 153982 549938 154066 550174
rect 154302 549938 154334 550174
rect 153714 549854 154334 549938
rect 153714 549618 153746 549854
rect 153982 549618 154066 549854
rect 154302 549618 154334 549854
rect 153714 513174 154334 549618
rect 153714 512938 153746 513174
rect 153982 512938 154066 513174
rect 154302 512938 154334 513174
rect 153714 512854 154334 512938
rect 153714 512618 153746 512854
rect 153982 512618 154066 512854
rect 154302 512618 154334 512854
rect 153714 476174 154334 512618
rect 153714 475938 153746 476174
rect 153982 475938 154066 476174
rect 154302 475938 154334 476174
rect 153714 475854 154334 475938
rect 153714 475618 153746 475854
rect 153982 475618 154066 475854
rect 154302 475618 154334 475854
rect 153714 439174 154334 475618
rect 153714 438938 153746 439174
rect 153982 438938 154066 439174
rect 154302 438938 154334 439174
rect 153714 438854 154334 438938
rect 153714 438618 153746 438854
rect 153982 438618 154066 438854
rect 154302 438618 154334 438854
rect 153714 402174 154334 438618
rect 153714 401938 153746 402174
rect 153982 401938 154066 402174
rect 154302 401938 154334 402174
rect 153714 401854 154334 401938
rect 153714 401618 153746 401854
rect 153982 401618 154066 401854
rect 154302 401618 154334 401854
rect 153714 365174 154334 401618
rect 153714 364938 153746 365174
rect 153982 364938 154066 365174
rect 154302 364938 154334 365174
rect 153714 364854 154334 364938
rect 153714 364618 153746 364854
rect 153982 364618 154066 364854
rect 154302 364618 154334 364854
rect 153714 328174 154334 364618
rect 153714 327938 153746 328174
rect 153982 327938 154066 328174
rect 154302 327938 154334 328174
rect 153714 327854 154334 327938
rect 153714 327618 153746 327854
rect 153982 327618 154066 327854
rect 154302 327618 154334 327854
rect 153714 291174 154334 327618
rect 153714 290938 153746 291174
rect 153982 290938 154066 291174
rect 154302 290938 154334 291174
rect 153714 290854 154334 290938
rect 153714 290618 153746 290854
rect 153982 290618 154066 290854
rect 154302 290618 154334 290854
rect 153714 254174 154334 290618
rect 153714 253938 153746 254174
rect 153982 253938 154066 254174
rect 154302 253938 154334 254174
rect 153714 253854 154334 253938
rect 153714 253618 153746 253854
rect 153982 253618 154066 253854
rect 154302 253618 154334 253854
rect 153714 217174 154334 253618
rect 153714 216938 153746 217174
rect 153982 216938 154066 217174
rect 154302 216938 154334 217174
rect 153714 216854 154334 216938
rect 153714 216618 153746 216854
rect 153982 216618 154066 216854
rect 154302 216618 154334 216854
rect 153714 180174 154334 216618
rect 153714 179938 153746 180174
rect 153982 179938 154066 180174
rect 154302 179938 154334 180174
rect 153714 179854 154334 179938
rect 153714 179618 153746 179854
rect 153982 179618 154066 179854
rect 154302 179618 154334 179854
rect 153714 143174 154334 179618
rect 153714 142938 153746 143174
rect 153982 142938 154066 143174
rect 154302 142938 154334 143174
rect 153714 142854 154334 142938
rect 153714 142618 153746 142854
rect 153982 142618 154066 142854
rect 154302 142618 154334 142854
rect 153714 106174 154334 142618
rect 153714 105938 153746 106174
rect 153982 105938 154066 106174
rect 154302 105938 154334 106174
rect 153714 105854 154334 105938
rect 153714 105618 153746 105854
rect 153982 105618 154066 105854
rect 154302 105618 154334 105854
rect 153714 69174 154334 105618
rect 153714 68938 153746 69174
rect 153982 68938 154066 69174
rect 154302 68938 154334 69174
rect 153714 68854 154334 68938
rect 153714 68618 153746 68854
rect 153982 68618 154066 68854
rect 154302 68618 154334 68854
rect 153714 32174 154334 68618
rect 177994 705798 178614 711590
rect 177994 705562 178026 705798
rect 178262 705562 178346 705798
rect 178582 705562 178614 705798
rect 177994 705478 178614 705562
rect 177994 705242 178026 705478
rect 178262 705242 178346 705478
rect 178582 705242 178614 705478
rect 177994 694454 178614 705242
rect 177994 694218 178026 694454
rect 178262 694218 178346 694454
rect 178582 694218 178614 694454
rect 177994 694134 178614 694218
rect 177994 693898 178026 694134
rect 178262 693898 178346 694134
rect 178582 693898 178614 694134
rect 177994 657454 178614 693898
rect 177994 657218 178026 657454
rect 178262 657218 178346 657454
rect 178582 657218 178614 657454
rect 177994 657134 178614 657218
rect 177994 656898 178026 657134
rect 178262 656898 178346 657134
rect 178582 656898 178614 657134
rect 177994 620454 178614 656898
rect 177994 620218 178026 620454
rect 178262 620218 178346 620454
rect 178582 620218 178614 620454
rect 177994 620134 178614 620218
rect 177994 619898 178026 620134
rect 178262 619898 178346 620134
rect 178582 619898 178614 620134
rect 177994 583454 178614 619898
rect 177994 583218 178026 583454
rect 178262 583218 178346 583454
rect 178582 583218 178614 583454
rect 177994 583134 178614 583218
rect 177994 582898 178026 583134
rect 178262 582898 178346 583134
rect 178582 582898 178614 583134
rect 177994 546454 178614 582898
rect 177994 546218 178026 546454
rect 178262 546218 178346 546454
rect 178582 546218 178614 546454
rect 177994 546134 178614 546218
rect 177994 545898 178026 546134
rect 178262 545898 178346 546134
rect 178582 545898 178614 546134
rect 177994 509454 178614 545898
rect 177994 509218 178026 509454
rect 178262 509218 178346 509454
rect 178582 509218 178614 509454
rect 177994 509134 178614 509218
rect 177994 508898 178026 509134
rect 178262 508898 178346 509134
rect 178582 508898 178614 509134
rect 177994 472454 178614 508898
rect 177994 472218 178026 472454
rect 178262 472218 178346 472454
rect 178582 472218 178614 472454
rect 177994 472134 178614 472218
rect 177994 471898 178026 472134
rect 178262 471898 178346 472134
rect 178582 471898 178614 472134
rect 177994 435454 178614 471898
rect 177994 435218 178026 435454
rect 178262 435218 178346 435454
rect 178582 435218 178614 435454
rect 177994 435134 178614 435218
rect 177994 434898 178026 435134
rect 178262 434898 178346 435134
rect 178582 434898 178614 435134
rect 177994 398454 178614 434898
rect 177994 398218 178026 398454
rect 178262 398218 178346 398454
rect 178582 398218 178614 398454
rect 177994 398134 178614 398218
rect 177994 397898 178026 398134
rect 178262 397898 178346 398134
rect 178582 397898 178614 398134
rect 177994 361454 178614 397898
rect 177994 361218 178026 361454
rect 178262 361218 178346 361454
rect 178582 361218 178614 361454
rect 177994 361134 178614 361218
rect 177994 360898 178026 361134
rect 178262 360898 178346 361134
rect 178582 360898 178614 361134
rect 177994 324454 178614 360898
rect 177994 324218 178026 324454
rect 178262 324218 178346 324454
rect 178582 324218 178614 324454
rect 177994 324134 178614 324218
rect 177994 323898 178026 324134
rect 178262 323898 178346 324134
rect 178582 323898 178614 324134
rect 177994 287454 178614 323898
rect 177994 287218 178026 287454
rect 178262 287218 178346 287454
rect 178582 287218 178614 287454
rect 177994 287134 178614 287218
rect 177994 286898 178026 287134
rect 178262 286898 178346 287134
rect 178582 286898 178614 287134
rect 177994 250454 178614 286898
rect 177994 250218 178026 250454
rect 178262 250218 178346 250454
rect 178582 250218 178614 250454
rect 177994 250134 178614 250218
rect 177994 249898 178026 250134
rect 178262 249898 178346 250134
rect 178582 249898 178614 250134
rect 177994 213454 178614 249898
rect 177994 213218 178026 213454
rect 178262 213218 178346 213454
rect 178582 213218 178614 213454
rect 177994 213134 178614 213218
rect 177994 212898 178026 213134
rect 178262 212898 178346 213134
rect 178582 212898 178614 213134
rect 177994 176454 178614 212898
rect 177994 176218 178026 176454
rect 178262 176218 178346 176454
rect 178582 176218 178614 176454
rect 177994 176134 178614 176218
rect 177994 175898 178026 176134
rect 178262 175898 178346 176134
rect 178582 175898 178614 176134
rect 177994 139454 178614 175898
rect 177994 139218 178026 139454
rect 178262 139218 178346 139454
rect 178582 139218 178614 139454
rect 177994 139134 178614 139218
rect 177994 138898 178026 139134
rect 178262 138898 178346 139134
rect 178582 138898 178614 139134
rect 177994 102454 178614 138898
rect 177994 102218 178026 102454
rect 178262 102218 178346 102454
rect 178582 102218 178614 102454
rect 177994 102134 178614 102218
rect 177994 101898 178026 102134
rect 178262 101898 178346 102134
rect 178582 101898 178614 102134
rect 177994 65454 178614 101898
rect 177994 65218 178026 65454
rect 178262 65218 178346 65454
rect 178582 65218 178614 65454
rect 177994 65134 178614 65218
rect 177994 64898 178026 65134
rect 178262 64898 178346 65134
rect 178582 64898 178614 65134
rect 153714 31938 153746 32174
rect 153982 31938 154066 32174
rect 154302 31938 154334 32174
rect 153714 31854 154334 31938
rect 153714 31618 153746 31854
rect 153982 31618 154066 31854
rect 154302 31618 154334 31854
rect 149994 28218 150026 28454
rect 150262 28218 150346 28454
rect 150582 28218 150614 28454
rect 149994 28134 150614 28218
rect 149994 27898 150026 28134
rect 150262 27898 150346 28134
rect 150582 27898 150614 28134
rect 121994 -1542 122026 -1306
rect 122262 -1542 122346 -1306
rect 122582 -1542 122614 -1306
rect 121994 -1626 122614 -1542
rect 121994 -1862 122026 -1626
rect 122262 -1862 122346 -1626
rect 122582 -1862 122614 -1626
rect 121994 -7654 122614 -1862
rect 149994 -1306 150614 27898
rect 152636 28454 152956 28486
rect 152636 28218 152678 28454
rect 152914 28218 152956 28454
rect 152636 28134 152956 28218
rect 152636 27898 152678 28134
rect 152914 27898 152956 28134
rect 152636 27866 152956 27898
rect 149994 -1542 150026 -1306
rect 150262 -1542 150346 -1306
rect 150582 -1542 150614 -1306
rect 149994 -1626 150614 -1542
rect 149994 -1862 150026 -1626
rect 150262 -1862 150346 -1626
rect 150582 -1862 150614 -1626
rect 149994 -7654 150614 -1862
rect 153714 -346 154334 31618
rect 156109 32174 156429 32206
rect 156109 31938 156151 32174
rect 156387 31938 156429 32174
rect 156109 31854 156429 31938
rect 156109 31618 156151 31854
rect 156387 31618 156429 31854
rect 156109 31586 156429 31618
rect 163055 32174 163375 32206
rect 163055 31938 163097 32174
rect 163333 31938 163375 32174
rect 163055 31854 163375 31938
rect 163055 31618 163097 31854
rect 163333 31618 163375 31854
rect 163055 31586 163375 31618
rect 172218 32174 172538 32206
rect 172218 31938 172260 32174
rect 172496 31938 172538 32174
rect 172218 31854 172538 31938
rect 172218 31618 172260 31854
rect 172496 31618 172538 31854
rect 172218 31586 172538 31618
rect 173166 32174 173486 32206
rect 173166 31938 173208 32174
rect 173444 31938 173486 32174
rect 173166 31854 173486 31938
rect 173166 31618 173208 31854
rect 173444 31618 173486 31854
rect 173166 31586 173486 31618
rect 174114 32174 174434 32206
rect 174114 31938 174156 32174
rect 174392 31938 174434 32174
rect 174114 31854 174434 31938
rect 174114 31618 174156 31854
rect 174392 31618 174434 31854
rect 174114 31586 174434 31618
rect 175062 32174 175382 32206
rect 175062 31938 175104 32174
rect 175340 31938 175382 32174
rect 175062 31854 175382 31938
rect 175062 31618 175104 31854
rect 175340 31618 175382 31854
rect 175062 31586 175382 31618
rect 159582 28454 159902 28486
rect 159582 28218 159624 28454
rect 159860 28218 159902 28454
rect 159582 28134 159902 28218
rect 159582 27898 159624 28134
rect 159860 27898 159902 28134
rect 159582 27866 159902 27898
rect 166528 28454 166848 28486
rect 166528 28218 166570 28454
rect 166806 28218 166848 28454
rect 166528 28134 166848 28218
rect 166528 27898 166570 28134
rect 166806 27898 166848 28134
rect 166528 27866 166848 27898
rect 172692 28454 173012 28486
rect 172692 28218 172734 28454
rect 172970 28218 173012 28454
rect 172692 28134 173012 28218
rect 172692 27898 172734 28134
rect 172970 27898 173012 28134
rect 172692 27866 173012 27898
rect 173640 28454 173960 28486
rect 173640 28218 173682 28454
rect 173918 28218 173960 28454
rect 173640 28134 173960 28218
rect 173640 27898 173682 28134
rect 173918 27898 173960 28134
rect 173640 27866 173960 27898
rect 174588 28454 174908 28486
rect 174588 28218 174630 28454
rect 174866 28218 174908 28454
rect 174588 28134 174908 28218
rect 174588 27898 174630 28134
rect 174866 27898 174908 28134
rect 174588 27866 174908 27898
rect 177994 28454 178614 64898
rect 177994 28218 178026 28454
rect 178262 28218 178346 28454
rect 178582 28218 178614 28454
rect 177994 28134 178614 28218
rect 177994 27898 178026 28134
rect 178262 27898 178346 28134
rect 178582 27898 178614 28134
rect 153714 -582 153746 -346
rect 153982 -582 154066 -346
rect 154302 -582 154334 -346
rect 153714 -666 154334 -582
rect 153714 -902 153746 -666
rect 153982 -902 154066 -666
rect 154302 -902 154334 -666
rect 153714 -7654 154334 -902
rect 177994 -1306 178614 27898
rect 177994 -1542 178026 -1306
rect 178262 -1542 178346 -1306
rect 178582 -1542 178614 -1306
rect 177994 -1626 178614 -1542
rect 177994 -1862 178026 -1626
rect 178262 -1862 178346 -1626
rect 178582 -1862 178614 -1626
rect 177994 -7654 178614 -1862
rect 181714 704838 182334 711590
rect 181714 704602 181746 704838
rect 181982 704602 182066 704838
rect 182302 704602 182334 704838
rect 181714 704518 182334 704602
rect 181714 704282 181746 704518
rect 181982 704282 182066 704518
rect 182302 704282 182334 704518
rect 181714 698174 182334 704282
rect 181714 697938 181746 698174
rect 181982 697938 182066 698174
rect 182302 697938 182334 698174
rect 181714 697854 182334 697938
rect 181714 697618 181746 697854
rect 181982 697618 182066 697854
rect 182302 697618 182334 697854
rect 181714 661174 182334 697618
rect 181714 660938 181746 661174
rect 181982 660938 182066 661174
rect 182302 660938 182334 661174
rect 181714 660854 182334 660938
rect 181714 660618 181746 660854
rect 181982 660618 182066 660854
rect 182302 660618 182334 660854
rect 181714 624174 182334 660618
rect 181714 623938 181746 624174
rect 181982 623938 182066 624174
rect 182302 623938 182334 624174
rect 181714 623854 182334 623938
rect 181714 623618 181746 623854
rect 181982 623618 182066 623854
rect 182302 623618 182334 623854
rect 181714 587174 182334 623618
rect 181714 586938 181746 587174
rect 181982 586938 182066 587174
rect 182302 586938 182334 587174
rect 181714 586854 182334 586938
rect 181714 586618 181746 586854
rect 181982 586618 182066 586854
rect 182302 586618 182334 586854
rect 181714 550174 182334 586618
rect 181714 549938 181746 550174
rect 181982 549938 182066 550174
rect 182302 549938 182334 550174
rect 181714 549854 182334 549938
rect 181714 549618 181746 549854
rect 181982 549618 182066 549854
rect 182302 549618 182334 549854
rect 181714 513174 182334 549618
rect 181714 512938 181746 513174
rect 181982 512938 182066 513174
rect 182302 512938 182334 513174
rect 181714 512854 182334 512938
rect 181714 512618 181746 512854
rect 181982 512618 182066 512854
rect 182302 512618 182334 512854
rect 181714 476174 182334 512618
rect 181714 475938 181746 476174
rect 181982 475938 182066 476174
rect 182302 475938 182334 476174
rect 181714 475854 182334 475938
rect 181714 475618 181746 475854
rect 181982 475618 182066 475854
rect 182302 475618 182334 475854
rect 181714 439174 182334 475618
rect 181714 438938 181746 439174
rect 181982 438938 182066 439174
rect 182302 438938 182334 439174
rect 181714 438854 182334 438938
rect 181714 438618 181746 438854
rect 181982 438618 182066 438854
rect 182302 438618 182334 438854
rect 181714 402174 182334 438618
rect 181714 401938 181746 402174
rect 181982 401938 182066 402174
rect 182302 401938 182334 402174
rect 181714 401854 182334 401938
rect 181714 401618 181746 401854
rect 181982 401618 182066 401854
rect 182302 401618 182334 401854
rect 181714 365174 182334 401618
rect 181714 364938 181746 365174
rect 181982 364938 182066 365174
rect 182302 364938 182334 365174
rect 181714 364854 182334 364938
rect 181714 364618 181746 364854
rect 181982 364618 182066 364854
rect 182302 364618 182334 364854
rect 181714 328174 182334 364618
rect 181714 327938 181746 328174
rect 181982 327938 182066 328174
rect 182302 327938 182334 328174
rect 181714 327854 182334 327938
rect 181714 327618 181746 327854
rect 181982 327618 182066 327854
rect 182302 327618 182334 327854
rect 181714 291174 182334 327618
rect 181714 290938 181746 291174
rect 181982 290938 182066 291174
rect 182302 290938 182334 291174
rect 181714 290854 182334 290938
rect 181714 290618 181746 290854
rect 181982 290618 182066 290854
rect 182302 290618 182334 290854
rect 181714 254174 182334 290618
rect 181714 253938 181746 254174
rect 181982 253938 182066 254174
rect 182302 253938 182334 254174
rect 181714 253854 182334 253938
rect 181714 253618 181746 253854
rect 181982 253618 182066 253854
rect 182302 253618 182334 253854
rect 181714 217174 182334 253618
rect 181714 216938 181746 217174
rect 181982 216938 182066 217174
rect 182302 216938 182334 217174
rect 181714 216854 182334 216938
rect 181714 216618 181746 216854
rect 181982 216618 182066 216854
rect 182302 216618 182334 216854
rect 181714 180174 182334 216618
rect 181714 179938 181746 180174
rect 181982 179938 182066 180174
rect 182302 179938 182334 180174
rect 181714 179854 182334 179938
rect 181714 179618 181746 179854
rect 181982 179618 182066 179854
rect 182302 179618 182334 179854
rect 181714 143174 182334 179618
rect 181714 142938 181746 143174
rect 181982 142938 182066 143174
rect 182302 142938 182334 143174
rect 181714 142854 182334 142938
rect 181714 142618 181746 142854
rect 181982 142618 182066 142854
rect 182302 142618 182334 142854
rect 181714 106174 182334 142618
rect 181714 105938 181746 106174
rect 181982 105938 182066 106174
rect 182302 105938 182334 106174
rect 181714 105854 182334 105938
rect 181714 105618 181746 105854
rect 181982 105618 182066 105854
rect 182302 105618 182334 105854
rect 181714 69174 182334 105618
rect 181714 68938 181746 69174
rect 181982 68938 182066 69174
rect 182302 68938 182334 69174
rect 181714 68854 182334 68938
rect 181714 68618 181746 68854
rect 181982 68618 182066 68854
rect 182302 68618 182334 68854
rect 181714 32174 182334 68618
rect 205994 705798 206614 711590
rect 205994 705562 206026 705798
rect 206262 705562 206346 705798
rect 206582 705562 206614 705798
rect 205994 705478 206614 705562
rect 205994 705242 206026 705478
rect 206262 705242 206346 705478
rect 206582 705242 206614 705478
rect 205994 694454 206614 705242
rect 205994 694218 206026 694454
rect 206262 694218 206346 694454
rect 206582 694218 206614 694454
rect 205994 694134 206614 694218
rect 205994 693898 206026 694134
rect 206262 693898 206346 694134
rect 206582 693898 206614 694134
rect 205994 657454 206614 693898
rect 205994 657218 206026 657454
rect 206262 657218 206346 657454
rect 206582 657218 206614 657454
rect 205994 657134 206614 657218
rect 205994 656898 206026 657134
rect 206262 656898 206346 657134
rect 206582 656898 206614 657134
rect 205994 620454 206614 656898
rect 205994 620218 206026 620454
rect 206262 620218 206346 620454
rect 206582 620218 206614 620454
rect 205994 620134 206614 620218
rect 205994 619898 206026 620134
rect 206262 619898 206346 620134
rect 206582 619898 206614 620134
rect 205994 583454 206614 619898
rect 205994 583218 206026 583454
rect 206262 583218 206346 583454
rect 206582 583218 206614 583454
rect 205994 583134 206614 583218
rect 205994 582898 206026 583134
rect 206262 582898 206346 583134
rect 206582 582898 206614 583134
rect 205994 546454 206614 582898
rect 205994 546218 206026 546454
rect 206262 546218 206346 546454
rect 206582 546218 206614 546454
rect 205994 546134 206614 546218
rect 205994 545898 206026 546134
rect 206262 545898 206346 546134
rect 206582 545898 206614 546134
rect 205994 509454 206614 545898
rect 205994 509218 206026 509454
rect 206262 509218 206346 509454
rect 206582 509218 206614 509454
rect 205994 509134 206614 509218
rect 205994 508898 206026 509134
rect 206262 508898 206346 509134
rect 206582 508898 206614 509134
rect 205994 472454 206614 508898
rect 205994 472218 206026 472454
rect 206262 472218 206346 472454
rect 206582 472218 206614 472454
rect 205994 472134 206614 472218
rect 205994 471898 206026 472134
rect 206262 471898 206346 472134
rect 206582 471898 206614 472134
rect 205994 435454 206614 471898
rect 205994 435218 206026 435454
rect 206262 435218 206346 435454
rect 206582 435218 206614 435454
rect 205994 435134 206614 435218
rect 205994 434898 206026 435134
rect 206262 434898 206346 435134
rect 206582 434898 206614 435134
rect 205994 398454 206614 434898
rect 205994 398218 206026 398454
rect 206262 398218 206346 398454
rect 206582 398218 206614 398454
rect 205994 398134 206614 398218
rect 205994 397898 206026 398134
rect 206262 397898 206346 398134
rect 206582 397898 206614 398134
rect 205994 361454 206614 397898
rect 205994 361218 206026 361454
rect 206262 361218 206346 361454
rect 206582 361218 206614 361454
rect 205994 361134 206614 361218
rect 205994 360898 206026 361134
rect 206262 360898 206346 361134
rect 206582 360898 206614 361134
rect 205994 324454 206614 360898
rect 205994 324218 206026 324454
rect 206262 324218 206346 324454
rect 206582 324218 206614 324454
rect 205994 324134 206614 324218
rect 205994 323898 206026 324134
rect 206262 323898 206346 324134
rect 206582 323898 206614 324134
rect 205994 287454 206614 323898
rect 205994 287218 206026 287454
rect 206262 287218 206346 287454
rect 206582 287218 206614 287454
rect 205994 287134 206614 287218
rect 205994 286898 206026 287134
rect 206262 286898 206346 287134
rect 206582 286898 206614 287134
rect 205994 250454 206614 286898
rect 205994 250218 206026 250454
rect 206262 250218 206346 250454
rect 206582 250218 206614 250454
rect 205994 250134 206614 250218
rect 205994 249898 206026 250134
rect 206262 249898 206346 250134
rect 206582 249898 206614 250134
rect 205994 213454 206614 249898
rect 205994 213218 206026 213454
rect 206262 213218 206346 213454
rect 206582 213218 206614 213454
rect 205994 213134 206614 213218
rect 205994 212898 206026 213134
rect 206262 212898 206346 213134
rect 206582 212898 206614 213134
rect 205994 176454 206614 212898
rect 205994 176218 206026 176454
rect 206262 176218 206346 176454
rect 206582 176218 206614 176454
rect 205994 176134 206614 176218
rect 205994 175898 206026 176134
rect 206262 175898 206346 176134
rect 206582 175898 206614 176134
rect 205994 139454 206614 175898
rect 205994 139218 206026 139454
rect 206262 139218 206346 139454
rect 206582 139218 206614 139454
rect 205994 139134 206614 139218
rect 205994 138898 206026 139134
rect 206262 138898 206346 139134
rect 206582 138898 206614 139134
rect 205994 102454 206614 138898
rect 205994 102218 206026 102454
rect 206262 102218 206346 102454
rect 206582 102218 206614 102454
rect 205994 102134 206614 102218
rect 205994 101898 206026 102134
rect 206262 101898 206346 102134
rect 206582 101898 206614 102134
rect 205994 65454 206614 101898
rect 205994 65218 206026 65454
rect 206262 65218 206346 65454
rect 206582 65218 206614 65454
rect 205994 65134 206614 65218
rect 205994 64898 206026 65134
rect 206262 64898 206346 65134
rect 206582 64898 206614 65134
rect 181714 31938 181746 32174
rect 181982 31938 182066 32174
rect 182302 31938 182334 32174
rect 181714 31854 182334 31938
rect 181714 31618 181746 31854
rect 181982 31618 182066 31854
rect 182302 31618 182334 31854
rect 181714 -346 182334 31618
rect 182417 32174 182737 32206
rect 182417 31938 182459 32174
rect 182695 31938 182737 32174
rect 182417 31854 182737 31938
rect 182417 31618 182459 31854
rect 182695 31618 182737 31854
rect 182417 31586 182737 31618
rect 189363 32174 189683 32206
rect 189363 31938 189405 32174
rect 189641 31938 189683 32174
rect 189363 31854 189683 31938
rect 189363 31618 189405 31854
rect 189641 31618 189683 31854
rect 189363 31586 189683 31618
rect 196309 32174 196629 32206
rect 196309 31938 196351 32174
rect 196587 31938 196629 32174
rect 196309 31854 196629 31938
rect 196309 31618 196351 31854
rect 196587 31618 196629 31854
rect 196309 31586 196629 31618
rect 203255 32174 203575 32206
rect 203255 31938 203297 32174
rect 203533 31938 203575 32174
rect 203255 31854 203575 31938
rect 203255 31618 203297 31854
rect 203533 31618 203575 31854
rect 203255 31586 203575 31618
rect 185890 28454 186210 28486
rect 185890 28218 185932 28454
rect 186168 28218 186210 28454
rect 185890 28134 186210 28218
rect 185890 27898 185932 28134
rect 186168 27898 186210 28134
rect 185890 27866 186210 27898
rect 192836 28454 193156 28486
rect 192836 28218 192878 28454
rect 193114 28218 193156 28454
rect 192836 28134 193156 28218
rect 192836 27898 192878 28134
rect 193114 27898 193156 28134
rect 192836 27866 193156 27898
rect 199782 28454 200102 28486
rect 199782 28218 199824 28454
rect 200060 28218 200102 28454
rect 199782 28134 200102 28218
rect 199782 27898 199824 28134
rect 200060 27898 200102 28134
rect 199782 27866 200102 27898
rect 205994 28454 206614 64898
rect 209714 704838 210334 711590
rect 209714 704602 209746 704838
rect 209982 704602 210066 704838
rect 210302 704602 210334 704838
rect 209714 704518 210334 704602
rect 209714 704282 209746 704518
rect 209982 704282 210066 704518
rect 210302 704282 210334 704518
rect 209714 698174 210334 704282
rect 209714 697938 209746 698174
rect 209982 697938 210066 698174
rect 210302 697938 210334 698174
rect 209714 697854 210334 697938
rect 209714 697618 209746 697854
rect 209982 697618 210066 697854
rect 210302 697618 210334 697854
rect 209714 661174 210334 697618
rect 209714 660938 209746 661174
rect 209982 660938 210066 661174
rect 210302 660938 210334 661174
rect 209714 660854 210334 660938
rect 209714 660618 209746 660854
rect 209982 660618 210066 660854
rect 210302 660618 210334 660854
rect 209714 624174 210334 660618
rect 209714 623938 209746 624174
rect 209982 623938 210066 624174
rect 210302 623938 210334 624174
rect 209714 623854 210334 623938
rect 209714 623618 209746 623854
rect 209982 623618 210066 623854
rect 210302 623618 210334 623854
rect 209714 587174 210334 623618
rect 209714 586938 209746 587174
rect 209982 586938 210066 587174
rect 210302 586938 210334 587174
rect 209714 586854 210334 586938
rect 209714 586618 209746 586854
rect 209982 586618 210066 586854
rect 210302 586618 210334 586854
rect 209714 550174 210334 586618
rect 209714 549938 209746 550174
rect 209982 549938 210066 550174
rect 210302 549938 210334 550174
rect 209714 549854 210334 549938
rect 209714 549618 209746 549854
rect 209982 549618 210066 549854
rect 210302 549618 210334 549854
rect 209714 513174 210334 549618
rect 209714 512938 209746 513174
rect 209982 512938 210066 513174
rect 210302 512938 210334 513174
rect 209714 512854 210334 512938
rect 209714 512618 209746 512854
rect 209982 512618 210066 512854
rect 210302 512618 210334 512854
rect 209714 476174 210334 512618
rect 209714 475938 209746 476174
rect 209982 475938 210066 476174
rect 210302 475938 210334 476174
rect 209714 475854 210334 475938
rect 209714 475618 209746 475854
rect 209982 475618 210066 475854
rect 210302 475618 210334 475854
rect 209714 439174 210334 475618
rect 209714 438938 209746 439174
rect 209982 438938 210066 439174
rect 210302 438938 210334 439174
rect 209714 438854 210334 438938
rect 209714 438618 209746 438854
rect 209982 438618 210066 438854
rect 210302 438618 210334 438854
rect 209714 402174 210334 438618
rect 209714 401938 209746 402174
rect 209982 401938 210066 402174
rect 210302 401938 210334 402174
rect 209714 401854 210334 401938
rect 209714 401618 209746 401854
rect 209982 401618 210066 401854
rect 210302 401618 210334 401854
rect 209714 365174 210334 401618
rect 209714 364938 209746 365174
rect 209982 364938 210066 365174
rect 210302 364938 210334 365174
rect 209714 364854 210334 364938
rect 209714 364618 209746 364854
rect 209982 364618 210066 364854
rect 210302 364618 210334 364854
rect 209714 328174 210334 364618
rect 209714 327938 209746 328174
rect 209982 327938 210066 328174
rect 210302 327938 210334 328174
rect 209714 327854 210334 327938
rect 209714 327618 209746 327854
rect 209982 327618 210066 327854
rect 210302 327618 210334 327854
rect 209714 291174 210334 327618
rect 209714 290938 209746 291174
rect 209982 290938 210066 291174
rect 210302 290938 210334 291174
rect 209714 290854 210334 290938
rect 209714 290618 209746 290854
rect 209982 290618 210066 290854
rect 210302 290618 210334 290854
rect 209714 254174 210334 290618
rect 209714 253938 209746 254174
rect 209982 253938 210066 254174
rect 210302 253938 210334 254174
rect 209714 253854 210334 253938
rect 209714 253618 209746 253854
rect 209982 253618 210066 253854
rect 210302 253618 210334 253854
rect 209714 217174 210334 253618
rect 209714 216938 209746 217174
rect 209982 216938 210066 217174
rect 210302 216938 210334 217174
rect 209714 216854 210334 216938
rect 209714 216618 209746 216854
rect 209982 216618 210066 216854
rect 210302 216618 210334 216854
rect 209714 180174 210334 216618
rect 209714 179938 209746 180174
rect 209982 179938 210066 180174
rect 210302 179938 210334 180174
rect 209714 179854 210334 179938
rect 209714 179618 209746 179854
rect 209982 179618 210066 179854
rect 210302 179618 210334 179854
rect 209714 143174 210334 179618
rect 209714 142938 209746 143174
rect 209982 142938 210066 143174
rect 210302 142938 210334 143174
rect 209714 142854 210334 142938
rect 209714 142618 209746 142854
rect 209982 142618 210066 142854
rect 210302 142618 210334 142854
rect 209714 106174 210334 142618
rect 209714 105938 209746 106174
rect 209982 105938 210066 106174
rect 210302 105938 210334 106174
rect 209714 105854 210334 105938
rect 209714 105618 209746 105854
rect 209982 105618 210066 105854
rect 210302 105618 210334 105854
rect 209714 69174 210334 105618
rect 209714 68938 209746 69174
rect 209982 68938 210066 69174
rect 210302 68938 210334 69174
rect 209714 68854 210334 68938
rect 209714 68618 209746 68854
rect 209982 68618 210066 68854
rect 210302 68618 210334 68854
rect 209714 32174 210334 68618
rect 233994 705798 234614 711590
rect 233994 705562 234026 705798
rect 234262 705562 234346 705798
rect 234582 705562 234614 705798
rect 233994 705478 234614 705562
rect 233994 705242 234026 705478
rect 234262 705242 234346 705478
rect 234582 705242 234614 705478
rect 233994 694454 234614 705242
rect 233994 694218 234026 694454
rect 234262 694218 234346 694454
rect 234582 694218 234614 694454
rect 233994 694134 234614 694218
rect 233994 693898 234026 694134
rect 234262 693898 234346 694134
rect 234582 693898 234614 694134
rect 233994 657454 234614 693898
rect 233994 657218 234026 657454
rect 234262 657218 234346 657454
rect 234582 657218 234614 657454
rect 233994 657134 234614 657218
rect 233994 656898 234026 657134
rect 234262 656898 234346 657134
rect 234582 656898 234614 657134
rect 233994 620454 234614 656898
rect 233994 620218 234026 620454
rect 234262 620218 234346 620454
rect 234582 620218 234614 620454
rect 233994 620134 234614 620218
rect 233994 619898 234026 620134
rect 234262 619898 234346 620134
rect 234582 619898 234614 620134
rect 233994 583454 234614 619898
rect 233994 583218 234026 583454
rect 234262 583218 234346 583454
rect 234582 583218 234614 583454
rect 233994 583134 234614 583218
rect 233994 582898 234026 583134
rect 234262 582898 234346 583134
rect 234582 582898 234614 583134
rect 233994 546454 234614 582898
rect 233994 546218 234026 546454
rect 234262 546218 234346 546454
rect 234582 546218 234614 546454
rect 233994 546134 234614 546218
rect 233994 545898 234026 546134
rect 234262 545898 234346 546134
rect 234582 545898 234614 546134
rect 233994 509454 234614 545898
rect 233994 509218 234026 509454
rect 234262 509218 234346 509454
rect 234582 509218 234614 509454
rect 233994 509134 234614 509218
rect 233994 508898 234026 509134
rect 234262 508898 234346 509134
rect 234582 508898 234614 509134
rect 233994 472454 234614 508898
rect 233994 472218 234026 472454
rect 234262 472218 234346 472454
rect 234582 472218 234614 472454
rect 233994 472134 234614 472218
rect 233994 471898 234026 472134
rect 234262 471898 234346 472134
rect 234582 471898 234614 472134
rect 233994 435454 234614 471898
rect 233994 435218 234026 435454
rect 234262 435218 234346 435454
rect 234582 435218 234614 435454
rect 233994 435134 234614 435218
rect 233994 434898 234026 435134
rect 234262 434898 234346 435134
rect 234582 434898 234614 435134
rect 233994 398454 234614 434898
rect 233994 398218 234026 398454
rect 234262 398218 234346 398454
rect 234582 398218 234614 398454
rect 233994 398134 234614 398218
rect 233994 397898 234026 398134
rect 234262 397898 234346 398134
rect 234582 397898 234614 398134
rect 233994 361454 234614 397898
rect 233994 361218 234026 361454
rect 234262 361218 234346 361454
rect 234582 361218 234614 361454
rect 233994 361134 234614 361218
rect 233994 360898 234026 361134
rect 234262 360898 234346 361134
rect 234582 360898 234614 361134
rect 233994 324454 234614 360898
rect 233994 324218 234026 324454
rect 234262 324218 234346 324454
rect 234582 324218 234614 324454
rect 233994 324134 234614 324218
rect 233994 323898 234026 324134
rect 234262 323898 234346 324134
rect 234582 323898 234614 324134
rect 233994 287454 234614 323898
rect 233994 287218 234026 287454
rect 234262 287218 234346 287454
rect 234582 287218 234614 287454
rect 233994 287134 234614 287218
rect 233994 286898 234026 287134
rect 234262 286898 234346 287134
rect 234582 286898 234614 287134
rect 233994 250454 234614 286898
rect 233994 250218 234026 250454
rect 234262 250218 234346 250454
rect 234582 250218 234614 250454
rect 233994 250134 234614 250218
rect 233994 249898 234026 250134
rect 234262 249898 234346 250134
rect 234582 249898 234614 250134
rect 233994 213454 234614 249898
rect 233994 213218 234026 213454
rect 234262 213218 234346 213454
rect 234582 213218 234614 213454
rect 233994 213134 234614 213218
rect 233994 212898 234026 213134
rect 234262 212898 234346 213134
rect 234582 212898 234614 213134
rect 233994 176454 234614 212898
rect 233994 176218 234026 176454
rect 234262 176218 234346 176454
rect 234582 176218 234614 176454
rect 233994 176134 234614 176218
rect 233994 175898 234026 176134
rect 234262 175898 234346 176134
rect 234582 175898 234614 176134
rect 233994 139454 234614 175898
rect 233994 139218 234026 139454
rect 234262 139218 234346 139454
rect 234582 139218 234614 139454
rect 233994 139134 234614 139218
rect 233994 138898 234026 139134
rect 234262 138898 234346 139134
rect 234582 138898 234614 139134
rect 233994 102454 234614 138898
rect 233994 102218 234026 102454
rect 234262 102218 234346 102454
rect 234582 102218 234614 102454
rect 233994 102134 234614 102218
rect 233994 101898 234026 102134
rect 234262 101898 234346 102134
rect 234582 101898 234614 102134
rect 233994 65454 234614 101898
rect 233994 65218 234026 65454
rect 234262 65218 234346 65454
rect 234582 65218 234614 65454
rect 233994 65134 234614 65218
rect 233994 64898 234026 65134
rect 234262 64898 234346 65134
rect 234582 64898 234614 65134
rect 233994 54481 234614 64898
rect 237714 704838 238334 711590
rect 237714 704602 237746 704838
rect 237982 704602 238066 704838
rect 238302 704602 238334 704838
rect 237714 704518 238334 704602
rect 237714 704282 237746 704518
rect 237982 704282 238066 704518
rect 238302 704282 238334 704518
rect 237714 698174 238334 704282
rect 237714 697938 237746 698174
rect 237982 697938 238066 698174
rect 238302 697938 238334 698174
rect 237714 697854 238334 697938
rect 237714 697618 237746 697854
rect 237982 697618 238066 697854
rect 238302 697618 238334 697854
rect 237714 661174 238334 697618
rect 237714 660938 237746 661174
rect 237982 660938 238066 661174
rect 238302 660938 238334 661174
rect 237714 660854 238334 660938
rect 237714 660618 237746 660854
rect 237982 660618 238066 660854
rect 238302 660618 238334 660854
rect 237714 624174 238334 660618
rect 237714 623938 237746 624174
rect 237982 623938 238066 624174
rect 238302 623938 238334 624174
rect 237714 623854 238334 623938
rect 237714 623618 237746 623854
rect 237982 623618 238066 623854
rect 238302 623618 238334 623854
rect 237714 587174 238334 623618
rect 237714 586938 237746 587174
rect 237982 586938 238066 587174
rect 238302 586938 238334 587174
rect 237714 586854 238334 586938
rect 237714 586618 237746 586854
rect 237982 586618 238066 586854
rect 238302 586618 238334 586854
rect 237714 550174 238334 586618
rect 237714 549938 237746 550174
rect 237982 549938 238066 550174
rect 238302 549938 238334 550174
rect 237714 549854 238334 549938
rect 237714 549618 237746 549854
rect 237982 549618 238066 549854
rect 238302 549618 238334 549854
rect 237714 513174 238334 549618
rect 237714 512938 237746 513174
rect 237982 512938 238066 513174
rect 238302 512938 238334 513174
rect 237714 512854 238334 512938
rect 237714 512618 237746 512854
rect 237982 512618 238066 512854
rect 238302 512618 238334 512854
rect 237714 476174 238334 512618
rect 237714 475938 237746 476174
rect 237982 475938 238066 476174
rect 238302 475938 238334 476174
rect 237714 475854 238334 475938
rect 237714 475618 237746 475854
rect 237982 475618 238066 475854
rect 238302 475618 238334 475854
rect 237714 439174 238334 475618
rect 237714 438938 237746 439174
rect 237982 438938 238066 439174
rect 238302 438938 238334 439174
rect 237714 438854 238334 438938
rect 237714 438618 237746 438854
rect 237982 438618 238066 438854
rect 238302 438618 238334 438854
rect 237714 402174 238334 438618
rect 237714 401938 237746 402174
rect 237982 401938 238066 402174
rect 238302 401938 238334 402174
rect 237714 401854 238334 401938
rect 237714 401618 237746 401854
rect 237982 401618 238066 401854
rect 238302 401618 238334 401854
rect 237714 365174 238334 401618
rect 237714 364938 237746 365174
rect 237982 364938 238066 365174
rect 238302 364938 238334 365174
rect 237714 364854 238334 364938
rect 237714 364618 237746 364854
rect 237982 364618 238066 364854
rect 238302 364618 238334 364854
rect 237714 328174 238334 364618
rect 237714 327938 237746 328174
rect 237982 327938 238066 328174
rect 238302 327938 238334 328174
rect 237714 327854 238334 327938
rect 237714 327618 237746 327854
rect 237982 327618 238066 327854
rect 238302 327618 238334 327854
rect 237714 291174 238334 327618
rect 237714 290938 237746 291174
rect 237982 290938 238066 291174
rect 238302 290938 238334 291174
rect 237714 290854 238334 290938
rect 237714 290618 237746 290854
rect 237982 290618 238066 290854
rect 238302 290618 238334 290854
rect 237714 254174 238334 290618
rect 237714 253938 237746 254174
rect 237982 253938 238066 254174
rect 238302 253938 238334 254174
rect 237714 253854 238334 253938
rect 237714 253618 237746 253854
rect 237982 253618 238066 253854
rect 238302 253618 238334 253854
rect 237714 217174 238334 253618
rect 237714 216938 237746 217174
rect 237982 216938 238066 217174
rect 238302 216938 238334 217174
rect 237714 216854 238334 216938
rect 237714 216618 237746 216854
rect 237982 216618 238066 216854
rect 238302 216618 238334 216854
rect 237714 180174 238334 216618
rect 237714 179938 237746 180174
rect 237982 179938 238066 180174
rect 238302 179938 238334 180174
rect 237714 179854 238334 179938
rect 237714 179618 237746 179854
rect 237982 179618 238066 179854
rect 238302 179618 238334 179854
rect 237714 143174 238334 179618
rect 237714 142938 237746 143174
rect 237982 142938 238066 143174
rect 238302 142938 238334 143174
rect 237714 142854 238334 142938
rect 237714 142618 237746 142854
rect 237982 142618 238066 142854
rect 238302 142618 238334 142854
rect 237714 106174 238334 142618
rect 237714 105938 237746 106174
rect 237982 105938 238066 106174
rect 238302 105938 238334 106174
rect 237714 105854 238334 105938
rect 237714 105618 237746 105854
rect 237982 105618 238066 105854
rect 238302 105618 238334 105854
rect 237714 69174 238334 105618
rect 237714 68938 237746 69174
rect 237982 68938 238066 69174
rect 238302 68938 238334 69174
rect 237714 68854 238334 68938
rect 237714 68618 237746 68854
rect 237982 68618 238066 68854
rect 238302 68618 238334 68854
rect 237714 54481 238334 68618
rect 261994 705798 262614 711590
rect 261994 705562 262026 705798
rect 262262 705562 262346 705798
rect 262582 705562 262614 705798
rect 261994 705478 262614 705562
rect 261994 705242 262026 705478
rect 262262 705242 262346 705478
rect 262582 705242 262614 705478
rect 261994 694454 262614 705242
rect 261994 694218 262026 694454
rect 262262 694218 262346 694454
rect 262582 694218 262614 694454
rect 261994 694134 262614 694218
rect 261994 693898 262026 694134
rect 262262 693898 262346 694134
rect 262582 693898 262614 694134
rect 261994 657454 262614 693898
rect 261994 657218 262026 657454
rect 262262 657218 262346 657454
rect 262582 657218 262614 657454
rect 261994 657134 262614 657218
rect 261994 656898 262026 657134
rect 262262 656898 262346 657134
rect 262582 656898 262614 657134
rect 261994 620454 262614 656898
rect 261994 620218 262026 620454
rect 262262 620218 262346 620454
rect 262582 620218 262614 620454
rect 261994 620134 262614 620218
rect 261994 619898 262026 620134
rect 262262 619898 262346 620134
rect 262582 619898 262614 620134
rect 261994 583454 262614 619898
rect 261994 583218 262026 583454
rect 262262 583218 262346 583454
rect 262582 583218 262614 583454
rect 261994 583134 262614 583218
rect 261994 582898 262026 583134
rect 262262 582898 262346 583134
rect 262582 582898 262614 583134
rect 261994 546454 262614 582898
rect 261994 546218 262026 546454
rect 262262 546218 262346 546454
rect 262582 546218 262614 546454
rect 261994 546134 262614 546218
rect 261994 545898 262026 546134
rect 262262 545898 262346 546134
rect 262582 545898 262614 546134
rect 261994 509454 262614 545898
rect 261994 509218 262026 509454
rect 262262 509218 262346 509454
rect 262582 509218 262614 509454
rect 261994 509134 262614 509218
rect 261994 508898 262026 509134
rect 262262 508898 262346 509134
rect 262582 508898 262614 509134
rect 261994 472454 262614 508898
rect 261994 472218 262026 472454
rect 262262 472218 262346 472454
rect 262582 472218 262614 472454
rect 261994 472134 262614 472218
rect 261994 471898 262026 472134
rect 262262 471898 262346 472134
rect 262582 471898 262614 472134
rect 261994 435454 262614 471898
rect 261994 435218 262026 435454
rect 262262 435218 262346 435454
rect 262582 435218 262614 435454
rect 261994 435134 262614 435218
rect 261994 434898 262026 435134
rect 262262 434898 262346 435134
rect 262582 434898 262614 435134
rect 261994 398454 262614 434898
rect 261994 398218 262026 398454
rect 262262 398218 262346 398454
rect 262582 398218 262614 398454
rect 261994 398134 262614 398218
rect 261994 397898 262026 398134
rect 262262 397898 262346 398134
rect 262582 397898 262614 398134
rect 261994 361454 262614 397898
rect 261994 361218 262026 361454
rect 262262 361218 262346 361454
rect 262582 361218 262614 361454
rect 261994 361134 262614 361218
rect 261994 360898 262026 361134
rect 262262 360898 262346 361134
rect 262582 360898 262614 361134
rect 261994 324454 262614 360898
rect 261994 324218 262026 324454
rect 262262 324218 262346 324454
rect 262582 324218 262614 324454
rect 261994 324134 262614 324218
rect 261994 323898 262026 324134
rect 262262 323898 262346 324134
rect 262582 323898 262614 324134
rect 261994 287454 262614 323898
rect 261994 287218 262026 287454
rect 262262 287218 262346 287454
rect 262582 287218 262614 287454
rect 261994 287134 262614 287218
rect 261994 286898 262026 287134
rect 262262 286898 262346 287134
rect 262582 286898 262614 287134
rect 261994 250454 262614 286898
rect 261994 250218 262026 250454
rect 262262 250218 262346 250454
rect 262582 250218 262614 250454
rect 261994 250134 262614 250218
rect 261994 249898 262026 250134
rect 262262 249898 262346 250134
rect 262582 249898 262614 250134
rect 261994 213454 262614 249898
rect 261994 213218 262026 213454
rect 262262 213218 262346 213454
rect 262582 213218 262614 213454
rect 261994 213134 262614 213218
rect 261994 212898 262026 213134
rect 262262 212898 262346 213134
rect 262582 212898 262614 213134
rect 261994 176454 262614 212898
rect 261994 176218 262026 176454
rect 262262 176218 262346 176454
rect 262582 176218 262614 176454
rect 261994 176134 262614 176218
rect 261994 175898 262026 176134
rect 262262 175898 262346 176134
rect 262582 175898 262614 176134
rect 261994 139454 262614 175898
rect 261994 139218 262026 139454
rect 262262 139218 262346 139454
rect 262582 139218 262614 139454
rect 261994 139134 262614 139218
rect 261994 138898 262026 139134
rect 262262 138898 262346 139134
rect 262582 138898 262614 139134
rect 261994 102454 262614 138898
rect 261994 102218 262026 102454
rect 262262 102218 262346 102454
rect 262582 102218 262614 102454
rect 261994 102134 262614 102218
rect 261994 101898 262026 102134
rect 262262 101898 262346 102134
rect 262582 101898 262614 102134
rect 261994 65454 262614 101898
rect 261994 65218 262026 65454
rect 262262 65218 262346 65454
rect 262582 65218 262614 65454
rect 261994 65134 262614 65218
rect 261994 64898 262026 65134
rect 262262 64898 262346 65134
rect 262582 64898 262614 65134
rect 261994 53393 262614 64898
rect 265714 704838 266334 711590
rect 265714 704602 265746 704838
rect 265982 704602 266066 704838
rect 266302 704602 266334 704838
rect 265714 704518 266334 704602
rect 265714 704282 265746 704518
rect 265982 704282 266066 704518
rect 266302 704282 266334 704518
rect 265714 698174 266334 704282
rect 265714 697938 265746 698174
rect 265982 697938 266066 698174
rect 266302 697938 266334 698174
rect 265714 697854 266334 697938
rect 265714 697618 265746 697854
rect 265982 697618 266066 697854
rect 266302 697618 266334 697854
rect 265714 661174 266334 697618
rect 265714 660938 265746 661174
rect 265982 660938 266066 661174
rect 266302 660938 266334 661174
rect 265714 660854 266334 660938
rect 265714 660618 265746 660854
rect 265982 660618 266066 660854
rect 266302 660618 266334 660854
rect 265714 624174 266334 660618
rect 265714 623938 265746 624174
rect 265982 623938 266066 624174
rect 266302 623938 266334 624174
rect 265714 623854 266334 623938
rect 265714 623618 265746 623854
rect 265982 623618 266066 623854
rect 266302 623618 266334 623854
rect 265714 587174 266334 623618
rect 265714 586938 265746 587174
rect 265982 586938 266066 587174
rect 266302 586938 266334 587174
rect 265714 586854 266334 586938
rect 265714 586618 265746 586854
rect 265982 586618 266066 586854
rect 266302 586618 266334 586854
rect 265714 550174 266334 586618
rect 265714 549938 265746 550174
rect 265982 549938 266066 550174
rect 266302 549938 266334 550174
rect 265714 549854 266334 549938
rect 265714 549618 265746 549854
rect 265982 549618 266066 549854
rect 266302 549618 266334 549854
rect 265714 513174 266334 549618
rect 265714 512938 265746 513174
rect 265982 512938 266066 513174
rect 266302 512938 266334 513174
rect 265714 512854 266334 512938
rect 265714 512618 265746 512854
rect 265982 512618 266066 512854
rect 266302 512618 266334 512854
rect 265714 476174 266334 512618
rect 265714 475938 265746 476174
rect 265982 475938 266066 476174
rect 266302 475938 266334 476174
rect 265714 475854 266334 475938
rect 265714 475618 265746 475854
rect 265982 475618 266066 475854
rect 266302 475618 266334 475854
rect 265714 439174 266334 475618
rect 265714 438938 265746 439174
rect 265982 438938 266066 439174
rect 266302 438938 266334 439174
rect 265714 438854 266334 438938
rect 265714 438618 265746 438854
rect 265982 438618 266066 438854
rect 266302 438618 266334 438854
rect 265714 402174 266334 438618
rect 265714 401938 265746 402174
rect 265982 401938 266066 402174
rect 266302 401938 266334 402174
rect 265714 401854 266334 401938
rect 265714 401618 265746 401854
rect 265982 401618 266066 401854
rect 266302 401618 266334 401854
rect 265714 365174 266334 401618
rect 265714 364938 265746 365174
rect 265982 364938 266066 365174
rect 266302 364938 266334 365174
rect 265714 364854 266334 364938
rect 265714 364618 265746 364854
rect 265982 364618 266066 364854
rect 266302 364618 266334 364854
rect 265714 328174 266334 364618
rect 265714 327938 265746 328174
rect 265982 327938 266066 328174
rect 266302 327938 266334 328174
rect 265714 327854 266334 327938
rect 265714 327618 265746 327854
rect 265982 327618 266066 327854
rect 266302 327618 266334 327854
rect 265714 291174 266334 327618
rect 265714 290938 265746 291174
rect 265982 290938 266066 291174
rect 266302 290938 266334 291174
rect 265714 290854 266334 290938
rect 265714 290618 265746 290854
rect 265982 290618 266066 290854
rect 266302 290618 266334 290854
rect 265714 254174 266334 290618
rect 265714 253938 265746 254174
rect 265982 253938 266066 254174
rect 266302 253938 266334 254174
rect 265714 253854 266334 253938
rect 265714 253618 265746 253854
rect 265982 253618 266066 253854
rect 266302 253618 266334 253854
rect 265714 217174 266334 253618
rect 265714 216938 265746 217174
rect 265982 216938 266066 217174
rect 266302 216938 266334 217174
rect 265714 216854 266334 216938
rect 265714 216618 265746 216854
rect 265982 216618 266066 216854
rect 266302 216618 266334 216854
rect 265714 180174 266334 216618
rect 265714 179938 265746 180174
rect 265982 179938 266066 180174
rect 266302 179938 266334 180174
rect 265714 179854 266334 179938
rect 265714 179618 265746 179854
rect 265982 179618 266066 179854
rect 266302 179618 266334 179854
rect 265714 143174 266334 179618
rect 265714 142938 265746 143174
rect 265982 142938 266066 143174
rect 266302 142938 266334 143174
rect 265714 142854 266334 142938
rect 265714 142618 265746 142854
rect 265982 142618 266066 142854
rect 266302 142618 266334 142854
rect 265714 106174 266334 142618
rect 265714 105938 265746 106174
rect 265982 105938 266066 106174
rect 266302 105938 266334 106174
rect 265714 105854 266334 105938
rect 265714 105618 265746 105854
rect 265982 105618 266066 105854
rect 266302 105618 266334 105854
rect 265714 69174 266334 105618
rect 265714 68938 265746 69174
rect 265982 68938 266066 69174
rect 266302 68938 266334 69174
rect 265714 68854 266334 68938
rect 265714 68618 265746 68854
rect 265982 68618 266066 68854
rect 266302 68618 266334 68854
rect 265714 53748 266334 68618
rect 289994 705798 290614 711590
rect 289994 705562 290026 705798
rect 290262 705562 290346 705798
rect 290582 705562 290614 705798
rect 289994 705478 290614 705562
rect 289994 705242 290026 705478
rect 290262 705242 290346 705478
rect 290582 705242 290614 705478
rect 289994 694454 290614 705242
rect 289994 694218 290026 694454
rect 290262 694218 290346 694454
rect 290582 694218 290614 694454
rect 289994 694134 290614 694218
rect 289994 693898 290026 694134
rect 290262 693898 290346 694134
rect 290582 693898 290614 694134
rect 289994 657454 290614 693898
rect 289994 657218 290026 657454
rect 290262 657218 290346 657454
rect 290582 657218 290614 657454
rect 289994 657134 290614 657218
rect 289994 656898 290026 657134
rect 290262 656898 290346 657134
rect 290582 656898 290614 657134
rect 289994 620454 290614 656898
rect 289994 620218 290026 620454
rect 290262 620218 290346 620454
rect 290582 620218 290614 620454
rect 289994 620134 290614 620218
rect 289994 619898 290026 620134
rect 290262 619898 290346 620134
rect 290582 619898 290614 620134
rect 289994 583454 290614 619898
rect 289994 583218 290026 583454
rect 290262 583218 290346 583454
rect 290582 583218 290614 583454
rect 289994 583134 290614 583218
rect 289994 582898 290026 583134
rect 290262 582898 290346 583134
rect 290582 582898 290614 583134
rect 289994 546454 290614 582898
rect 289994 546218 290026 546454
rect 290262 546218 290346 546454
rect 290582 546218 290614 546454
rect 289994 546134 290614 546218
rect 289994 545898 290026 546134
rect 290262 545898 290346 546134
rect 290582 545898 290614 546134
rect 289994 509454 290614 545898
rect 289994 509218 290026 509454
rect 290262 509218 290346 509454
rect 290582 509218 290614 509454
rect 289994 509134 290614 509218
rect 289994 508898 290026 509134
rect 290262 508898 290346 509134
rect 290582 508898 290614 509134
rect 289994 472454 290614 508898
rect 289994 472218 290026 472454
rect 290262 472218 290346 472454
rect 290582 472218 290614 472454
rect 289994 472134 290614 472218
rect 289994 471898 290026 472134
rect 290262 471898 290346 472134
rect 290582 471898 290614 472134
rect 289994 435454 290614 471898
rect 289994 435218 290026 435454
rect 290262 435218 290346 435454
rect 290582 435218 290614 435454
rect 289994 435134 290614 435218
rect 289994 434898 290026 435134
rect 290262 434898 290346 435134
rect 290582 434898 290614 435134
rect 289994 398454 290614 434898
rect 289994 398218 290026 398454
rect 290262 398218 290346 398454
rect 290582 398218 290614 398454
rect 289994 398134 290614 398218
rect 289994 397898 290026 398134
rect 290262 397898 290346 398134
rect 290582 397898 290614 398134
rect 289994 361454 290614 397898
rect 289994 361218 290026 361454
rect 290262 361218 290346 361454
rect 290582 361218 290614 361454
rect 289994 361134 290614 361218
rect 289994 360898 290026 361134
rect 290262 360898 290346 361134
rect 290582 360898 290614 361134
rect 289994 324454 290614 360898
rect 289994 324218 290026 324454
rect 290262 324218 290346 324454
rect 290582 324218 290614 324454
rect 289994 324134 290614 324218
rect 289994 323898 290026 324134
rect 290262 323898 290346 324134
rect 290582 323898 290614 324134
rect 289994 287454 290614 323898
rect 289994 287218 290026 287454
rect 290262 287218 290346 287454
rect 290582 287218 290614 287454
rect 289994 287134 290614 287218
rect 289994 286898 290026 287134
rect 290262 286898 290346 287134
rect 290582 286898 290614 287134
rect 289994 250454 290614 286898
rect 289994 250218 290026 250454
rect 290262 250218 290346 250454
rect 290582 250218 290614 250454
rect 289994 250134 290614 250218
rect 289994 249898 290026 250134
rect 290262 249898 290346 250134
rect 290582 249898 290614 250134
rect 289994 213454 290614 249898
rect 289994 213218 290026 213454
rect 290262 213218 290346 213454
rect 290582 213218 290614 213454
rect 289994 213134 290614 213218
rect 289994 212898 290026 213134
rect 290262 212898 290346 213134
rect 290582 212898 290614 213134
rect 289994 176454 290614 212898
rect 289994 176218 290026 176454
rect 290262 176218 290346 176454
rect 290582 176218 290614 176454
rect 289994 176134 290614 176218
rect 289994 175898 290026 176134
rect 290262 175898 290346 176134
rect 290582 175898 290614 176134
rect 289994 139454 290614 175898
rect 289994 139218 290026 139454
rect 290262 139218 290346 139454
rect 290582 139218 290614 139454
rect 289994 139134 290614 139218
rect 289994 138898 290026 139134
rect 290262 138898 290346 139134
rect 290582 138898 290614 139134
rect 289994 102454 290614 138898
rect 289994 102218 290026 102454
rect 290262 102218 290346 102454
rect 290582 102218 290614 102454
rect 289994 102134 290614 102218
rect 289994 101898 290026 102134
rect 290262 101898 290346 102134
rect 290582 101898 290614 102134
rect 289994 65454 290614 101898
rect 289994 65218 290026 65454
rect 290262 65218 290346 65454
rect 290582 65218 290614 65454
rect 289994 65134 290614 65218
rect 289994 64898 290026 65134
rect 290262 64898 290346 65134
rect 290582 64898 290614 65134
rect 209714 31938 209746 32174
rect 209982 31938 210066 32174
rect 210302 31938 210334 32174
rect 209714 31854 210334 31938
rect 209714 31618 209746 31854
rect 209982 31618 210066 31854
rect 210302 31618 210334 31854
rect 205994 28218 206026 28454
rect 206262 28218 206346 28454
rect 206582 28218 206614 28454
rect 205994 28134 206614 28218
rect 205994 27898 206026 28134
rect 206262 27898 206346 28134
rect 206582 27898 206614 28134
rect 181714 -582 181746 -346
rect 181982 -582 182066 -346
rect 182302 -582 182334 -346
rect 181714 -666 182334 -582
rect 181714 -902 181746 -666
rect 181982 -902 182066 -666
rect 182302 -902 182334 -666
rect 181714 -7654 182334 -902
rect 205994 -1306 206614 27898
rect 206728 28454 207048 28486
rect 206728 28218 206770 28454
rect 207006 28218 207048 28454
rect 206728 28134 207048 28218
rect 206728 27898 206770 28134
rect 207006 27898 207048 28134
rect 206728 27866 207048 27898
rect 205994 -1542 206026 -1306
rect 206262 -1542 206346 -1306
rect 206582 -1542 206614 -1306
rect 205994 -1626 206614 -1542
rect 205994 -1862 206026 -1626
rect 206262 -1862 206346 -1626
rect 206582 -1862 206614 -1626
rect 205994 -7654 206614 -1862
rect 209714 -346 210334 31618
rect 212418 32174 212738 32206
rect 212418 31938 212460 32174
rect 212696 31938 212738 32174
rect 212418 31854 212738 31938
rect 212418 31618 212460 31854
rect 212696 31618 212738 31854
rect 212418 31586 212738 31618
rect 213366 32174 213686 32206
rect 213366 31938 213408 32174
rect 213644 31938 213686 32174
rect 213366 31854 213686 31938
rect 213366 31618 213408 31854
rect 213644 31618 213686 31854
rect 213366 31586 213686 31618
rect 214314 32174 214634 32206
rect 214314 31938 214356 32174
rect 214592 31938 214634 32174
rect 214314 31854 214634 31938
rect 214314 31618 214356 31854
rect 214592 31618 214634 31854
rect 214314 31586 214634 31618
rect 215262 32174 215582 32206
rect 215262 31938 215304 32174
rect 215540 31938 215582 32174
rect 215262 31854 215582 31938
rect 215262 31618 215304 31854
rect 215540 31618 215582 31854
rect 215262 31586 215582 31618
rect 222617 32174 222937 32206
rect 222617 31938 222659 32174
rect 222895 31938 222937 32174
rect 222617 31854 222937 31938
rect 222617 31618 222659 31854
rect 222895 31618 222937 31854
rect 222617 31586 222937 31618
rect 229563 32174 229883 32206
rect 229563 31938 229605 32174
rect 229841 31938 229883 32174
rect 229563 31854 229883 31938
rect 229563 31618 229605 31854
rect 229841 31618 229883 31854
rect 229563 31586 229883 31618
rect 236509 32174 236829 32206
rect 236509 31938 236551 32174
rect 236787 31938 236829 32174
rect 236509 31854 236829 31938
rect 236509 31618 236551 31854
rect 236787 31618 236829 31854
rect 236509 31586 236829 31618
rect 243455 32174 243775 32206
rect 243455 31938 243497 32174
rect 243733 31938 243775 32174
rect 243455 31854 243775 31938
rect 243455 31618 243497 31854
rect 243733 31618 243775 31854
rect 243455 31586 243775 31618
rect 252618 32174 252938 32206
rect 252618 31938 252660 32174
rect 252896 31938 252938 32174
rect 252618 31854 252938 31938
rect 252618 31618 252660 31854
rect 252896 31618 252938 31854
rect 252618 31586 252938 31618
rect 253566 32174 253886 32206
rect 253566 31938 253608 32174
rect 253844 31938 253886 32174
rect 253566 31854 253886 31938
rect 253566 31618 253608 31854
rect 253844 31618 253886 31854
rect 253566 31586 253886 31618
rect 254514 32174 254834 32206
rect 254514 31938 254556 32174
rect 254792 31938 254834 32174
rect 254514 31854 254834 31938
rect 254514 31618 254556 31854
rect 254792 31618 254834 31854
rect 254514 31586 254834 31618
rect 255462 32174 255782 32206
rect 255462 31938 255504 32174
rect 255740 31938 255782 32174
rect 255462 31854 255782 31938
rect 255462 31618 255504 31854
rect 255740 31618 255782 31854
rect 255462 31586 255782 31618
rect 262817 32174 263137 32206
rect 262817 31938 262859 32174
rect 263095 31938 263137 32174
rect 262817 31854 263137 31938
rect 262817 31618 262859 31854
rect 263095 31618 263137 31854
rect 262817 31586 263137 31618
rect 269763 32174 270083 32206
rect 269763 31938 269805 32174
rect 270041 31938 270083 32174
rect 269763 31854 270083 31938
rect 269763 31618 269805 31854
rect 270041 31618 270083 31854
rect 269763 31586 270083 31618
rect 276709 32174 277029 32206
rect 276709 31938 276751 32174
rect 276987 31938 277029 32174
rect 276709 31854 277029 31938
rect 276709 31618 276751 31854
rect 276987 31618 277029 31854
rect 276709 31586 277029 31618
rect 283655 32174 283975 32206
rect 283655 31938 283697 32174
rect 283933 31938 283975 32174
rect 283655 31854 283975 31938
rect 283655 31618 283697 31854
rect 283933 31618 283975 31854
rect 283655 31586 283975 31618
rect 212892 28454 213212 28486
rect 212892 28218 212934 28454
rect 213170 28218 213212 28454
rect 212892 28134 213212 28218
rect 212892 27898 212934 28134
rect 213170 27898 213212 28134
rect 212892 27866 213212 27898
rect 213840 28454 214160 28486
rect 213840 28218 213882 28454
rect 214118 28218 214160 28454
rect 213840 28134 214160 28218
rect 213840 27898 213882 28134
rect 214118 27898 214160 28134
rect 213840 27866 214160 27898
rect 214788 28454 215108 28486
rect 214788 28218 214830 28454
rect 215066 28218 215108 28454
rect 214788 28134 215108 28218
rect 214788 27898 214830 28134
rect 215066 27898 215108 28134
rect 214788 27866 215108 27898
rect 226090 28454 226410 28486
rect 226090 28218 226132 28454
rect 226368 28218 226410 28454
rect 226090 28134 226410 28218
rect 226090 27898 226132 28134
rect 226368 27898 226410 28134
rect 226090 27866 226410 27898
rect 233036 28454 233356 28486
rect 233036 28218 233078 28454
rect 233314 28218 233356 28454
rect 233036 28134 233356 28218
rect 233036 27898 233078 28134
rect 233314 27898 233356 28134
rect 233036 27866 233356 27898
rect 239982 28454 240302 28486
rect 239982 28218 240024 28454
rect 240260 28218 240302 28454
rect 239982 28134 240302 28218
rect 239982 27898 240024 28134
rect 240260 27898 240302 28134
rect 239982 27866 240302 27898
rect 246928 28454 247248 28486
rect 246928 28218 246970 28454
rect 247206 28218 247248 28454
rect 246928 28134 247248 28218
rect 246928 27898 246970 28134
rect 247206 27898 247248 28134
rect 246928 27866 247248 27898
rect 253092 28454 253412 28486
rect 253092 28218 253134 28454
rect 253370 28218 253412 28454
rect 253092 28134 253412 28218
rect 253092 27898 253134 28134
rect 253370 27898 253412 28134
rect 253092 27866 253412 27898
rect 254040 28454 254360 28486
rect 254040 28218 254082 28454
rect 254318 28218 254360 28454
rect 254040 28134 254360 28218
rect 254040 27898 254082 28134
rect 254318 27898 254360 28134
rect 254040 27866 254360 27898
rect 254988 28454 255308 28486
rect 254988 28218 255030 28454
rect 255266 28218 255308 28454
rect 254988 28134 255308 28218
rect 254988 27898 255030 28134
rect 255266 27898 255308 28134
rect 254988 27866 255308 27898
rect 266290 28454 266610 28486
rect 266290 28218 266332 28454
rect 266568 28218 266610 28454
rect 266290 28134 266610 28218
rect 266290 27898 266332 28134
rect 266568 27898 266610 28134
rect 266290 27866 266610 27898
rect 273236 28454 273556 28486
rect 273236 28218 273278 28454
rect 273514 28218 273556 28454
rect 273236 28134 273556 28218
rect 273236 27898 273278 28134
rect 273514 27898 273556 28134
rect 273236 27866 273556 27898
rect 280182 28454 280502 28486
rect 280182 28218 280224 28454
rect 280460 28218 280502 28454
rect 280182 28134 280502 28218
rect 280182 27898 280224 28134
rect 280460 27898 280502 28134
rect 280182 27866 280502 27898
rect 287128 28454 287448 28486
rect 287128 28218 287170 28454
rect 287406 28218 287448 28454
rect 287128 28134 287448 28218
rect 287128 27898 287170 28134
rect 287406 27898 287448 28134
rect 287128 27866 287448 27898
rect 289994 28454 290614 64898
rect 289994 28218 290026 28454
rect 290262 28218 290346 28454
rect 290582 28218 290614 28454
rect 289994 28134 290614 28218
rect 289994 27898 290026 28134
rect 290262 27898 290346 28134
rect 290582 27898 290614 28134
rect 209714 -582 209746 -346
rect 209982 -582 210066 -346
rect 210302 -582 210334 -346
rect 209714 -666 210334 -582
rect 209714 -902 209746 -666
rect 209982 -902 210066 -666
rect 210302 -902 210334 -666
rect 209714 -7654 210334 -902
rect 289994 -1306 290614 27898
rect 289994 -1542 290026 -1306
rect 290262 -1542 290346 -1306
rect 290582 -1542 290614 -1306
rect 289994 -1626 290614 -1542
rect 289994 -1862 290026 -1626
rect 290262 -1862 290346 -1626
rect 290582 -1862 290614 -1626
rect 289994 -7654 290614 -1862
rect 293714 704838 294334 711590
rect 293714 704602 293746 704838
rect 293982 704602 294066 704838
rect 294302 704602 294334 704838
rect 293714 704518 294334 704602
rect 293714 704282 293746 704518
rect 293982 704282 294066 704518
rect 294302 704282 294334 704518
rect 293714 698174 294334 704282
rect 293714 697938 293746 698174
rect 293982 697938 294066 698174
rect 294302 697938 294334 698174
rect 293714 697854 294334 697938
rect 293714 697618 293746 697854
rect 293982 697618 294066 697854
rect 294302 697618 294334 697854
rect 293714 661174 294334 697618
rect 293714 660938 293746 661174
rect 293982 660938 294066 661174
rect 294302 660938 294334 661174
rect 293714 660854 294334 660938
rect 293714 660618 293746 660854
rect 293982 660618 294066 660854
rect 294302 660618 294334 660854
rect 293714 624174 294334 660618
rect 293714 623938 293746 624174
rect 293982 623938 294066 624174
rect 294302 623938 294334 624174
rect 293714 623854 294334 623938
rect 293714 623618 293746 623854
rect 293982 623618 294066 623854
rect 294302 623618 294334 623854
rect 293714 587174 294334 623618
rect 293714 586938 293746 587174
rect 293982 586938 294066 587174
rect 294302 586938 294334 587174
rect 293714 586854 294334 586938
rect 293714 586618 293746 586854
rect 293982 586618 294066 586854
rect 294302 586618 294334 586854
rect 293714 550174 294334 586618
rect 293714 549938 293746 550174
rect 293982 549938 294066 550174
rect 294302 549938 294334 550174
rect 293714 549854 294334 549938
rect 293714 549618 293746 549854
rect 293982 549618 294066 549854
rect 294302 549618 294334 549854
rect 293714 513174 294334 549618
rect 293714 512938 293746 513174
rect 293982 512938 294066 513174
rect 294302 512938 294334 513174
rect 293714 512854 294334 512938
rect 293714 512618 293746 512854
rect 293982 512618 294066 512854
rect 294302 512618 294334 512854
rect 293714 476174 294334 512618
rect 293714 475938 293746 476174
rect 293982 475938 294066 476174
rect 294302 475938 294334 476174
rect 293714 475854 294334 475938
rect 293714 475618 293746 475854
rect 293982 475618 294066 475854
rect 294302 475618 294334 475854
rect 293714 439174 294334 475618
rect 293714 438938 293746 439174
rect 293982 438938 294066 439174
rect 294302 438938 294334 439174
rect 293714 438854 294334 438938
rect 293714 438618 293746 438854
rect 293982 438618 294066 438854
rect 294302 438618 294334 438854
rect 293714 402174 294334 438618
rect 293714 401938 293746 402174
rect 293982 401938 294066 402174
rect 294302 401938 294334 402174
rect 293714 401854 294334 401938
rect 293714 401618 293746 401854
rect 293982 401618 294066 401854
rect 294302 401618 294334 401854
rect 293714 365174 294334 401618
rect 293714 364938 293746 365174
rect 293982 364938 294066 365174
rect 294302 364938 294334 365174
rect 293714 364854 294334 364938
rect 293714 364618 293746 364854
rect 293982 364618 294066 364854
rect 294302 364618 294334 364854
rect 293714 328174 294334 364618
rect 293714 327938 293746 328174
rect 293982 327938 294066 328174
rect 294302 327938 294334 328174
rect 293714 327854 294334 327938
rect 293714 327618 293746 327854
rect 293982 327618 294066 327854
rect 294302 327618 294334 327854
rect 293714 291174 294334 327618
rect 293714 290938 293746 291174
rect 293982 290938 294066 291174
rect 294302 290938 294334 291174
rect 293714 290854 294334 290938
rect 293714 290618 293746 290854
rect 293982 290618 294066 290854
rect 294302 290618 294334 290854
rect 293714 254174 294334 290618
rect 293714 253938 293746 254174
rect 293982 253938 294066 254174
rect 294302 253938 294334 254174
rect 293714 253854 294334 253938
rect 293714 253618 293746 253854
rect 293982 253618 294066 253854
rect 294302 253618 294334 253854
rect 293714 217174 294334 253618
rect 293714 216938 293746 217174
rect 293982 216938 294066 217174
rect 294302 216938 294334 217174
rect 293714 216854 294334 216938
rect 293714 216618 293746 216854
rect 293982 216618 294066 216854
rect 294302 216618 294334 216854
rect 293714 180174 294334 216618
rect 293714 179938 293746 180174
rect 293982 179938 294066 180174
rect 294302 179938 294334 180174
rect 293714 179854 294334 179938
rect 293714 179618 293746 179854
rect 293982 179618 294066 179854
rect 294302 179618 294334 179854
rect 293714 143174 294334 179618
rect 293714 142938 293746 143174
rect 293982 142938 294066 143174
rect 294302 142938 294334 143174
rect 293714 142854 294334 142938
rect 293714 142618 293746 142854
rect 293982 142618 294066 142854
rect 294302 142618 294334 142854
rect 293714 106174 294334 142618
rect 293714 105938 293746 106174
rect 293982 105938 294066 106174
rect 294302 105938 294334 106174
rect 293714 105854 294334 105938
rect 293714 105618 293746 105854
rect 293982 105618 294066 105854
rect 294302 105618 294334 105854
rect 293714 69174 294334 105618
rect 293714 68938 293746 69174
rect 293982 68938 294066 69174
rect 294302 68938 294334 69174
rect 293714 68854 294334 68938
rect 293714 68618 293746 68854
rect 293982 68618 294066 68854
rect 294302 68618 294334 68854
rect 293714 32174 294334 68618
rect 293714 31938 293746 32174
rect 293982 31938 294066 32174
rect 294302 31938 294334 32174
rect 293714 31854 294334 31938
rect 293714 31618 293746 31854
rect 293982 31618 294066 31854
rect 294302 31618 294334 31854
rect 293714 -346 294334 31618
rect 293714 -582 293746 -346
rect 293982 -582 294066 -346
rect 294302 -582 294334 -346
rect 293714 -666 294334 -582
rect 293714 -902 293746 -666
rect 293982 -902 294066 -666
rect 294302 -902 294334 -666
rect 293714 -7654 294334 -902
rect 317994 705798 318614 711590
rect 317994 705562 318026 705798
rect 318262 705562 318346 705798
rect 318582 705562 318614 705798
rect 317994 705478 318614 705562
rect 317994 705242 318026 705478
rect 318262 705242 318346 705478
rect 318582 705242 318614 705478
rect 317994 694454 318614 705242
rect 317994 694218 318026 694454
rect 318262 694218 318346 694454
rect 318582 694218 318614 694454
rect 317994 694134 318614 694218
rect 317994 693898 318026 694134
rect 318262 693898 318346 694134
rect 318582 693898 318614 694134
rect 317994 657454 318614 693898
rect 317994 657218 318026 657454
rect 318262 657218 318346 657454
rect 318582 657218 318614 657454
rect 317994 657134 318614 657218
rect 317994 656898 318026 657134
rect 318262 656898 318346 657134
rect 318582 656898 318614 657134
rect 317994 620454 318614 656898
rect 317994 620218 318026 620454
rect 318262 620218 318346 620454
rect 318582 620218 318614 620454
rect 317994 620134 318614 620218
rect 317994 619898 318026 620134
rect 318262 619898 318346 620134
rect 318582 619898 318614 620134
rect 317994 583454 318614 619898
rect 317994 583218 318026 583454
rect 318262 583218 318346 583454
rect 318582 583218 318614 583454
rect 317994 583134 318614 583218
rect 317994 582898 318026 583134
rect 318262 582898 318346 583134
rect 318582 582898 318614 583134
rect 317994 546454 318614 582898
rect 317994 546218 318026 546454
rect 318262 546218 318346 546454
rect 318582 546218 318614 546454
rect 317994 546134 318614 546218
rect 317994 545898 318026 546134
rect 318262 545898 318346 546134
rect 318582 545898 318614 546134
rect 317994 509454 318614 545898
rect 317994 509218 318026 509454
rect 318262 509218 318346 509454
rect 318582 509218 318614 509454
rect 317994 509134 318614 509218
rect 317994 508898 318026 509134
rect 318262 508898 318346 509134
rect 318582 508898 318614 509134
rect 317994 472454 318614 508898
rect 317994 472218 318026 472454
rect 318262 472218 318346 472454
rect 318582 472218 318614 472454
rect 317994 472134 318614 472218
rect 317994 471898 318026 472134
rect 318262 471898 318346 472134
rect 318582 471898 318614 472134
rect 317994 435454 318614 471898
rect 317994 435218 318026 435454
rect 318262 435218 318346 435454
rect 318582 435218 318614 435454
rect 317994 435134 318614 435218
rect 317994 434898 318026 435134
rect 318262 434898 318346 435134
rect 318582 434898 318614 435134
rect 317994 398454 318614 434898
rect 317994 398218 318026 398454
rect 318262 398218 318346 398454
rect 318582 398218 318614 398454
rect 317994 398134 318614 398218
rect 317994 397898 318026 398134
rect 318262 397898 318346 398134
rect 318582 397898 318614 398134
rect 317994 361454 318614 397898
rect 317994 361218 318026 361454
rect 318262 361218 318346 361454
rect 318582 361218 318614 361454
rect 317994 361134 318614 361218
rect 317994 360898 318026 361134
rect 318262 360898 318346 361134
rect 318582 360898 318614 361134
rect 317994 324454 318614 360898
rect 317994 324218 318026 324454
rect 318262 324218 318346 324454
rect 318582 324218 318614 324454
rect 317994 324134 318614 324218
rect 317994 323898 318026 324134
rect 318262 323898 318346 324134
rect 318582 323898 318614 324134
rect 317994 287454 318614 323898
rect 317994 287218 318026 287454
rect 318262 287218 318346 287454
rect 318582 287218 318614 287454
rect 317994 287134 318614 287218
rect 317994 286898 318026 287134
rect 318262 286898 318346 287134
rect 318582 286898 318614 287134
rect 317994 250454 318614 286898
rect 317994 250218 318026 250454
rect 318262 250218 318346 250454
rect 318582 250218 318614 250454
rect 317994 250134 318614 250218
rect 317994 249898 318026 250134
rect 318262 249898 318346 250134
rect 318582 249898 318614 250134
rect 317994 213454 318614 249898
rect 317994 213218 318026 213454
rect 318262 213218 318346 213454
rect 318582 213218 318614 213454
rect 317994 213134 318614 213218
rect 317994 212898 318026 213134
rect 318262 212898 318346 213134
rect 318582 212898 318614 213134
rect 317994 176454 318614 212898
rect 317994 176218 318026 176454
rect 318262 176218 318346 176454
rect 318582 176218 318614 176454
rect 317994 176134 318614 176218
rect 317994 175898 318026 176134
rect 318262 175898 318346 176134
rect 318582 175898 318614 176134
rect 317994 139454 318614 175898
rect 317994 139218 318026 139454
rect 318262 139218 318346 139454
rect 318582 139218 318614 139454
rect 317994 139134 318614 139218
rect 317994 138898 318026 139134
rect 318262 138898 318346 139134
rect 318582 138898 318614 139134
rect 317994 102454 318614 138898
rect 317994 102218 318026 102454
rect 318262 102218 318346 102454
rect 318582 102218 318614 102454
rect 317994 102134 318614 102218
rect 317994 101898 318026 102134
rect 318262 101898 318346 102134
rect 318582 101898 318614 102134
rect 317994 65454 318614 101898
rect 317994 65218 318026 65454
rect 318262 65218 318346 65454
rect 318582 65218 318614 65454
rect 317994 65134 318614 65218
rect 317994 64898 318026 65134
rect 318262 64898 318346 65134
rect 318582 64898 318614 65134
rect 317994 28454 318614 64898
rect 317994 28218 318026 28454
rect 318262 28218 318346 28454
rect 318582 28218 318614 28454
rect 317994 28134 318614 28218
rect 317994 27898 318026 28134
rect 318262 27898 318346 28134
rect 318582 27898 318614 28134
rect 317994 -1306 318614 27898
rect 317994 -1542 318026 -1306
rect 318262 -1542 318346 -1306
rect 318582 -1542 318614 -1306
rect 317994 -1626 318614 -1542
rect 317994 -1862 318026 -1626
rect 318262 -1862 318346 -1626
rect 318582 -1862 318614 -1626
rect 317994 -7654 318614 -1862
rect 321714 704838 322334 711590
rect 321714 704602 321746 704838
rect 321982 704602 322066 704838
rect 322302 704602 322334 704838
rect 321714 704518 322334 704602
rect 321714 704282 321746 704518
rect 321982 704282 322066 704518
rect 322302 704282 322334 704518
rect 321714 698174 322334 704282
rect 321714 697938 321746 698174
rect 321982 697938 322066 698174
rect 322302 697938 322334 698174
rect 321714 697854 322334 697938
rect 321714 697618 321746 697854
rect 321982 697618 322066 697854
rect 322302 697618 322334 697854
rect 321714 661174 322334 697618
rect 321714 660938 321746 661174
rect 321982 660938 322066 661174
rect 322302 660938 322334 661174
rect 321714 660854 322334 660938
rect 321714 660618 321746 660854
rect 321982 660618 322066 660854
rect 322302 660618 322334 660854
rect 321714 624174 322334 660618
rect 321714 623938 321746 624174
rect 321982 623938 322066 624174
rect 322302 623938 322334 624174
rect 321714 623854 322334 623938
rect 321714 623618 321746 623854
rect 321982 623618 322066 623854
rect 322302 623618 322334 623854
rect 321714 587174 322334 623618
rect 321714 586938 321746 587174
rect 321982 586938 322066 587174
rect 322302 586938 322334 587174
rect 321714 586854 322334 586938
rect 321714 586618 321746 586854
rect 321982 586618 322066 586854
rect 322302 586618 322334 586854
rect 321714 550174 322334 586618
rect 321714 549938 321746 550174
rect 321982 549938 322066 550174
rect 322302 549938 322334 550174
rect 321714 549854 322334 549938
rect 321714 549618 321746 549854
rect 321982 549618 322066 549854
rect 322302 549618 322334 549854
rect 321714 513174 322334 549618
rect 321714 512938 321746 513174
rect 321982 512938 322066 513174
rect 322302 512938 322334 513174
rect 321714 512854 322334 512938
rect 321714 512618 321746 512854
rect 321982 512618 322066 512854
rect 322302 512618 322334 512854
rect 321714 476174 322334 512618
rect 321714 475938 321746 476174
rect 321982 475938 322066 476174
rect 322302 475938 322334 476174
rect 321714 475854 322334 475938
rect 321714 475618 321746 475854
rect 321982 475618 322066 475854
rect 322302 475618 322334 475854
rect 321714 439174 322334 475618
rect 321714 438938 321746 439174
rect 321982 438938 322066 439174
rect 322302 438938 322334 439174
rect 321714 438854 322334 438938
rect 321714 438618 321746 438854
rect 321982 438618 322066 438854
rect 322302 438618 322334 438854
rect 321714 402174 322334 438618
rect 321714 401938 321746 402174
rect 321982 401938 322066 402174
rect 322302 401938 322334 402174
rect 321714 401854 322334 401938
rect 321714 401618 321746 401854
rect 321982 401618 322066 401854
rect 322302 401618 322334 401854
rect 321714 365174 322334 401618
rect 321714 364938 321746 365174
rect 321982 364938 322066 365174
rect 322302 364938 322334 365174
rect 321714 364854 322334 364938
rect 321714 364618 321746 364854
rect 321982 364618 322066 364854
rect 322302 364618 322334 364854
rect 321714 328174 322334 364618
rect 321714 327938 321746 328174
rect 321982 327938 322066 328174
rect 322302 327938 322334 328174
rect 321714 327854 322334 327938
rect 321714 327618 321746 327854
rect 321982 327618 322066 327854
rect 322302 327618 322334 327854
rect 321714 291174 322334 327618
rect 321714 290938 321746 291174
rect 321982 290938 322066 291174
rect 322302 290938 322334 291174
rect 321714 290854 322334 290938
rect 321714 290618 321746 290854
rect 321982 290618 322066 290854
rect 322302 290618 322334 290854
rect 321714 254174 322334 290618
rect 321714 253938 321746 254174
rect 321982 253938 322066 254174
rect 322302 253938 322334 254174
rect 321714 253854 322334 253938
rect 321714 253618 321746 253854
rect 321982 253618 322066 253854
rect 322302 253618 322334 253854
rect 321714 217174 322334 253618
rect 321714 216938 321746 217174
rect 321982 216938 322066 217174
rect 322302 216938 322334 217174
rect 321714 216854 322334 216938
rect 321714 216618 321746 216854
rect 321982 216618 322066 216854
rect 322302 216618 322334 216854
rect 321714 180174 322334 216618
rect 321714 179938 321746 180174
rect 321982 179938 322066 180174
rect 322302 179938 322334 180174
rect 321714 179854 322334 179938
rect 321714 179618 321746 179854
rect 321982 179618 322066 179854
rect 322302 179618 322334 179854
rect 321714 143174 322334 179618
rect 321714 142938 321746 143174
rect 321982 142938 322066 143174
rect 322302 142938 322334 143174
rect 321714 142854 322334 142938
rect 321714 142618 321746 142854
rect 321982 142618 322066 142854
rect 322302 142618 322334 142854
rect 321714 106174 322334 142618
rect 321714 105938 321746 106174
rect 321982 105938 322066 106174
rect 322302 105938 322334 106174
rect 321714 105854 322334 105938
rect 321714 105618 321746 105854
rect 321982 105618 322066 105854
rect 322302 105618 322334 105854
rect 321714 69174 322334 105618
rect 321714 68938 321746 69174
rect 321982 68938 322066 69174
rect 322302 68938 322334 69174
rect 321714 68854 322334 68938
rect 321714 68618 321746 68854
rect 321982 68618 322066 68854
rect 322302 68618 322334 68854
rect 321714 32174 322334 68618
rect 321714 31938 321746 32174
rect 321982 31938 322066 32174
rect 322302 31938 322334 32174
rect 321714 31854 322334 31938
rect 321714 31618 321746 31854
rect 321982 31618 322066 31854
rect 322302 31618 322334 31854
rect 321714 -346 322334 31618
rect 321714 -582 321746 -346
rect 321982 -582 322066 -346
rect 322302 -582 322334 -346
rect 321714 -666 322334 -582
rect 321714 -902 321746 -666
rect 321982 -902 322066 -666
rect 322302 -902 322334 -666
rect 321714 -7654 322334 -902
rect 345994 705798 346614 711590
rect 345994 705562 346026 705798
rect 346262 705562 346346 705798
rect 346582 705562 346614 705798
rect 345994 705478 346614 705562
rect 345994 705242 346026 705478
rect 346262 705242 346346 705478
rect 346582 705242 346614 705478
rect 345994 694454 346614 705242
rect 345994 694218 346026 694454
rect 346262 694218 346346 694454
rect 346582 694218 346614 694454
rect 345994 694134 346614 694218
rect 345994 693898 346026 694134
rect 346262 693898 346346 694134
rect 346582 693898 346614 694134
rect 345994 657454 346614 693898
rect 345994 657218 346026 657454
rect 346262 657218 346346 657454
rect 346582 657218 346614 657454
rect 345994 657134 346614 657218
rect 345994 656898 346026 657134
rect 346262 656898 346346 657134
rect 346582 656898 346614 657134
rect 345994 620454 346614 656898
rect 345994 620218 346026 620454
rect 346262 620218 346346 620454
rect 346582 620218 346614 620454
rect 345994 620134 346614 620218
rect 345994 619898 346026 620134
rect 346262 619898 346346 620134
rect 346582 619898 346614 620134
rect 345994 583454 346614 619898
rect 345994 583218 346026 583454
rect 346262 583218 346346 583454
rect 346582 583218 346614 583454
rect 345994 583134 346614 583218
rect 345994 582898 346026 583134
rect 346262 582898 346346 583134
rect 346582 582898 346614 583134
rect 345994 546454 346614 582898
rect 345994 546218 346026 546454
rect 346262 546218 346346 546454
rect 346582 546218 346614 546454
rect 345994 546134 346614 546218
rect 345994 545898 346026 546134
rect 346262 545898 346346 546134
rect 346582 545898 346614 546134
rect 345994 509454 346614 545898
rect 345994 509218 346026 509454
rect 346262 509218 346346 509454
rect 346582 509218 346614 509454
rect 345994 509134 346614 509218
rect 345994 508898 346026 509134
rect 346262 508898 346346 509134
rect 346582 508898 346614 509134
rect 345994 472454 346614 508898
rect 345994 472218 346026 472454
rect 346262 472218 346346 472454
rect 346582 472218 346614 472454
rect 345994 472134 346614 472218
rect 345994 471898 346026 472134
rect 346262 471898 346346 472134
rect 346582 471898 346614 472134
rect 345994 435454 346614 471898
rect 345994 435218 346026 435454
rect 346262 435218 346346 435454
rect 346582 435218 346614 435454
rect 345994 435134 346614 435218
rect 345994 434898 346026 435134
rect 346262 434898 346346 435134
rect 346582 434898 346614 435134
rect 345994 398454 346614 434898
rect 345994 398218 346026 398454
rect 346262 398218 346346 398454
rect 346582 398218 346614 398454
rect 345994 398134 346614 398218
rect 345994 397898 346026 398134
rect 346262 397898 346346 398134
rect 346582 397898 346614 398134
rect 345994 361454 346614 397898
rect 345994 361218 346026 361454
rect 346262 361218 346346 361454
rect 346582 361218 346614 361454
rect 345994 361134 346614 361218
rect 345994 360898 346026 361134
rect 346262 360898 346346 361134
rect 346582 360898 346614 361134
rect 345994 324454 346614 360898
rect 345994 324218 346026 324454
rect 346262 324218 346346 324454
rect 346582 324218 346614 324454
rect 345994 324134 346614 324218
rect 345994 323898 346026 324134
rect 346262 323898 346346 324134
rect 346582 323898 346614 324134
rect 345994 287454 346614 323898
rect 345994 287218 346026 287454
rect 346262 287218 346346 287454
rect 346582 287218 346614 287454
rect 345994 287134 346614 287218
rect 345994 286898 346026 287134
rect 346262 286898 346346 287134
rect 346582 286898 346614 287134
rect 345994 250454 346614 286898
rect 345994 250218 346026 250454
rect 346262 250218 346346 250454
rect 346582 250218 346614 250454
rect 345994 250134 346614 250218
rect 345994 249898 346026 250134
rect 346262 249898 346346 250134
rect 346582 249898 346614 250134
rect 345994 213454 346614 249898
rect 345994 213218 346026 213454
rect 346262 213218 346346 213454
rect 346582 213218 346614 213454
rect 345994 213134 346614 213218
rect 345994 212898 346026 213134
rect 346262 212898 346346 213134
rect 346582 212898 346614 213134
rect 345994 176454 346614 212898
rect 345994 176218 346026 176454
rect 346262 176218 346346 176454
rect 346582 176218 346614 176454
rect 345994 176134 346614 176218
rect 345994 175898 346026 176134
rect 346262 175898 346346 176134
rect 346582 175898 346614 176134
rect 345994 139454 346614 175898
rect 345994 139218 346026 139454
rect 346262 139218 346346 139454
rect 346582 139218 346614 139454
rect 345994 139134 346614 139218
rect 345994 138898 346026 139134
rect 346262 138898 346346 139134
rect 346582 138898 346614 139134
rect 345994 102454 346614 138898
rect 345994 102218 346026 102454
rect 346262 102218 346346 102454
rect 346582 102218 346614 102454
rect 345994 102134 346614 102218
rect 345994 101898 346026 102134
rect 346262 101898 346346 102134
rect 346582 101898 346614 102134
rect 345994 65454 346614 101898
rect 345994 65218 346026 65454
rect 346262 65218 346346 65454
rect 346582 65218 346614 65454
rect 345994 65134 346614 65218
rect 345994 64898 346026 65134
rect 346262 64898 346346 65134
rect 346582 64898 346614 65134
rect 345994 28454 346614 64898
rect 345994 28218 346026 28454
rect 346262 28218 346346 28454
rect 346582 28218 346614 28454
rect 345994 28134 346614 28218
rect 345994 27898 346026 28134
rect 346262 27898 346346 28134
rect 346582 27898 346614 28134
rect 345994 -1306 346614 27898
rect 345994 -1542 346026 -1306
rect 346262 -1542 346346 -1306
rect 346582 -1542 346614 -1306
rect 345994 -1626 346614 -1542
rect 345994 -1862 346026 -1626
rect 346262 -1862 346346 -1626
rect 346582 -1862 346614 -1626
rect 345994 -7654 346614 -1862
rect 349714 704838 350334 711590
rect 349714 704602 349746 704838
rect 349982 704602 350066 704838
rect 350302 704602 350334 704838
rect 349714 704518 350334 704602
rect 349714 704282 349746 704518
rect 349982 704282 350066 704518
rect 350302 704282 350334 704518
rect 349714 698174 350334 704282
rect 349714 697938 349746 698174
rect 349982 697938 350066 698174
rect 350302 697938 350334 698174
rect 349714 697854 350334 697938
rect 349714 697618 349746 697854
rect 349982 697618 350066 697854
rect 350302 697618 350334 697854
rect 349714 661174 350334 697618
rect 349714 660938 349746 661174
rect 349982 660938 350066 661174
rect 350302 660938 350334 661174
rect 349714 660854 350334 660938
rect 349714 660618 349746 660854
rect 349982 660618 350066 660854
rect 350302 660618 350334 660854
rect 349714 624174 350334 660618
rect 349714 623938 349746 624174
rect 349982 623938 350066 624174
rect 350302 623938 350334 624174
rect 349714 623854 350334 623938
rect 349714 623618 349746 623854
rect 349982 623618 350066 623854
rect 350302 623618 350334 623854
rect 349714 587174 350334 623618
rect 349714 586938 349746 587174
rect 349982 586938 350066 587174
rect 350302 586938 350334 587174
rect 349714 586854 350334 586938
rect 349714 586618 349746 586854
rect 349982 586618 350066 586854
rect 350302 586618 350334 586854
rect 349714 550174 350334 586618
rect 349714 549938 349746 550174
rect 349982 549938 350066 550174
rect 350302 549938 350334 550174
rect 349714 549854 350334 549938
rect 349714 549618 349746 549854
rect 349982 549618 350066 549854
rect 350302 549618 350334 549854
rect 349714 513174 350334 549618
rect 349714 512938 349746 513174
rect 349982 512938 350066 513174
rect 350302 512938 350334 513174
rect 349714 512854 350334 512938
rect 349714 512618 349746 512854
rect 349982 512618 350066 512854
rect 350302 512618 350334 512854
rect 349714 476174 350334 512618
rect 349714 475938 349746 476174
rect 349982 475938 350066 476174
rect 350302 475938 350334 476174
rect 349714 475854 350334 475938
rect 349714 475618 349746 475854
rect 349982 475618 350066 475854
rect 350302 475618 350334 475854
rect 349714 439174 350334 475618
rect 349714 438938 349746 439174
rect 349982 438938 350066 439174
rect 350302 438938 350334 439174
rect 349714 438854 350334 438938
rect 349714 438618 349746 438854
rect 349982 438618 350066 438854
rect 350302 438618 350334 438854
rect 349714 402174 350334 438618
rect 349714 401938 349746 402174
rect 349982 401938 350066 402174
rect 350302 401938 350334 402174
rect 349714 401854 350334 401938
rect 349714 401618 349746 401854
rect 349982 401618 350066 401854
rect 350302 401618 350334 401854
rect 349714 365174 350334 401618
rect 349714 364938 349746 365174
rect 349982 364938 350066 365174
rect 350302 364938 350334 365174
rect 349714 364854 350334 364938
rect 349714 364618 349746 364854
rect 349982 364618 350066 364854
rect 350302 364618 350334 364854
rect 349714 328174 350334 364618
rect 349714 327938 349746 328174
rect 349982 327938 350066 328174
rect 350302 327938 350334 328174
rect 349714 327854 350334 327938
rect 349714 327618 349746 327854
rect 349982 327618 350066 327854
rect 350302 327618 350334 327854
rect 349714 291174 350334 327618
rect 349714 290938 349746 291174
rect 349982 290938 350066 291174
rect 350302 290938 350334 291174
rect 349714 290854 350334 290938
rect 349714 290618 349746 290854
rect 349982 290618 350066 290854
rect 350302 290618 350334 290854
rect 349714 254174 350334 290618
rect 349714 253938 349746 254174
rect 349982 253938 350066 254174
rect 350302 253938 350334 254174
rect 349714 253854 350334 253938
rect 349714 253618 349746 253854
rect 349982 253618 350066 253854
rect 350302 253618 350334 253854
rect 349714 217174 350334 253618
rect 349714 216938 349746 217174
rect 349982 216938 350066 217174
rect 350302 216938 350334 217174
rect 349714 216854 350334 216938
rect 349714 216618 349746 216854
rect 349982 216618 350066 216854
rect 350302 216618 350334 216854
rect 349714 180174 350334 216618
rect 349714 179938 349746 180174
rect 349982 179938 350066 180174
rect 350302 179938 350334 180174
rect 349714 179854 350334 179938
rect 349714 179618 349746 179854
rect 349982 179618 350066 179854
rect 350302 179618 350334 179854
rect 349714 143174 350334 179618
rect 349714 142938 349746 143174
rect 349982 142938 350066 143174
rect 350302 142938 350334 143174
rect 349714 142854 350334 142938
rect 349714 142618 349746 142854
rect 349982 142618 350066 142854
rect 350302 142618 350334 142854
rect 349714 106174 350334 142618
rect 349714 105938 349746 106174
rect 349982 105938 350066 106174
rect 350302 105938 350334 106174
rect 349714 105854 350334 105938
rect 349714 105618 349746 105854
rect 349982 105618 350066 105854
rect 350302 105618 350334 105854
rect 349714 69174 350334 105618
rect 349714 68938 349746 69174
rect 349982 68938 350066 69174
rect 350302 68938 350334 69174
rect 349714 68854 350334 68938
rect 349714 68618 349746 68854
rect 349982 68618 350066 68854
rect 350302 68618 350334 68854
rect 349714 32174 350334 68618
rect 349714 31938 349746 32174
rect 349982 31938 350066 32174
rect 350302 31938 350334 32174
rect 349714 31854 350334 31938
rect 349714 31618 349746 31854
rect 349982 31618 350066 31854
rect 350302 31618 350334 31854
rect 349714 -346 350334 31618
rect 349714 -582 349746 -346
rect 349982 -582 350066 -346
rect 350302 -582 350334 -346
rect 349714 -666 350334 -582
rect 349714 -902 349746 -666
rect 349982 -902 350066 -666
rect 350302 -902 350334 -666
rect 349714 -7654 350334 -902
rect 373994 705798 374614 711590
rect 373994 705562 374026 705798
rect 374262 705562 374346 705798
rect 374582 705562 374614 705798
rect 373994 705478 374614 705562
rect 373994 705242 374026 705478
rect 374262 705242 374346 705478
rect 374582 705242 374614 705478
rect 373994 694454 374614 705242
rect 373994 694218 374026 694454
rect 374262 694218 374346 694454
rect 374582 694218 374614 694454
rect 373994 694134 374614 694218
rect 373994 693898 374026 694134
rect 374262 693898 374346 694134
rect 374582 693898 374614 694134
rect 373994 657454 374614 693898
rect 373994 657218 374026 657454
rect 374262 657218 374346 657454
rect 374582 657218 374614 657454
rect 373994 657134 374614 657218
rect 373994 656898 374026 657134
rect 374262 656898 374346 657134
rect 374582 656898 374614 657134
rect 373994 620454 374614 656898
rect 373994 620218 374026 620454
rect 374262 620218 374346 620454
rect 374582 620218 374614 620454
rect 373994 620134 374614 620218
rect 373994 619898 374026 620134
rect 374262 619898 374346 620134
rect 374582 619898 374614 620134
rect 373994 583454 374614 619898
rect 373994 583218 374026 583454
rect 374262 583218 374346 583454
rect 374582 583218 374614 583454
rect 373994 583134 374614 583218
rect 373994 582898 374026 583134
rect 374262 582898 374346 583134
rect 374582 582898 374614 583134
rect 373994 546454 374614 582898
rect 373994 546218 374026 546454
rect 374262 546218 374346 546454
rect 374582 546218 374614 546454
rect 373994 546134 374614 546218
rect 373994 545898 374026 546134
rect 374262 545898 374346 546134
rect 374582 545898 374614 546134
rect 373994 509454 374614 545898
rect 373994 509218 374026 509454
rect 374262 509218 374346 509454
rect 374582 509218 374614 509454
rect 373994 509134 374614 509218
rect 373994 508898 374026 509134
rect 374262 508898 374346 509134
rect 374582 508898 374614 509134
rect 373994 472454 374614 508898
rect 373994 472218 374026 472454
rect 374262 472218 374346 472454
rect 374582 472218 374614 472454
rect 373994 472134 374614 472218
rect 373994 471898 374026 472134
rect 374262 471898 374346 472134
rect 374582 471898 374614 472134
rect 373994 435454 374614 471898
rect 373994 435218 374026 435454
rect 374262 435218 374346 435454
rect 374582 435218 374614 435454
rect 373994 435134 374614 435218
rect 373994 434898 374026 435134
rect 374262 434898 374346 435134
rect 374582 434898 374614 435134
rect 373994 398454 374614 434898
rect 373994 398218 374026 398454
rect 374262 398218 374346 398454
rect 374582 398218 374614 398454
rect 373994 398134 374614 398218
rect 373994 397898 374026 398134
rect 374262 397898 374346 398134
rect 374582 397898 374614 398134
rect 373994 361454 374614 397898
rect 373994 361218 374026 361454
rect 374262 361218 374346 361454
rect 374582 361218 374614 361454
rect 373994 361134 374614 361218
rect 373994 360898 374026 361134
rect 374262 360898 374346 361134
rect 374582 360898 374614 361134
rect 373994 324454 374614 360898
rect 373994 324218 374026 324454
rect 374262 324218 374346 324454
rect 374582 324218 374614 324454
rect 373994 324134 374614 324218
rect 373994 323898 374026 324134
rect 374262 323898 374346 324134
rect 374582 323898 374614 324134
rect 373994 287454 374614 323898
rect 373994 287218 374026 287454
rect 374262 287218 374346 287454
rect 374582 287218 374614 287454
rect 373994 287134 374614 287218
rect 373994 286898 374026 287134
rect 374262 286898 374346 287134
rect 374582 286898 374614 287134
rect 373994 250454 374614 286898
rect 373994 250218 374026 250454
rect 374262 250218 374346 250454
rect 374582 250218 374614 250454
rect 373994 250134 374614 250218
rect 373994 249898 374026 250134
rect 374262 249898 374346 250134
rect 374582 249898 374614 250134
rect 373994 213454 374614 249898
rect 373994 213218 374026 213454
rect 374262 213218 374346 213454
rect 374582 213218 374614 213454
rect 373994 213134 374614 213218
rect 373994 212898 374026 213134
rect 374262 212898 374346 213134
rect 374582 212898 374614 213134
rect 373994 176454 374614 212898
rect 373994 176218 374026 176454
rect 374262 176218 374346 176454
rect 374582 176218 374614 176454
rect 373994 176134 374614 176218
rect 373994 175898 374026 176134
rect 374262 175898 374346 176134
rect 374582 175898 374614 176134
rect 373994 139454 374614 175898
rect 373994 139218 374026 139454
rect 374262 139218 374346 139454
rect 374582 139218 374614 139454
rect 373994 139134 374614 139218
rect 373994 138898 374026 139134
rect 374262 138898 374346 139134
rect 374582 138898 374614 139134
rect 373994 102454 374614 138898
rect 373994 102218 374026 102454
rect 374262 102218 374346 102454
rect 374582 102218 374614 102454
rect 373994 102134 374614 102218
rect 373994 101898 374026 102134
rect 374262 101898 374346 102134
rect 374582 101898 374614 102134
rect 373994 65454 374614 101898
rect 373994 65218 374026 65454
rect 374262 65218 374346 65454
rect 374582 65218 374614 65454
rect 373994 65134 374614 65218
rect 373994 64898 374026 65134
rect 374262 64898 374346 65134
rect 374582 64898 374614 65134
rect 373994 28454 374614 64898
rect 373994 28218 374026 28454
rect 374262 28218 374346 28454
rect 374582 28218 374614 28454
rect 373994 28134 374614 28218
rect 373994 27898 374026 28134
rect 374262 27898 374346 28134
rect 374582 27898 374614 28134
rect 373994 -1306 374614 27898
rect 373994 -1542 374026 -1306
rect 374262 -1542 374346 -1306
rect 374582 -1542 374614 -1306
rect 373994 -1626 374614 -1542
rect 373994 -1862 374026 -1626
rect 374262 -1862 374346 -1626
rect 374582 -1862 374614 -1626
rect 373994 -7654 374614 -1862
rect 377714 704838 378334 711590
rect 377714 704602 377746 704838
rect 377982 704602 378066 704838
rect 378302 704602 378334 704838
rect 377714 704518 378334 704602
rect 377714 704282 377746 704518
rect 377982 704282 378066 704518
rect 378302 704282 378334 704518
rect 377714 698174 378334 704282
rect 377714 697938 377746 698174
rect 377982 697938 378066 698174
rect 378302 697938 378334 698174
rect 377714 697854 378334 697938
rect 377714 697618 377746 697854
rect 377982 697618 378066 697854
rect 378302 697618 378334 697854
rect 377714 661174 378334 697618
rect 377714 660938 377746 661174
rect 377982 660938 378066 661174
rect 378302 660938 378334 661174
rect 377714 660854 378334 660938
rect 377714 660618 377746 660854
rect 377982 660618 378066 660854
rect 378302 660618 378334 660854
rect 377714 624174 378334 660618
rect 377714 623938 377746 624174
rect 377982 623938 378066 624174
rect 378302 623938 378334 624174
rect 377714 623854 378334 623938
rect 377714 623618 377746 623854
rect 377982 623618 378066 623854
rect 378302 623618 378334 623854
rect 377714 587174 378334 623618
rect 377714 586938 377746 587174
rect 377982 586938 378066 587174
rect 378302 586938 378334 587174
rect 377714 586854 378334 586938
rect 377714 586618 377746 586854
rect 377982 586618 378066 586854
rect 378302 586618 378334 586854
rect 377714 550174 378334 586618
rect 377714 549938 377746 550174
rect 377982 549938 378066 550174
rect 378302 549938 378334 550174
rect 377714 549854 378334 549938
rect 377714 549618 377746 549854
rect 377982 549618 378066 549854
rect 378302 549618 378334 549854
rect 377714 513174 378334 549618
rect 377714 512938 377746 513174
rect 377982 512938 378066 513174
rect 378302 512938 378334 513174
rect 377714 512854 378334 512938
rect 377714 512618 377746 512854
rect 377982 512618 378066 512854
rect 378302 512618 378334 512854
rect 377714 476174 378334 512618
rect 377714 475938 377746 476174
rect 377982 475938 378066 476174
rect 378302 475938 378334 476174
rect 377714 475854 378334 475938
rect 377714 475618 377746 475854
rect 377982 475618 378066 475854
rect 378302 475618 378334 475854
rect 377714 439174 378334 475618
rect 377714 438938 377746 439174
rect 377982 438938 378066 439174
rect 378302 438938 378334 439174
rect 377714 438854 378334 438938
rect 377714 438618 377746 438854
rect 377982 438618 378066 438854
rect 378302 438618 378334 438854
rect 377714 402174 378334 438618
rect 377714 401938 377746 402174
rect 377982 401938 378066 402174
rect 378302 401938 378334 402174
rect 377714 401854 378334 401938
rect 377714 401618 377746 401854
rect 377982 401618 378066 401854
rect 378302 401618 378334 401854
rect 377714 365174 378334 401618
rect 377714 364938 377746 365174
rect 377982 364938 378066 365174
rect 378302 364938 378334 365174
rect 377714 364854 378334 364938
rect 377714 364618 377746 364854
rect 377982 364618 378066 364854
rect 378302 364618 378334 364854
rect 377714 328174 378334 364618
rect 377714 327938 377746 328174
rect 377982 327938 378066 328174
rect 378302 327938 378334 328174
rect 377714 327854 378334 327938
rect 377714 327618 377746 327854
rect 377982 327618 378066 327854
rect 378302 327618 378334 327854
rect 377714 291174 378334 327618
rect 377714 290938 377746 291174
rect 377982 290938 378066 291174
rect 378302 290938 378334 291174
rect 377714 290854 378334 290938
rect 377714 290618 377746 290854
rect 377982 290618 378066 290854
rect 378302 290618 378334 290854
rect 377714 254174 378334 290618
rect 377714 253938 377746 254174
rect 377982 253938 378066 254174
rect 378302 253938 378334 254174
rect 377714 253854 378334 253938
rect 377714 253618 377746 253854
rect 377982 253618 378066 253854
rect 378302 253618 378334 253854
rect 377714 217174 378334 253618
rect 377714 216938 377746 217174
rect 377982 216938 378066 217174
rect 378302 216938 378334 217174
rect 377714 216854 378334 216938
rect 377714 216618 377746 216854
rect 377982 216618 378066 216854
rect 378302 216618 378334 216854
rect 377714 180174 378334 216618
rect 377714 179938 377746 180174
rect 377982 179938 378066 180174
rect 378302 179938 378334 180174
rect 377714 179854 378334 179938
rect 377714 179618 377746 179854
rect 377982 179618 378066 179854
rect 378302 179618 378334 179854
rect 377714 143174 378334 179618
rect 377714 142938 377746 143174
rect 377982 142938 378066 143174
rect 378302 142938 378334 143174
rect 377714 142854 378334 142938
rect 377714 142618 377746 142854
rect 377982 142618 378066 142854
rect 378302 142618 378334 142854
rect 377714 106174 378334 142618
rect 377714 105938 377746 106174
rect 377982 105938 378066 106174
rect 378302 105938 378334 106174
rect 377714 105854 378334 105938
rect 377714 105618 377746 105854
rect 377982 105618 378066 105854
rect 378302 105618 378334 105854
rect 377714 69174 378334 105618
rect 377714 68938 377746 69174
rect 377982 68938 378066 69174
rect 378302 68938 378334 69174
rect 377714 68854 378334 68938
rect 377714 68618 377746 68854
rect 377982 68618 378066 68854
rect 378302 68618 378334 68854
rect 377714 32174 378334 68618
rect 377714 31938 377746 32174
rect 377982 31938 378066 32174
rect 378302 31938 378334 32174
rect 377714 31854 378334 31938
rect 377714 31618 377746 31854
rect 377982 31618 378066 31854
rect 378302 31618 378334 31854
rect 377714 -346 378334 31618
rect 377714 -582 377746 -346
rect 377982 -582 378066 -346
rect 378302 -582 378334 -346
rect 377714 -666 378334 -582
rect 377714 -902 377746 -666
rect 377982 -902 378066 -666
rect 378302 -902 378334 -666
rect 377714 -7654 378334 -902
rect 401994 705798 402614 711590
rect 401994 705562 402026 705798
rect 402262 705562 402346 705798
rect 402582 705562 402614 705798
rect 401994 705478 402614 705562
rect 401994 705242 402026 705478
rect 402262 705242 402346 705478
rect 402582 705242 402614 705478
rect 401994 694454 402614 705242
rect 401994 694218 402026 694454
rect 402262 694218 402346 694454
rect 402582 694218 402614 694454
rect 401994 694134 402614 694218
rect 401994 693898 402026 694134
rect 402262 693898 402346 694134
rect 402582 693898 402614 694134
rect 401994 657454 402614 693898
rect 401994 657218 402026 657454
rect 402262 657218 402346 657454
rect 402582 657218 402614 657454
rect 401994 657134 402614 657218
rect 401994 656898 402026 657134
rect 402262 656898 402346 657134
rect 402582 656898 402614 657134
rect 401994 620454 402614 656898
rect 401994 620218 402026 620454
rect 402262 620218 402346 620454
rect 402582 620218 402614 620454
rect 401994 620134 402614 620218
rect 401994 619898 402026 620134
rect 402262 619898 402346 620134
rect 402582 619898 402614 620134
rect 401994 583454 402614 619898
rect 401994 583218 402026 583454
rect 402262 583218 402346 583454
rect 402582 583218 402614 583454
rect 401994 583134 402614 583218
rect 401994 582898 402026 583134
rect 402262 582898 402346 583134
rect 402582 582898 402614 583134
rect 401994 546454 402614 582898
rect 401994 546218 402026 546454
rect 402262 546218 402346 546454
rect 402582 546218 402614 546454
rect 401994 546134 402614 546218
rect 401994 545898 402026 546134
rect 402262 545898 402346 546134
rect 402582 545898 402614 546134
rect 401994 509454 402614 545898
rect 401994 509218 402026 509454
rect 402262 509218 402346 509454
rect 402582 509218 402614 509454
rect 401994 509134 402614 509218
rect 401994 508898 402026 509134
rect 402262 508898 402346 509134
rect 402582 508898 402614 509134
rect 401994 472454 402614 508898
rect 401994 472218 402026 472454
rect 402262 472218 402346 472454
rect 402582 472218 402614 472454
rect 401994 472134 402614 472218
rect 401994 471898 402026 472134
rect 402262 471898 402346 472134
rect 402582 471898 402614 472134
rect 401994 435454 402614 471898
rect 401994 435218 402026 435454
rect 402262 435218 402346 435454
rect 402582 435218 402614 435454
rect 401994 435134 402614 435218
rect 401994 434898 402026 435134
rect 402262 434898 402346 435134
rect 402582 434898 402614 435134
rect 401994 398454 402614 434898
rect 401994 398218 402026 398454
rect 402262 398218 402346 398454
rect 402582 398218 402614 398454
rect 401994 398134 402614 398218
rect 401994 397898 402026 398134
rect 402262 397898 402346 398134
rect 402582 397898 402614 398134
rect 401994 361454 402614 397898
rect 401994 361218 402026 361454
rect 402262 361218 402346 361454
rect 402582 361218 402614 361454
rect 401994 361134 402614 361218
rect 401994 360898 402026 361134
rect 402262 360898 402346 361134
rect 402582 360898 402614 361134
rect 401994 324454 402614 360898
rect 401994 324218 402026 324454
rect 402262 324218 402346 324454
rect 402582 324218 402614 324454
rect 401994 324134 402614 324218
rect 401994 323898 402026 324134
rect 402262 323898 402346 324134
rect 402582 323898 402614 324134
rect 401994 287454 402614 323898
rect 401994 287218 402026 287454
rect 402262 287218 402346 287454
rect 402582 287218 402614 287454
rect 401994 287134 402614 287218
rect 401994 286898 402026 287134
rect 402262 286898 402346 287134
rect 402582 286898 402614 287134
rect 401994 250454 402614 286898
rect 401994 250218 402026 250454
rect 402262 250218 402346 250454
rect 402582 250218 402614 250454
rect 401994 250134 402614 250218
rect 401994 249898 402026 250134
rect 402262 249898 402346 250134
rect 402582 249898 402614 250134
rect 401994 213454 402614 249898
rect 401994 213218 402026 213454
rect 402262 213218 402346 213454
rect 402582 213218 402614 213454
rect 401994 213134 402614 213218
rect 401994 212898 402026 213134
rect 402262 212898 402346 213134
rect 402582 212898 402614 213134
rect 401994 176454 402614 212898
rect 401994 176218 402026 176454
rect 402262 176218 402346 176454
rect 402582 176218 402614 176454
rect 401994 176134 402614 176218
rect 401994 175898 402026 176134
rect 402262 175898 402346 176134
rect 402582 175898 402614 176134
rect 401994 139454 402614 175898
rect 401994 139218 402026 139454
rect 402262 139218 402346 139454
rect 402582 139218 402614 139454
rect 401994 139134 402614 139218
rect 401994 138898 402026 139134
rect 402262 138898 402346 139134
rect 402582 138898 402614 139134
rect 401994 102454 402614 138898
rect 401994 102218 402026 102454
rect 402262 102218 402346 102454
rect 402582 102218 402614 102454
rect 401994 102134 402614 102218
rect 401994 101898 402026 102134
rect 402262 101898 402346 102134
rect 402582 101898 402614 102134
rect 401994 65454 402614 101898
rect 401994 65218 402026 65454
rect 402262 65218 402346 65454
rect 402582 65218 402614 65454
rect 401994 65134 402614 65218
rect 401994 64898 402026 65134
rect 402262 64898 402346 65134
rect 402582 64898 402614 65134
rect 401994 28454 402614 64898
rect 401994 28218 402026 28454
rect 402262 28218 402346 28454
rect 402582 28218 402614 28454
rect 401994 28134 402614 28218
rect 401994 27898 402026 28134
rect 402262 27898 402346 28134
rect 402582 27898 402614 28134
rect 401994 -1306 402614 27898
rect 401994 -1542 402026 -1306
rect 402262 -1542 402346 -1306
rect 402582 -1542 402614 -1306
rect 401994 -1626 402614 -1542
rect 401994 -1862 402026 -1626
rect 402262 -1862 402346 -1626
rect 402582 -1862 402614 -1626
rect 401994 -7654 402614 -1862
rect 405714 704838 406334 711590
rect 405714 704602 405746 704838
rect 405982 704602 406066 704838
rect 406302 704602 406334 704838
rect 405714 704518 406334 704602
rect 405714 704282 405746 704518
rect 405982 704282 406066 704518
rect 406302 704282 406334 704518
rect 405714 698174 406334 704282
rect 405714 697938 405746 698174
rect 405982 697938 406066 698174
rect 406302 697938 406334 698174
rect 405714 697854 406334 697938
rect 405714 697618 405746 697854
rect 405982 697618 406066 697854
rect 406302 697618 406334 697854
rect 405714 661174 406334 697618
rect 405714 660938 405746 661174
rect 405982 660938 406066 661174
rect 406302 660938 406334 661174
rect 405714 660854 406334 660938
rect 405714 660618 405746 660854
rect 405982 660618 406066 660854
rect 406302 660618 406334 660854
rect 405714 624174 406334 660618
rect 405714 623938 405746 624174
rect 405982 623938 406066 624174
rect 406302 623938 406334 624174
rect 405714 623854 406334 623938
rect 405714 623618 405746 623854
rect 405982 623618 406066 623854
rect 406302 623618 406334 623854
rect 405714 587174 406334 623618
rect 405714 586938 405746 587174
rect 405982 586938 406066 587174
rect 406302 586938 406334 587174
rect 405714 586854 406334 586938
rect 405714 586618 405746 586854
rect 405982 586618 406066 586854
rect 406302 586618 406334 586854
rect 405714 550174 406334 586618
rect 405714 549938 405746 550174
rect 405982 549938 406066 550174
rect 406302 549938 406334 550174
rect 405714 549854 406334 549938
rect 405714 549618 405746 549854
rect 405982 549618 406066 549854
rect 406302 549618 406334 549854
rect 405714 513174 406334 549618
rect 405714 512938 405746 513174
rect 405982 512938 406066 513174
rect 406302 512938 406334 513174
rect 405714 512854 406334 512938
rect 405714 512618 405746 512854
rect 405982 512618 406066 512854
rect 406302 512618 406334 512854
rect 405714 476174 406334 512618
rect 405714 475938 405746 476174
rect 405982 475938 406066 476174
rect 406302 475938 406334 476174
rect 405714 475854 406334 475938
rect 405714 475618 405746 475854
rect 405982 475618 406066 475854
rect 406302 475618 406334 475854
rect 405714 439174 406334 475618
rect 405714 438938 405746 439174
rect 405982 438938 406066 439174
rect 406302 438938 406334 439174
rect 405714 438854 406334 438938
rect 405714 438618 405746 438854
rect 405982 438618 406066 438854
rect 406302 438618 406334 438854
rect 405714 402174 406334 438618
rect 405714 401938 405746 402174
rect 405982 401938 406066 402174
rect 406302 401938 406334 402174
rect 405714 401854 406334 401938
rect 405714 401618 405746 401854
rect 405982 401618 406066 401854
rect 406302 401618 406334 401854
rect 405714 365174 406334 401618
rect 405714 364938 405746 365174
rect 405982 364938 406066 365174
rect 406302 364938 406334 365174
rect 405714 364854 406334 364938
rect 405714 364618 405746 364854
rect 405982 364618 406066 364854
rect 406302 364618 406334 364854
rect 405714 328174 406334 364618
rect 405714 327938 405746 328174
rect 405982 327938 406066 328174
rect 406302 327938 406334 328174
rect 405714 327854 406334 327938
rect 405714 327618 405746 327854
rect 405982 327618 406066 327854
rect 406302 327618 406334 327854
rect 405714 291174 406334 327618
rect 405714 290938 405746 291174
rect 405982 290938 406066 291174
rect 406302 290938 406334 291174
rect 405714 290854 406334 290938
rect 405714 290618 405746 290854
rect 405982 290618 406066 290854
rect 406302 290618 406334 290854
rect 405714 254174 406334 290618
rect 405714 253938 405746 254174
rect 405982 253938 406066 254174
rect 406302 253938 406334 254174
rect 405714 253854 406334 253938
rect 405714 253618 405746 253854
rect 405982 253618 406066 253854
rect 406302 253618 406334 253854
rect 405714 217174 406334 253618
rect 405714 216938 405746 217174
rect 405982 216938 406066 217174
rect 406302 216938 406334 217174
rect 405714 216854 406334 216938
rect 405714 216618 405746 216854
rect 405982 216618 406066 216854
rect 406302 216618 406334 216854
rect 405714 180174 406334 216618
rect 405714 179938 405746 180174
rect 405982 179938 406066 180174
rect 406302 179938 406334 180174
rect 405714 179854 406334 179938
rect 405714 179618 405746 179854
rect 405982 179618 406066 179854
rect 406302 179618 406334 179854
rect 405714 143174 406334 179618
rect 405714 142938 405746 143174
rect 405982 142938 406066 143174
rect 406302 142938 406334 143174
rect 405714 142854 406334 142938
rect 405714 142618 405746 142854
rect 405982 142618 406066 142854
rect 406302 142618 406334 142854
rect 405714 106174 406334 142618
rect 405714 105938 405746 106174
rect 405982 105938 406066 106174
rect 406302 105938 406334 106174
rect 405714 105854 406334 105938
rect 405714 105618 405746 105854
rect 405982 105618 406066 105854
rect 406302 105618 406334 105854
rect 405714 69174 406334 105618
rect 405714 68938 405746 69174
rect 405982 68938 406066 69174
rect 406302 68938 406334 69174
rect 405714 68854 406334 68938
rect 405714 68618 405746 68854
rect 405982 68618 406066 68854
rect 406302 68618 406334 68854
rect 405714 32174 406334 68618
rect 405714 31938 405746 32174
rect 405982 31938 406066 32174
rect 406302 31938 406334 32174
rect 405714 31854 406334 31938
rect 405714 31618 405746 31854
rect 405982 31618 406066 31854
rect 406302 31618 406334 31854
rect 405714 -346 406334 31618
rect 405714 -582 405746 -346
rect 405982 -582 406066 -346
rect 406302 -582 406334 -346
rect 405714 -666 406334 -582
rect 405714 -902 405746 -666
rect 405982 -902 406066 -666
rect 406302 -902 406334 -666
rect 405714 -7654 406334 -902
rect 429994 705798 430614 711590
rect 429994 705562 430026 705798
rect 430262 705562 430346 705798
rect 430582 705562 430614 705798
rect 429994 705478 430614 705562
rect 429994 705242 430026 705478
rect 430262 705242 430346 705478
rect 430582 705242 430614 705478
rect 429994 694454 430614 705242
rect 429994 694218 430026 694454
rect 430262 694218 430346 694454
rect 430582 694218 430614 694454
rect 429994 694134 430614 694218
rect 429994 693898 430026 694134
rect 430262 693898 430346 694134
rect 430582 693898 430614 694134
rect 429994 657454 430614 693898
rect 429994 657218 430026 657454
rect 430262 657218 430346 657454
rect 430582 657218 430614 657454
rect 429994 657134 430614 657218
rect 429994 656898 430026 657134
rect 430262 656898 430346 657134
rect 430582 656898 430614 657134
rect 429994 620454 430614 656898
rect 429994 620218 430026 620454
rect 430262 620218 430346 620454
rect 430582 620218 430614 620454
rect 429994 620134 430614 620218
rect 429994 619898 430026 620134
rect 430262 619898 430346 620134
rect 430582 619898 430614 620134
rect 429994 583454 430614 619898
rect 429994 583218 430026 583454
rect 430262 583218 430346 583454
rect 430582 583218 430614 583454
rect 429994 583134 430614 583218
rect 429994 582898 430026 583134
rect 430262 582898 430346 583134
rect 430582 582898 430614 583134
rect 429994 546454 430614 582898
rect 429994 546218 430026 546454
rect 430262 546218 430346 546454
rect 430582 546218 430614 546454
rect 429994 546134 430614 546218
rect 429994 545898 430026 546134
rect 430262 545898 430346 546134
rect 430582 545898 430614 546134
rect 429994 509454 430614 545898
rect 429994 509218 430026 509454
rect 430262 509218 430346 509454
rect 430582 509218 430614 509454
rect 429994 509134 430614 509218
rect 429994 508898 430026 509134
rect 430262 508898 430346 509134
rect 430582 508898 430614 509134
rect 429994 472454 430614 508898
rect 429994 472218 430026 472454
rect 430262 472218 430346 472454
rect 430582 472218 430614 472454
rect 429994 472134 430614 472218
rect 429994 471898 430026 472134
rect 430262 471898 430346 472134
rect 430582 471898 430614 472134
rect 429994 435454 430614 471898
rect 429994 435218 430026 435454
rect 430262 435218 430346 435454
rect 430582 435218 430614 435454
rect 429994 435134 430614 435218
rect 429994 434898 430026 435134
rect 430262 434898 430346 435134
rect 430582 434898 430614 435134
rect 429994 398454 430614 434898
rect 429994 398218 430026 398454
rect 430262 398218 430346 398454
rect 430582 398218 430614 398454
rect 429994 398134 430614 398218
rect 429994 397898 430026 398134
rect 430262 397898 430346 398134
rect 430582 397898 430614 398134
rect 429994 361454 430614 397898
rect 429994 361218 430026 361454
rect 430262 361218 430346 361454
rect 430582 361218 430614 361454
rect 429994 361134 430614 361218
rect 429994 360898 430026 361134
rect 430262 360898 430346 361134
rect 430582 360898 430614 361134
rect 429994 324454 430614 360898
rect 429994 324218 430026 324454
rect 430262 324218 430346 324454
rect 430582 324218 430614 324454
rect 429994 324134 430614 324218
rect 429994 323898 430026 324134
rect 430262 323898 430346 324134
rect 430582 323898 430614 324134
rect 429994 287454 430614 323898
rect 429994 287218 430026 287454
rect 430262 287218 430346 287454
rect 430582 287218 430614 287454
rect 429994 287134 430614 287218
rect 429994 286898 430026 287134
rect 430262 286898 430346 287134
rect 430582 286898 430614 287134
rect 429994 250454 430614 286898
rect 429994 250218 430026 250454
rect 430262 250218 430346 250454
rect 430582 250218 430614 250454
rect 429994 250134 430614 250218
rect 429994 249898 430026 250134
rect 430262 249898 430346 250134
rect 430582 249898 430614 250134
rect 429994 213454 430614 249898
rect 429994 213218 430026 213454
rect 430262 213218 430346 213454
rect 430582 213218 430614 213454
rect 429994 213134 430614 213218
rect 429994 212898 430026 213134
rect 430262 212898 430346 213134
rect 430582 212898 430614 213134
rect 429994 176454 430614 212898
rect 429994 176218 430026 176454
rect 430262 176218 430346 176454
rect 430582 176218 430614 176454
rect 429994 176134 430614 176218
rect 429994 175898 430026 176134
rect 430262 175898 430346 176134
rect 430582 175898 430614 176134
rect 429994 139454 430614 175898
rect 429994 139218 430026 139454
rect 430262 139218 430346 139454
rect 430582 139218 430614 139454
rect 429994 139134 430614 139218
rect 429994 138898 430026 139134
rect 430262 138898 430346 139134
rect 430582 138898 430614 139134
rect 429994 102454 430614 138898
rect 429994 102218 430026 102454
rect 430262 102218 430346 102454
rect 430582 102218 430614 102454
rect 429994 102134 430614 102218
rect 429994 101898 430026 102134
rect 430262 101898 430346 102134
rect 430582 101898 430614 102134
rect 429994 65454 430614 101898
rect 429994 65218 430026 65454
rect 430262 65218 430346 65454
rect 430582 65218 430614 65454
rect 429994 65134 430614 65218
rect 429994 64898 430026 65134
rect 430262 64898 430346 65134
rect 430582 64898 430614 65134
rect 429994 28454 430614 64898
rect 429994 28218 430026 28454
rect 430262 28218 430346 28454
rect 430582 28218 430614 28454
rect 429994 28134 430614 28218
rect 429994 27898 430026 28134
rect 430262 27898 430346 28134
rect 430582 27898 430614 28134
rect 429994 -1306 430614 27898
rect 429994 -1542 430026 -1306
rect 430262 -1542 430346 -1306
rect 430582 -1542 430614 -1306
rect 429994 -1626 430614 -1542
rect 429994 -1862 430026 -1626
rect 430262 -1862 430346 -1626
rect 430582 -1862 430614 -1626
rect 429994 -7654 430614 -1862
rect 433714 704838 434334 711590
rect 433714 704602 433746 704838
rect 433982 704602 434066 704838
rect 434302 704602 434334 704838
rect 433714 704518 434334 704602
rect 433714 704282 433746 704518
rect 433982 704282 434066 704518
rect 434302 704282 434334 704518
rect 433714 698174 434334 704282
rect 433714 697938 433746 698174
rect 433982 697938 434066 698174
rect 434302 697938 434334 698174
rect 433714 697854 434334 697938
rect 433714 697618 433746 697854
rect 433982 697618 434066 697854
rect 434302 697618 434334 697854
rect 433714 661174 434334 697618
rect 433714 660938 433746 661174
rect 433982 660938 434066 661174
rect 434302 660938 434334 661174
rect 433714 660854 434334 660938
rect 433714 660618 433746 660854
rect 433982 660618 434066 660854
rect 434302 660618 434334 660854
rect 433714 624174 434334 660618
rect 433714 623938 433746 624174
rect 433982 623938 434066 624174
rect 434302 623938 434334 624174
rect 433714 623854 434334 623938
rect 433714 623618 433746 623854
rect 433982 623618 434066 623854
rect 434302 623618 434334 623854
rect 433714 587174 434334 623618
rect 433714 586938 433746 587174
rect 433982 586938 434066 587174
rect 434302 586938 434334 587174
rect 433714 586854 434334 586938
rect 433714 586618 433746 586854
rect 433982 586618 434066 586854
rect 434302 586618 434334 586854
rect 433714 550174 434334 586618
rect 433714 549938 433746 550174
rect 433982 549938 434066 550174
rect 434302 549938 434334 550174
rect 433714 549854 434334 549938
rect 433714 549618 433746 549854
rect 433982 549618 434066 549854
rect 434302 549618 434334 549854
rect 433714 513174 434334 549618
rect 433714 512938 433746 513174
rect 433982 512938 434066 513174
rect 434302 512938 434334 513174
rect 433714 512854 434334 512938
rect 433714 512618 433746 512854
rect 433982 512618 434066 512854
rect 434302 512618 434334 512854
rect 433714 476174 434334 512618
rect 433714 475938 433746 476174
rect 433982 475938 434066 476174
rect 434302 475938 434334 476174
rect 433714 475854 434334 475938
rect 433714 475618 433746 475854
rect 433982 475618 434066 475854
rect 434302 475618 434334 475854
rect 433714 439174 434334 475618
rect 433714 438938 433746 439174
rect 433982 438938 434066 439174
rect 434302 438938 434334 439174
rect 433714 438854 434334 438938
rect 433714 438618 433746 438854
rect 433982 438618 434066 438854
rect 434302 438618 434334 438854
rect 433714 402174 434334 438618
rect 433714 401938 433746 402174
rect 433982 401938 434066 402174
rect 434302 401938 434334 402174
rect 433714 401854 434334 401938
rect 433714 401618 433746 401854
rect 433982 401618 434066 401854
rect 434302 401618 434334 401854
rect 433714 365174 434334 401618
rect 433714 364938 433746 365174
rect 433982 364938 434066 365174
rect 434302 364938 434334 365174
rect 433714 364854 434334 364938
rect 433714 364618 433746 364854
rect 433982 364618 434066 364854
rect 434302 364618 434334 364854
rect 433714 328174 434334 364618
rect 433714 327938 433746 328174
rect 433982 327938 434066 328174
rect 434302 327938 434334 328174
rect 433714 327854 434334 327938
rect 433714 327618 433746 327854
rect 433982 327618 434066 327854
rect 434302 327618 434334 327854
rect 433714 291174 434334 327618
rect 433714 290938 433746 291174
rect 433982 290938 434066 291174
rect 434302 290938 434334 291174
rect 433714 290854 434334 290938
rect 433714 290618 433746 290854
rect 433982 290618 434066 290854
rect 434302 290618 434334 290854
rect 433714 254174 434334 290618
rect 433714 253938 433746 254174
rect 433982 253938 434066 254174
rect 434302 253938 434334 254174
rect 433714 253854 434334 253938
rect 433714 253618 433746 253854
rect 433982 253618 434066 253854
rect 434302 253618 434334 253854
rect 433714 217174 434334 253618
rect 433714 216938 433746 217174
rect 433982 216938 434066 217174
rect 434302 216938 434334 217174
rect 433714 216854 434334 216938
rect 433714 216618 433746 216854
rect 433982 216618 434066 216854
rect 434302 216618 434334 216854
rect 433714 180174 434334 216618
rect 433714 179938 433746 180174
rect 433982 179938 434066 180174
rect 434302 179938 434334 180174
rect 433714 179854 434334 179938
rect 433714 179618 433746 179854
rect 433982 179618 434066 179854
rect 434302 179618 434334 179854
rect 433714 143174 434334 179618
rect 433714 142938 433746 143174
rect 433982 142938 434066 143174
rect 434302 142938 434334 143174
rect 433714 142854 434334 142938
rect 433714 142618 433746 142854
rect 433982 142618 434066 142854
rect 434302 142618 434334 142854
rect 433714 106174 434334 142618
rect 433714 105938 433746 106174
rect 433982 105938 434066 106174
rect 434302 105938 434334 106174
rect 433714 105854 434334 105938
rect 433714 105618 433746 105854
rect 433982 105618 434066 105854
rect 434302 105618 434334 105854
rect 433714 69174 434334 105618
rect 433714 68938 433746 69174
rect 433982 68938 434066 69174
rect 434302 68938 434334 69174
rect 433714 68854 434334 68938
rect 433714 68618 433746 68854
rect 433982 68618 434066 68854
rect 434302 68618 434334 68854
rect 433714 32174 434334 68618
rect 433714 31938 433746 32174
rect 433982 31938 434066 32174
rect 434302 31938 434334 32174
rect 433714 31854 434334 31938
rect 433714 31618 433746 31854
rect 433982 31618 434066 31854
rect 434302 31618 434334 31854
rect 433714 -346 434334 31618
rect 433714 -582 433746 -346
rect 433982 -582 434066 -346
rect 434302 -582 434334 -346
rect 433714 -666 434334 -582
rect 433714 -902 433746 -666
rect 433982 -902 434066 -666
rect 434302 -902 434334 -666
rect 433714 -7654 434334 -902
rect 457994 705798 458614 711590
rect 457994 705562 458026 705798
rect 458262 705562 458346 705798
rect 458582 705562 458614 705798
rect 457994 705478 458614 705562
rect 457994 705242 458026 705478
rect 458262 705242 458346 705478
rect 458582 705242 458614 705478
rect 457994 694454 458614 705242
rect 457994 694218 458026 694454
rect 458262 694218 458346 694454
rect 458582 694218 458614 694454
rect 457994 694134 458614 694218
rect 457994 693898 458026 694134
rect 458262 693898 458346 694134
rect 458582 693898 458614 694134
rect 457994 657454 458614 693898
rect 457994 657218 458026 657454
rect 458262 657218 458346 657454
rect 458582 657218 458614 657454
rect 457994 657134 458614 657218
rect 457994 656898 458026 657134
rect 458262 656898 458346 657134
rect 458582 656898 458614 657134
rect 457994 620454 458614 656898
rect 457994 620218 458026 620454
rect 458262 620218 458346 620454
rect 458582 620218 458614 620454
rect 457994 620134 458614 620218
rect 457994 619898 458026 620134
rect 458262 619898 458346 620134
rect 458582 619898 458614 620134
rect 457994 583454 458614 619898
rect 457994 583218 458026 583454
rect 458262 583218 458346 583454
rect 458582 583218 458614 583454
rect 457994 583134 458614 583218
rect 457994 582898 458026 583134
rect 458262 582898 458346 583134
rect 458582 582898 458614 583134
rect 457994 546454 458614 582898
rect 457994 546218 458026 546454
rect 458262 546218 458346 546454
rect 458582 546218 458614 546454
rect 457994 546134 458614 546218
rect 457994 545898 458026 546134
rect 458262 545898 458346 546134
rect 458582 545898 458614 546134
rect 457994 509454 458614 545898
rect 457994 509218 458026 509454
rect 458262 509218 458346 509454
rect 458582 509218 458614 509454
rect 457994 509134 458614 509218
rect 457994 508898 458026 509134
rect 458262 508898 458346 509134
rect 458582 508898 458614 509134
rect 457994 472454 458614 508898
rect 457994 472218 458026 472454
rect 458262 472218 458346 472454
rect 458582 472218 458614 472454
rect 457994 472134 458614 472218
rect 457994 471898 458026 472134
rect 458262 471898 458346 472134
rect 458582 471898 458614 472134
rect 457994 435454 458614 471898
rect 457994 435218 458026 435454
rect 458262 435218 458346 435454
rect 458582 435218 458614 435454
rect 457994 435134 458614 435218
rect 457994 434898 458026 435134
rect 458262 434898 458346 435134
rect 458582 434898 458614 435134
rect 457994 398454 458614 434898
rect 457994 398218 458026 398454
rect 458262 398218 458346 398454
rect 458582 398218 458614 398454
rect 457994 398134 458614 398218
rect 457994 397898 458026 398134
rect 458262 397898 458346 398134
rect 458582 397898 458614 398134
rect 457994 361454 458614 397898
rect 457994 361218 458026 361454
rect 458262 361218 458346 361454
rect 458582 361218 458614 361454
rect 457994 361134 458614 361218
rect 457994 360898 458026 361134
rect 458262 360898 458346 361134
rect 458582 360898 458614 361134
rect 457994 324454 458614 360898
rect 457994 324218 458026 324454
rect 458262 324218 458346 324454
rect 458582 324218 458614 324454
rect 457994 324134 458614 324218
rect 457994 323898 458026 324134
rect 458262 323898 458346 324134
rect 458582 323898 458614 324134
rect 457994 287454 458614 323898
rect 457994 287218 458026 287454
rect 458262 287218 458346 287454
rect 458582 287218 458614 287454
rect 457994 287134 458614 287218
rect 457994 286898 458026 287134
rect 458262 286898 458346 287134
rect 458582 286898 458614 287134
rect 457994 250454 458614 286898
rect 457994 250218 458026 250454
rect 458262 250218 458346 250454
rect 458582 250218 458614 250454
rect 457994 250134 458614 250218
rect 457994 249898 458026 250134
rect 458262 249898 458346 250134
rect 458582 249898 458614 250134
rect 457994 213454 458614 249898
rect 457994 213218 458026 213454
rect 458262 213218 458346 213454
rect 458582 213218 458614 213454
rect 457994 213134 458614 213218
rect 457994 212898 458026 213134
rect 458262 212898 458346 213134
rect 458582 212898 458614 213134
rect 457994 176454 458614 212898
rect 457994 176218 458026 176454
rect 458262 176218 458346 176454
rect 458582 176218 458614 176454
rect 457994 176134 458614 176218
rect 457994 175898 458026 176134
rect 458262 175898 458346 176134
rect 458582 175898 458614 176134
rect 457994 139454 458614 175898
rect 457994 139218 458026 139454
rect 458262 139218 458346 139454
rect 458582 139218 458614 139454
rect 457994 139134 458614 139218
rect 457994 138898 458026 139134
rect 458262 138898 458346 139134
rect 458582 138898 458614 139134
rect 457994 102454 458614 138898
rect 457994 102218 458026 102454
rect 458262 102218 458346 102454
rect 458582 102218 458614 102454
rect 457994 102134 458614 102218
rect 457994 101898 458026 102134
rect 458262 101898 458346 102134
rect 458582 101898 458614 102134
rect 457994 65454 458614 101898
rect 457994 65218 458026 65454
rect 458262 65218 458346 65454
rect 458582 65218 458614 65454
rect 457994 65134 458614 65218
rect 457994 64898 458026 65134
rect 458262 64898 458346 65134
rect 458582 64898 458614 65134
rect 457994 28454 458614 64898
rect 457994 28218 458026 28454
rect 458262 28218 458346 28454
rect 458582 28218 458614 28454
rect 457994 28134 458614 28218
rect 457994 27898 458026 28134
rect 458262 27898 458346 28134
rect 458582 27898 458614 28134
rect 457994 -1306 458614 27898
rect 457994 -1542 458026 -1306
rect 458262 -1542 458346 -1306
rect 458582 -1542 458614 -1306
rect 457994 -1626 458614 -1542
rect 457994 -1862 458026 -1626
rect 458262 -1862 458346 -1626
rect 458582 -1862 458614 -1626
rect 457994 -7654 458614 -1862
rect 461714 704838 462334 711590
rect 461714 704602 461746 704838
rect 461982 704602 462066 704838
rect 462302 704602 462334 704838
rect 461714 704518 462334 704602
rect 461714 704282 461746 704518
rect 461982 704282 462066 704518
rect 462302 704282 462334 704518
rect 461714 698174 462334 704282
rect 461714 697938 461746 698174
rect 461982 697938 462066 698174
rect 462302 697938 462334 698174
rect 461714 697854 462334 697938
rect 461714 697618 461746 697854
rect 461982 697618 462066 697854
rect 462302 697618 462334 697854
rect 461714 661174 462334 697618
rect 461714 660938 461746 661174
rect 461982 660938 462066 661174
rect 462302 660938 462334 661174
rect 461714 660854 462334 660938
rect 461714 660618 461746 660854
rect 461982 660618 462066 660854
rect 462302 660618 462334 660854
rect 461714 624174 462334 660618
rect 461714 623938 461746 624174
rect 461982 623938 462066 624174
rect 462302 623938 462334 624174
rect 461714 623854 462334 623938
rect 461714 623618 461746 623854
rect 461982 623618 462066 623854
rect 462302 623618 462334 623854
rect 461714 587174 462334 623618
rect 461714 586938 461746 587174
rect 461982 586938 462066 587174
rect 462302 586938 462334 587174
rect 461714 586854 462334 586938
rect 461714 586618 461746 586854
rect 461982 586618 462066 586854
rect 462302 586618 462334 586854
rect 461714 550174 462334 586618
rect 461714 549938 461746 550174
rect 461982 549938 462066 550174
rect 462302 549938 462334 550174
rect 461714 549854 462334 549938
rect 461714 549618 461746 549854
rect 461982 549618 462066 549854
rect 462302 549618 462334 549854
rect 461714 513174 462334 549618
rect 461714 512938 461746 513174
rect 461982 512938 462066 513174
rect 462302 512938 462334 513174
rect 461714 512854 462334 512938
rect 461714 512618 461746 512854
rect 461982 512618 462066 512854
rect 462302 512618 462334 512854
rect 461714 476174 462334 512618
rect 461714 475938 461746 476174
rect 461982 475938 462066 476174
rect 462302 475938 462334 476174
rect 461714 475854 462334 475938
rect 461714 475618 461746 475854
rect 461982 475618 462066 475854
rect 462302 475618 462334 475854
rect 461714 439174 462334 475618
rect 461714 438938 461746 439174
rect 461982 438938 462066 439174
rect 462302 438938 462334 439174
rect 461714 438854 462334 438938
rect 461714 438618 461746 438854
rect 461982 438618 462066 438854
rect 462302 438618 462334 438854
rect 461714 402174 462334 438618
rect 461714 401938 461746 402174
rect 461982 401938 462066 402174
rect 462302 401938 462334 402174
rect 461714 401854 462334 401938
rect 461714 401618 461746 401854
rect 461982 401618 462066 401854
rect 462302 401618 462334 401854
rect 461714 365174 462334 401618
rect 461714 364938 461746 365174
rect 461982 364938 462066 365174
rect 462302 364938 462334 365174
rect 461714 364854 462334 364938
rect 461714 364618 461746 364854
rect 461982 364618 462066 364854
rect 462302 364618 462334 364854
rect 461714 328174 462334 364618
rect 461714 327938 461746 328174
rect 461982 327938 462066 328174
rect 462302 327938 462334 328174
rect 461714 327854 462334 327938
rect 461714 327618 461746 327854
rect 461982 327618 462066 327854
rect 462302 327618 462334 327854
rect 461714 291174 462334 327618
rect 461714 290938 461746 291174
rect 461982 290938 462066 291174
rect 462302 290938 462334 291174
rect 461714 290854 462334 290938
rect 461714 290618 461746 290854
rect 461982 290618 462066 290854
rect 462302 290618 462334 290854
rect 461714 254174 462334 290618
rect 461714 253938 461746 254174
rect 461982 253938 462066 254174
rect 462302 253938 462334 254174
rect 461714 253854 462334 253938
rect 461714 253618 461746 253854
rect 461982 253618 462066 253854
rect 462302 253618 462334 253854
rect 461714 217174 462334 253618
rect 461714 216938 461746 217174
rect 461982 216938 462066 217174
rect 462302 216938 462334 217174
rect 461714 216854 462334 216938
rect 461714 216618 461746 216854
rect 461982 216618 462066 216854
rect 462302 216618 462334 216854
rect 461714 180174 462334 216618
rect 461714 179938 461746 180174
rect 461982 179938 462066 180174
rect 462302 179938 462334 180174
rect 461714 179854 462334 179938
rect 461714 179618 461746 179854
rect 461982 179618 462066 179854
rect 462302 179618 462334 179854
rect 461714 143174 462334 179618
rect 461714 142938 461746 143174
rect 461982 142938 462066 143174
rect 462302 142938 462334 143174
rect 461714 142854 462334 142938
rect 461714 142618 461746 142854
rect 461982 142618 462066 142854
rect 462302 142618 462334 142854
rect 461714 106174 462334 142618
rect 461714 105938 461746 106174
rect 461982 105938 462066 106174
rect 462302 105938 462334 106174
rect 461714 105854 462334 105938
rect 461714 105618 461746 105854
rect 461982 105618 462066 105854
rect 462302 105618 462334 105854
rect 461714 69174 462334 105618
rect 461714 68938 461746 69174
rect 461982 68938 462066 69174
rect 462302 68938 462334 69174
rect 461714 68854 462334 68938
rect 461714 68618 461746 68854
rect 461982 68618 462066 68854
rect 462302 68618 462334 68854
rect 461714 32174 462334 68618
rect 461714 31938 461746 32174
rect 461982 31938 462066 32174
rect 462302 31938 462334 32174
rect 461714 31854 462334 31938
rect 461714 31618 461746 31854
rect 461982 31618 462066 31854
rect 462302 31618 462334 31854
rect 461714 -346 462334 31618
rect 461714 -582 461746 -346
rect 461982 -582 462066 -346
rect 462302 -582 462334 -346
rect 461714 -666 462334 -582
rect 461714 -902 461746 -666
rect 461982 -902 462066 -666
rect 462302 -902 462334 -666
rect 461714 -7654 462334 -902
rect 485994 705798 486614 711590
rect 485994 705562 486026 705798
rect 486262 705562 486346 705798
rect 486582 705562 486614 705798
rect 485994 705478 486614 705562
rect 485994 705242 486026 705478
rect 486262 705242 486346 705478
rect 486582 705242 486614 705478
rect 485994 694454 486614 705242
rect 485994 694218 486026 694454
rect 486262 694218 486346 694454
rect 486582 694218 486614 694454
rect 485994 694134 486614 694218
rect 485994 693898 486026 694134
rect 486262 693898 486346 694134
rect 486582 693898 486614 694134
rect 485994 657454 486614 693898
rect 485994 657218 486026 657454
rect 486262 657218 486346 657454
rect 486582 657218 486614 657454
rect 485994 657134 486614 657218
rect 485994 656898 486026 657134
rect 486262 656898 486346 657134
rect 486582 656898 486614 657134
rect 485994 620454 486614 656898
rect 485994 620218 486026 620454
rect 486262 620218 486346 620454
rect 486582 620218 486614 620454
rect 485994 620134 486614 620218
rect 485994 619898 486026 620134
rect 486262 619898 486346 620134
rect 486582 619898 486614 620134
rect 485994 583454 486614 619898
rect 485994 583218 486026 583454
rect 486262 583218 486346 583454
rect 486582 583218 486614 583454
rect 485994 583134 486614 583218
rect 485994 582898 486026 583134
rect 486262 582898 486346 583134
rect 486582 582898 486614 583134
rect 485994 546454 486614 582898
rect 485994 546218 486026 546454
rect 486262 546218 486346 546454
rect 486582 546218 486614 546454
rect 485994 546134 486614 546218
rect 485994 545898 486026 546134
rect 486262 545898 486346 546134
rect 486582 545898 486614 546134
rect 485994 509454 486614 545898
rect 485994 509218 486026 509454
rect 486262 509218 486346 509454
rect 486582 509218 486614 509454
rect 485994 509134 486614 509218
rect 485994 508898 486026 509134
rect 486262 508898 486346 509134
rect 486582 508898 486614 509134
rect 485994 472454 486614 508898
rect 485994 472218 486026 472454
rect 486262 472218 486346 472454
rect 486582 472218 486614 472454
rect 485994 472134 486614 472218
rect 485994 471898 486026 472134
rect 486262 471898 486346 472134
rect 486582 471898 486614 472134
rect 485994 435454 486614 471898
rect 485994 435218 486026 435454
rect 486262 435218 486346 435454
rect 486582 435218 486614 435454
rect 485994 435134 486614 435218
rect 485994 434898 486026 435134
rect 486262 434898 486346 435134
rect 486582 434898 486614 435134
rect 485994 398454 486614 434898
rect 485994 398218 486026 398454
rect 486262 398218 486346 398454
rect 486582 398218 486614 398454
rect 485994 398134 486614 398218
rect 485994 397898 486026 398134
rect 486262 397898 486346 398134
rect 486582 397898 486614 398134
rect 485994 361454 486614 397898
rect 485994 361218 486026 361454
rect 486262 361218 486346 361454
rect 486582 361218 486614 361454
rect 485994 361134 486614 361218
rect 485994 360898 486026 361134
rect 486262 360898 486346 361134
rect 486582 360898 486614 361134
rect 485994 324454 486614 360898
rect 485994 324218 486026 324454
rect 486262 324218 486346 324454
rect 486582 324218 486614 324454
rect 485994 324134 486614 324218
rect 485994 323898 486026 324134
rect 486262 323898 486346 324134
rect 486582 323898 486614 324134
rect 485994 287454 486614 323898
rect 485994 287218 486026 287454
rect 486262 287218 486346 287454
rect 486582 287218 486614 287454
rect 485994 287134 486614 287218
rect 485994 286898 486026 287134
rect 486262 286898 486346 287134
rect 486582 286898 486614 287134
rect 485994 250454 486614 286898
rect 485994 250218 486026 250454
rect 486262 250218 486346 250454
rect 486582 250218 486614 250454
rect 485994 250134 486614 250218
rect 485994 249898 486026 250134
rect 486262 249898 486346 250134
rect 486582 249898 486614 250134
rect 485994 213454 486614 249898
rect 485994 213218 486026 213454
rect 486262 213218 486346 213454
rect 486582 213218 486614 213454
rect 485994 213134 486614 213218
rect 485994 212898 486026 213134
rect 486262 212898 486346 213134
rect 486582 212898 486614 213134
rect 485994 176454 486614 212898
rect 485994 176218 486026 176454
rect 486262 176218 486346 176454
rect 486582 176218 486614 176454
rect 485994 176134 486614 176218
rect 485994 175898 486026 176134
rect 486262 175898 486346 176134
rect 486582 175898 486614 176134
rect 485994 139454 486614 175898
rect 485994 139218 486026 139454
rect 486262 139218 486346 139454
rect 486582 139218 486614 139454
rect 485994 139134 486614 139218
rect 485994 138898 486026 139134
rect 486262 138898 486346 139134
rect 486582 138898 486614 139134
rect 485994 102454 486614 138898
rect 485994 102218 486026 102454
rect 486262 102218 486346 102454
rect 486582 102218 486614 102454
rect 485994 102134 486614 102218
rect 485994 101898 486026 102134
rect 486262 101898 486346 102134
rect 486582 101898 486614 102134
rect 485994 65454 486614 101898
rect 485994 65218 486026 65454
rect 486262 65218 486346 65454
rect 486582 65218 486614 65454
rect 485994 65134 486614 65218
rect 485994 64898 486026 65134
rect 486262 64898 486346 65134
rect 486582 64898 486614 65134
rect 485994 28454 486614 64898
rect 485994 28218 486026 28454
rect 486262 28218 486346 28454
rect 486582 28218 486614 28454
rect 485994 28134 486614 28218
rect 485994 27898 486026 28134
rect 486262 27898 486346 28134
rect 486582 27898 486614 28134
rect 485994 -1306 486614 27898
rect 485994 -1542 486026 -1306
rect 486262 -1542 486346 -1306
rect 486582 -1542 486614 -1306
rect 485994 -1626 486614 -1542
rect 485994 -1862 486026 -1626
rect 486262 -1862 486346 -1626
rect 486582 -1862 486614 -1626
rect 485994 -7654 486614 -1862
rect 489714 704838 490334 711590
rect 489714 704602 489746 704838
rect 489982 704602 490066 704838
rect 490302 704602 490334 704838
rect 489714 704518 490334 704602
rect 489714 704282 489746 704518
rect 489982 704282 490066 704518
rect 490302 704282 490334 704518
rect 489714 698174 490334 704282
rect 489714 697938 489746 698174
rect 489982 697938 490066 698174
rect 490302 697938 490334 698174
rect 489714 697854 490334 697938
rect 489714 697618 489746 697854
rect 489982 697618 490066 697854
rect 490302 697618 490334 697854
rect 489714 661174 490334 697618
rect 489714 660938 489746 661174
rect 489982 660938 490066 661174
rect 490302 660938 490334 661174
rect 489714 660854 490334 660938
rect 489714 660618 489746 660854
rect 489982 660618 490066 660854
rect 490302 660618 490334 660854
rect 489714 624174 490334 660618
rect 489714 623938 489746 624174
rect 489982 623938 490066 624174
rect 490302 623938 490334 624174
rect 489714 623854 490334 623938
rect 489714 623618 489746 623854
rect 489982 623618 490066 623854
rect 490302 623618 490334 623854
rect 489714 587174 490334 623618
rect 489714 586938 489746 587174
rect 489982 586938 490066 587174
rect 490302 586938 490334 587174
rect 489714 586854 490334 586938
rect 489714 586618 489746 586854
rect 489982 586618 490066 586854
rect 490302 586618 490334 586854
rect 489714 550174 490334 586618
rect 489714 549938 489746 550174
rect 489982 549938 490066 550174
rect 490302 549938 490334 550174
rect 489714 549854 490334 549938
rect 489714 549618 489746 549854
rect 489982 549618 490066 549854
rect 490302 549618 490334 549854
rect 489714 513174 490334 549618
rect 489714 512938 489746 513174
rect 489982 512938 490066 513174
rect 490302 512938 490334 513174
rect 489714 512854 490334 512938
rect 489714 512618 489746 512854
rect 489982 512618 490066 512854
rect 490302 512618 490334 512854
rect 489714 476174 490334 512618
rect 489714 475938 489746 476174
rect 489982 475938 490066 476174
rect 490302 475938 490334 476174
rect 489714 475854 490334 475938
rect 489714 475618 489746 475854
rect 489982 475618 490066 475854
rect 490302 475618 490334 475854
rect 489714 439174 490334 475618
rect 489714 438938 489746 439174
rect 489982 438938 490066 439174
rect 490302 438938 490334 439174
rect 489714 438854 490334 438938
rect 489714 438618 489746 438854
rect 489982 438618 490066 438854
rect 490302 438618 490334 438854
rect 489714 402174 490334 438618
rect 489714 401938 489746 402174
rect 489982 401938 490066 402174
rect 490302 401938 490334 402174
rect 489714 401854 490334 401938
rect 489714 401618 489746 401854
rect 489982 401618 490066 401854
rect 490302 401618 490334 401854
rect 489714 365174 490334 401618
rect 489714 364938 489746 365174
rect 489982 364938 490066 365174
rect 490302 364938 490334 365174
rect 489714 364854 490334 364938
rect 489714 364618 489746 364854
rect 489982 364618 490066 364854
rect 490302 364618 490334 364854
rect 489714 328174 490334 364618
rect 489714 327938 489746 328174
rect 489982 327938 490066 328174
rect 490302 327938 490334 328174
rect 489714 327854 490334 327938
rect 489714 327618 489746 327854
rect 489982 327618 490066 327854
rect 490302 327618 490334 327854
rect 489714 291174 490334 327618
rect 489714 290938 489746 291174
rect 489982 290938 490066 291174
rect 490302 290938 490334 291174
rect 489714 290854 490334 290938
rect 489714 290618 489746 290854
rect 489982 290618 490066 290854
rect 490302 290618 490334 290854
rect 489714 254174 490334 290618
rect 489714 253938 489746 254174
rect 489982 253938 490066 254174
rect 490302 253938 490334 254174
rect 489714 253854 490334 253938
rect 489714 253618 489746 253854
rect 489982 253618 490066 253854
rect 490302 253618 490334 253854
rect 489714 217174 490334 253618
rect 489714 216938 489746 217174
rect 489982 216938 490066 217174
rect 490302 216938 490334 217174
rect 489714 216854 490334 216938
rect 489714 216618 489746 216854
rect 489982 216618 490066 216854
rect 490302 216618 490334 216854
rect 489714 180174 490334 216618
rect 489714 179938 489746 180174
rect 489982 179938 490066 180174
rect 490302 179938 490334 180174
rect 489714 179854 490334 179938
rect 489714 179618 489746 179854
rect 489982 179618 490066 179854
rect 490302 179618 490334 179854
rect 489714 143174 490334 179618
rect 489714 142938 489746 143174
rect 489982 142938 490066 143174
rect 490302 142938 490334 143174
rect 489714 142854 490334 142938
rect 489714 142618 489746 142854
rect 489982 142618 490066 142854
rect 490302 142618 490334 142854
rect 489714 106174 490334 142618
rect 489714 105938 489746 106174
rect 489982 105938 490066 106174
rect 490302 105938 490334 106174
rect 489714 105854 490334 105938
rect 489714 105618 489746 105854
rect 489982 105618 490066 105854
rect 490302 105618 490334 105854
rect 489714 69174 490334 105618
rect 489714 68938 489746 69174
rect 489982 68938 490066 69174
rect 490302 68938 490334 69174
rect 489714 68854 490334 68938
rect 489714 68618 489746 68854
rect 489982 68618 490066 68854
rect 490302 68618 490334 68854
rect 489714 32174 490334 68618
rect 489714 31938 489746 32174
rect 489982 31938 490066 32174
rect 490302 31938 490334 32174
rect 489714 31854 490334 31938
rect 489714 31618 489746 31854
rect 489982 31618 490066 31854
rect 490302 31618 490334 31854
rect 489714 -346 490334 31618
rect 489714 -582 489746 -346
rect 489982 -582 490066 -346
rect 490302 -582 490334 -346
rect 489714 -666 490334 -582
rect 489714 -902 489746 -666
rect 489982 -902 490066 -666
rect 490302 -902 490334 -666
rect 489714 -7654 490334 -902
rect 513994 705798 514614 711590
rect 513994 705562 514026 705798
rect 514262 705562 514346 705798
rect 514582 705562 514614 705798
rect 513994 705478 514614 705562
rect 513994 705242 514026 705478
rect 514262 705242 514346 705478
rect 514582 705242 514614 705478
rect 513994 694454 514614 705242
rect 513994 694218 514026 694454
rect 514262 694218 514346 694454
rect 514582 694218 514614 694454
rect 513994 694134 514614 694218
rect 513994 693898 514026 694134
rect 514262 693898 514346 694134
rect 514582 693898 514614 694134
rect 513994 657454 514614 693898
rect 513994 657218 514026 657454
rect 514262 657218 514346 657454
rect 514582 657218 514614 657454
rect 513994 657134 514614 657218
rect 513994 656898 514026 657134
rect 514262 656898 514346 657134
rect 514582 656898 514614 657134
rect 513994 620454 514614 656898
rect 513994 620218 514026 620454
rect 514262 620218 514346 620454
rect 514582 620218 514614 620454
rect 513994 620134 514614 620218
rect 513994 619898 514026 620134
rect 514262 619898 514346 620134
rect 514582 619898 514614 620134
rect 513994 583454 514614 619898
rect 513994 583218 514026 583454
rect 514262 583218 514346 583454
rect 514582 583218 514614 583454
rect 513994 583134 514614 583218
rect 513994 582898 514026 583134
rect 514262 582898 514346 583134
rect 514582 582898 514614 583134
rect 513994 546454 514614 582898
rect 513994 546218 514026 546454
rect 514262 546218 514346 546454
rect 514582 546218 514614 546454
rect 513994 546134 514614 546218
rect 513994 545898 514026 546134
rect 514262 545898 514346 546134
rect 514582 545898 514614 546134
rect 513994 509454 514614 545898
rect 513994 509218 514026 509454
rect 514262 509218 514346 509454
rect 514582 509218 514614 509454
rect 513994 509134 514614 509218
rect 513994 508898 514026 509134
rect 514262 508898 514346 509134
rect 514582 508898 514614 509134
rect 513994 472454 514614 508898
rect 513994 472218 514026 472454
rect 514262 472218 514346 472454
rect 514582 472218 514614 472454
rect 513994 472134 514614 472218
rect 513994 471898 514026 472134
rect 514262 471898 514346 472134
rect 514582 471898 514614 472134
rect 513994 435454 514614 471898
rect 513994 435218 514026 435454
rect 514262 435218 514346 435454
rect 514582 435218 514614 435454
rect 513994 435134 514614 435218
rect 513994 434898 514026 435134
rect 514262 434898 514346 435134
rect 514582 434898 514614 435134
rect 513994 398454 514614 434898
rect 513994 398218 514026 398454
rect 514262 398218 514346 398454
rect 514582 398218 514614 398454
rect 513994 398134 514614 398218
rect 513994 397898 514026 398134
rect 514262 397898 514346 398134
rect 514582 397898 514614 398134
rect 513994 361454 514614 397898
rect 513994 361218 514026 361454
rect 514262 361218 514346 361454
rect 514582 361218 514614 361454
rect 513994 361134 514614 361218
rect 513994 360898 514026 361134
rect 514262 360898 514346 361134
rect 514582 360898 514614 361134
rect 513994 324454 514614 360898
rect 513994 324218 514026 324454
rect 514262 324218 514346 324454
rect 514582 324218 514614 324454
rect 513994 324134 514614 324218
rect 513994 323898 514026 324134
rect 514262 323898 514346 324134
rect 514582 323898 514614 324134
rect 513994 287454 514614 323898
rect 513994 287218 514026 287454
rect 514262 287218 514346 287454
rect 514582 287218 514614 287454
rect 513994 287134 514614 287218
rect 513994 286898 514026 287134
rect 514262 286898 514346 287134
rect 514582 286898 514614 287134
rect 513994 250454 514614 286898
rect 513994 250218 514026 250454
rect 514262 250218 514346 250454
rect 514582 250218 514614 250454
rect 513994 250134 514614 250218
rect 513994 249898 514026 250134
rect 514262 249898 514346 250134
rect 514582 249898 514614 250134
rect 513994 213454 514614 249898
rect 513994 213218 514026 213454
rect 514262 213218 514346 213454
rect 514582 213218 514614 213454
rect 513994 213134 514614 213218
rect 513994 212898 514026 213134
rect 514262 212898 514346 213134
rect 514582 212898 514614 213134
rect 513994 176454 514614 212898
rect 513994 176218 514026 176454
rect 514262 176218 514346 176454
rect 514582 176218 514614 176454
rect 513994 176134 514614 176218
rect 513994 175898 514026 176134
rect 514262 175898 514346 176134
rect 514582 175898 514614 176134
rect 513994 139454 514614 175898
rect 513994 139218 514026 139454
rect 514262 139218 514346 139454
rect 514582 139218 514614 139454
rect 513994 139134 514614 139218
rect 513994 138898 514026 139134
rect 514262 138898 514346 139134
rect 514582 138898 514614 139134
rect 513994 102454 514614 138898
rect 513994 102218 514026 102454
rect 514262 102218 514346 102454
rect 514582 102218 514614 102454
rect 513994 102134 514614 102218
rect 513994 101898 514026 102134
rect 514262 101898 514346 102134
rect 514582 101898 514614 102134
rect 513994 65454 514614 101898
rect 513994 65218 514026 65454
rect 514262 65218 514346 65454
rect 514582 65218 514614 65454
rect 513994 65134 514614 65218
rect 513994 64898 514026 65134
rect 514262 64898 514346 65134
rect 514582 64898 514614 65134
rect 513994 28454 514614 64898
rect 513994 28218 514026 28454
rect 514262 28218 514346 28454
rect 514582 28218 514614 28454
rect 513994 28134 514614 28218
rect 513994 27898 514026 28134
rect 514262 27898 514346 28134
rect 514582 27898 514614 28134
rect 513994 -1306 514614 27898
rect 513994 -1542 514026 -1306
rect 514262 -1542 514346 -1306
rect 514582 -1542 514614 -1306
rect 513994 -1626 514614 -1542
rect 513994 -1862 514026 -1626
rect 514262 -1862 514346 -1626
rect 514582 -1862 514614 -1626
rect 513994 -7654 514614 -1862
rect 517714 704838 518334 711590
rect 517714 704602 517746 704838
rect 517982 704602 518066 704838
rect 518302 704602 518334 704838
rect 517714 704518 518334 704602
rect 517714 704282 517746 704518
rect 517982 704282 518066 704518
rect 518302 704282 518334 704518
rect 517714 698174 518334 704282
rect 517714 697938 517746 698174
rect 517982 697938 518066 698174
rect 518302 697938 518334 698174
rect 517714 697854 518334 697938
rect 517714 697618 517746 697854
rect 517982 697618 518066 697854
rect 518302 697618 518334 697854
rect 517714 661174 518334 697618
rect 517714 660938 517746 661174
rect 517982 660938 518066 661174
rect 518302 660938 518334 661174
rect 517714 660854 518334 660938
rect 517714 660618 517746 660854
rect 517982 660618 518066 660854
rect 518302 660618 518334 660854
rect 517714 624174 518334 660618
rect 517714 623938 517746 624174
rect 517982 623938 518066 624174
rect 518302 623938 518334 624174
rect 517714 623854 518334 623938
rect 517714 623618 517746 623854
rect 517982 623618 518066 623854
rect 518302 623618 518334 623854
rect 517714 587174 518334 623618
rect 517714 586938 517746 587174
rect 517982 586938 518066 587174
rect 518302 586938 518334 587174
rect 517714 586854 518334 586938
rect 517714 586618 517746 586854
rect 517982 586618 518066 586854
rect 518302 586618 518334 586854
rect 517714 550174 518334 586618
rect 517714 549938 517746 550174
rect 517982 549938 518066 550174
rect 518302 549938 518334 550174
rect 517714 549854 518334 549938
rect 517714 549618 517746 549854
rect 517982 549618 518066 549854
rect 518302 549618 518334 549854
rect 517714 513174 518334 549618
rect 517714 512938 517746 513174
rect 517982 512938 518066 513174
rect 518302 512938 518334 513174
rect 517714 512854 518334 512938
rect 517714 512618 517746 512854
rect 517982 512618 518066 512854
rect 518302 512618 518334 512854
rect 517714 476174 518334 512618
rect 517714 475938 517746 476174
rect 517982 475938 518066 476174
rect 518302 475938 518334 476174
rect 517714 475854 518334 475938
rect 517714 475618 517746 475854
rect 517982 475618 518066 475854
rect 518302 475618 518334 475854
rect 517714 439174 518334 475618
rect 517714 438938 517746 439174
rect 517982 438938 518066 439174
rect 518302 438938 518334 439174
rect 517714 438854 518334 438938
rect 517714 438618 517746 438854
rect 517982 438618 518066 438854
rect 518302 438618 518334 438854
rect 517714 402174 518334 438618
rect 517714 401938 517746 402174
rect 517982 401938 518066 402174
rect 518302 401938 518334 402174
rect 517714 401854 518334 401938
rect 517714 401618 517746 401854
rect 517982 401618 518066 401854
rect 518302 401618 518334 401854
rect 517714 365174 518334 401618
rect 517714 364938 517746 365174
rect 517982 364938 518066 365174
rect 518302 364938 518334 365174
rect 517714 364854 518334 364938
rect 517714 364618 517746 364854
rect 517982 364618 518066 364854
rect 518302 364618 518334 364854
rect 517714 328174 518334 364618
rect 517714 327938 517746 328174
rect 517982 327938 518066 328174
rect 518302 327938 518334 328174
rect 517714 327854 518334 327938
rect 517714 327618 517746 327854
rect 517982 327618 518066 327854
rect 518302 327618 518334 327854
rect 517714 291174 518334 327618
rect 517714 290938 517746 291174
rect 517982 290938 518066 291174
rect 518302 290938 518334 291174
rect 517714 290854 518334 290938
rect 517714 290618 517746 290854
rect 517982 290618 518066 290854
rect 518302 290618 518334 290854
rect 517714 254174 518334 290618
rect 517714 253938 517746 254174
rect 517982 253938 518066 254174
rect 518302 253938 518334 254174
rect 517714 253854 518334 253938
rect 517714 253618 517746 253854
rect 517982 253618 518066 253854
rect 518302 253618 518334 253854
rect 517714 217174 518334 253618
rect 517714 216938 517746 217174
rect 517982 216938 518066 217174
rect 518302 216938 518334 217174
rect 517714 216854 518334 216938
rect 517714 216618 517746 216854
rect 517982 216618 518066 216854
rect 518302 216618 518334 216854
rect 517714 180174 518334 216618
rect 517714 179938 517746 180174
rect 517982 179938 518066 180174
rect 518302 179938 518334 180174
rect 517714 179854 518334 179938
rect 517714 179618 517746 179854
rect 517982 179618 518066 179854
rect 518302 179618 518334 179854
rect 517714 143174 518334 179618
rect 517714 142938 517746 143174
rect 517982 142938 518066 143174
rect 518302 142938 518334 143174
rect 517714 142854 518334 142938
rect 517714 142618 517746 142854
rect 517982 142618 518066 142854
rect 518302 142618 518334 142854
rect 517714 106174 518334 142618
rect 517714 105938 517746 106174
rect 517982 105938 518066 106174
rect 518302 105938 518334 106174
rect 517714 105854 518334 105938
rect 517714 105618 517746 105854
rect 517982 105618 518066 105854
rect 518302 105618 518334 105854
rect 517714 69174 518334 105618
rect 517714 68938 517746 69174
rect 517982 68938 518066 69174
rect 518302 68938 518334 69174
rect 517714 68854 518334 68938
rect 517714 68618 517746 68854
rect 517982 68618 518066 68854
rect 518302 68618 518334 68854
rect 517714 32174 518334 68618
rect 517714 31938 517746 32174
rect 517982 31938 518066 32174
rect 518302 31938 518334 32174
rect 517714 31854 518334 31938
rect 517714 31618 517746 31854
rect 517982 31618 518066 31854
rect 518302 31618 518334 31854
rect 517714 -346 518334 31618
rect 517714 -582 517746 -346
rect 517982 -582 518066 -346
rect 518302 -582 518334 -346
rect 517714 -666 518334 -582
rect 517714 -902 517746 -666
rect 517982 -902 518066 -666
rect 518302 -902 518334 -666
rect 517714 -7654 518334 -902
rect 541994 705798 542614 711590
rect 541994 705562 542026 705798
rect 542262 705562 542346 705798
rect 542582 705562 542614 705798
rect 541994 705478 542614 705562
rect 541994 705242 542026 705478
rect 542262 705242 542346 705478
rect 542582 705242 542614 705478
rect 541994 694454 542614 705242
rect 541994 694218 542026 694454
rect 542262 694218 542346 694454
rect 542582 694218 542614 694454
rect 541994 694134 542614 694218
rect 541994 693898 542026 694134
rect 542262 693898 542346 694134
rect 542582 693898 542614 694134
rect 541994 657454 542614 693898
rect 541994 657218 542026 657454
rect 542262 657218 542346 657454
rect 542582 657218 542614 657454
rect 541994 657134 542614 657218
rect 541994 656898 542026 657134
rect 542262 656898 542346 657134
rect 542582 656898 542614 657134
rect 541994 620454 542614 656898
rect 541994 620218 542026 620454
rect 542262 620218 542346 620454
rect 542582 620218 542614 620454
rect 541994 620134 542614 620218
rect 541994 619898 542026 620134
rect 542262 619898 542346 620134
rect 542582 619898 542614 620134
rect 541994 583454 542614 619898
rect 541994 583218 542026 583454
rect 542262 583218 542346 583454
rect 542582 583218 542614 583454
rect 541994 583134 542614 583218
rect 541994 582898 542026 583134
rect 542262 582898 542346 583134
rect 542582 582898 542614 583134
rect 541994 546454 542614 582898
rect 541994 546218 542026 546454
rect 542262 546218 542346 546454
rect 542582 546218 542614 546454
rect 541994 546134 542614 546218
rect 541994 545898 542026 546134
rect 542262 545898 542346 546134
rect 542582 545898 542614 546134
rect 541994 509454 542614 545898
rect 541994 509218 542026 509454
rect 542262 509218 542346 509454
rect 542582 509218 542614 509454
rect 541994 509134 542614 509218
rect 541994 508898 542026 509134
rect 542262 508898 542346 509134
rect 542582 508898 542614 509134
rect 541994 472454 542614 508898
rect 541994 472218 542026 472454
rect 542262 472218 542346 472454
rect 542582 472218 542614 472454
rect 541994 472134 542614 472218
rect 541994 471898 542026 472134
rect 542262 471898 542346 472134
rect 542582 471898 542614 472134
rect 541994 435454 542614 471898
rect 541994 435218 542026 435454
rect 542262 435218 542346 435454
rect 542582 435218 542614 435454
rect 541994 435134 542614 435218
rect 541994 434898 542026 435134
rect 542262 434898 542346 435134
rect 542582 434898 542614 435134
rect 541994 398454 542614 434898
rect 541994 398218 542026 398454
rect 542262 398218 542346 398454
rect 542582 398218 542614 398454
rect 541994 398134 542614 398218
rect 541994 397898 542026 398134
rect 542262 397898 542346 398134
rect 542582 397898 542614 398134
rect 541994 361454 542614 397898
rect 541994 361218 542026 361454
rect 542262 361218 542346 361454
rect 542582 361218 542614 361454
rect 541994 361134 542614 361218
rect 541994 360898 542026 361134
rect 542262 360898 542346 361134
rect 542582 360898 542614 361134
rect 541994 324454 542614 360898
rect 541994 324218 542026 324454
rect 542262 324218 542346 324454
rect 542582 324218 542614 324454
rect 541994 324134 542614 324218
rect 541994 323898 542026 324134
rect 542262 323898 542346 324134
rect 542582 323898 542614 324134
rect 541994 287454 542614 323898
rect 541994 287218 542026 287454
rect 542262 287218 542346 287454
rect 542582 287218 542614 287454
rect 541994 287134 542614 287218
rect 541994 286898 542026 287134
rect 542262 286898 542346 287134
rect 542582 286898 542614 287134
rect 541994 250454 542614 286898
rect 541994 250218 542026 250454
rect 542262 250218 542346 250454
rect 542582 250218 542614 250454
rect 541994 250134 542614 250218
rect 541994 249898 542026 250134
rect 542262 249898 542346 250134
rect 542582 249898 542614 250134
rect 541994 213454 542614 249898
rect 541994 213218 542026 213454
rect 542262 213218 542346 213454
rect 542582 213218 542614 213454
rect 541994 213134 542614 213218
rect 541994 212898 542026 213134
rect 542262 212898 542346 213134
rect 542582 212898 542614 213134
rect 541994 176454 542614 212898
rect 541994 176218 542026 176454
rect 542262 176218 542346 176454
rect 542582 176218 542614 176454
rect 541994 176134 542614 176218
rect 541994 175898 542026 176134
rect 542262 175898 542346 176134
rect 542582 175898 542614 176134
rect 541994 139454 542614 175898
rect 541994 139218 542026 139454
rect 542262 139218 542346 139454
rect 542582 139218 542614 139454
rect 541994 139134 542614 139218
rect 541994 138898 542026 139134
rect 542262 138898 542346 139134
rect 542582 138898 542614 139134
rect 541994 102454 542614 138898
rect 541994 102218 542026 102454
rect 542262 102218 542346 102454
rect 542582 102218 542614 102454
rect 541994 102134 542614 102218
rect 541994 101898 542026 102134
rect 542262 101898 542346 102134
rect 542582 101898 542614 102134
rect 541994 65454 542614 101898
rect 541994 65218 542026 65454
rect 542262 65218 542346 65454
rect 542582 65218 542614 65454
rect 541994 65134 542614 65218
rect 541994 64898 542026 65134
rect 542262 64898 542346 65134
rect 542582 64898 542614 65134
rect 541994 28454 542614 64898
rect 541994 28218 542026 28454
rect 542262 28218 542346 28454
rect 542582 28218 542614 28454
rect 541994 28134 542614 28218
rect 541994 27898 542026 28134
rect 542262 27898 542346 28134
rect 542582 27898 542614 28134
rect 541994 -1306 542614 27898
rect 541994 -1542 542026 -1306
rect 542262 -1542 542346 -1306
rect 542582 -1542 542614 -1306
rect 541994 -1626 542614 -1542
rect 541994 -1862 542026 -1626
rect 542262 -1862 542346 -1626
rect 542582 -1862 542614 -1626
rect 541994 -7654 542614 -1862
rect 545714 704838 546334 711590
rect 545714 704602 545746 704838
rect 545982 704602 546066 704838
rect 546302 704602 546334 704838
rect 545714 704518 546334 704602
rect 545714 704282 545746 704518
rect 545982 704282 546066 704518
rect 546302 704282 546334 704518
rect 545714 698174 546334 704282
rect 545714 697938 545746 698174
rect 545982 697938 546066 698174
rect 546302 697938 546334 698174
rect 545714 697854 546334 697938
rect 545714 697618 545746 697854
rect 545982 697618 546066 697854
rect 546302 697618 546334 697854
rect 545714 661174 546334 697618
rect 545714 660938 545746 661174
rect 545982 660938 546066 661174
rect 546302 660938 546334 661174
rect 545714 660854 546334 660938
rect 545714 660618 545746 660854
rect 545982 660618 546066 660854
rect 546302 660618 546334 660854
rect 545714 624174 546334 660618
rect 545714 623938 545746 624174
rect 545982 623938 546066 624174
rect 546302 623938 546334 624174
rect 545714 623854 546334 623938
rect 545714 623618 545746 623854
rect 545982 623618 546066 623854
rect 546302 623618 546334 623854
rect 545714 587174 546334 623618
rect 545714 586938 545746 587174
rect 545982 586938 546066 587174
rect 546302 586938 546334 587174
rect 545714 586854 546334 586938
rect 545714 586618 545746 586854
rect 545982 586618 546066 586854
rect 546302 586618 546334 586854
rect 545714 550174 546334 586618
rect 545714 549938 545746 550174
rect 545982 549938 546066 550174
rect 546302 549938 546334 550174
rect 545714 549854 546334 549938
rect 545714 549618 545746 549854
rect 545982 549618 546066 549854
rect 546302 549618 546334 549854
rect 545714 513174 546334 549618
rect 545714 512938 545746 513174
rect 545982 512938 546066 513174
rect 546302 512938 546334 513174
rect 545714 512854 546334 512938
rect 545714 512618 545746 512854
rect 545982 512618 546066 512854
rect 546302 512618 546334 512854
rect 545714 476174 546334 512618
rect 545714 475938 545746 476174
rect 545982 475938 546066 476174
rect 546302 475938 546334 476174
rect 545714 475854 546334 475938
rect 545714 475618 545746 475854
rect 545982 475618 546066 475854
rect 546302 475618 546334 475854
rect 545714 439174 546334 475618
rect 545714 438938 545746 439174
rect 545982 438938 546066 439174
rect 546302 438938 546334 439174
rect 545714 438854 546334 438938
rect 545714 438618 545746 438854
rect 545982 438618 546066 438854
rect 546302 438618 546334 438854
rect 545714 402174 546334 438618
rect 545714 401938 545746 402174
rect 545982 401938 546066 402174
rect 546302 401938 546334 402174
rect 545714 401854 546334 401938
rect 545714 401618 545746 401854
rect 545982 401618 546066 401854
rect 546302 401618 546334 401854
rect 545714 365174 546334 401618
rect 545714 364938 545746 365174
rect 545982 364938 546066 365174
rect 546302 364938 546334 365174
rect 545714 364854 546334 364938
rect 545714 364618 545746 364854
rect 545982 364618 546066 364854
rect 546302 364618 546334 364854
rect 545714 328174 546334 364618
rect 545714 327938 545746 328174
rect 545982 327938 546066 328174
rect 546302 327938 546334 328174
rect 545714 327854 546334 327938
rect 545714 327618 545746 327854
rect 545982 327618 546066 327854
rect 546302 327618 546334 327854
rect 545714 291174 546334 327618
rect 545714 290938 545746 291174
rect 545982 290938 546066 291174
rect 546302 290938 546334 291174
rect 545714 290854 546334 290938
rect 545714 290618 545746 290854
rect 545982 290618 546066 290854
rect 546302 290618 546334 290854
rect 545714 254174 546334 290618
rect 545714 253938 545746 254174
rect 545982 253938 546066 254174
rect 546302 253938 546334 254174
rect 545714 253854 546334 253938
rect 545714 253618 545746 253854
rect 545982 253618 546066 253854
rect 546302 253618 546334 253854
rect 545714 217174 546334 253618
rect 545714 216938 545746 217174
rect 545982 216938 546066 217174
rect 546302 216938 546334 217174
rect 545714 216854 546334 216938
rect 545714 216618 545746 216854
rect 545982 216618 546066 216854
rect 546302 216618 546334 216854
rect 545714 180174 546334 216618
rect 545714 179938 545746 180174
rect 545982 179938 546066 180174
rect 546302 179938 546334 180174
rect 545714 179854 546334 179938
rect 545714 179618 545746 179854
rect 545982 179618 546066 179854
rect 546302 179618 546334 179854
rect 545714 143174 546334 179618
rect 545714 142938 545746 143174
rect 545982 142938 546066 143174
rect 546302 142938 546334 143174
rect 545714 142854 546334 142938
rect 545714 142618 545746 142854
rect 545982 142618 546066 142854
rect 546302 142618 546334 142854
rect 545714 106174 546334 142618
rect 545714 105938 545746 106174
rect 545982 105938 546066 106174
rect 546302 105938 546334 106174
rect 545714 105854 546334 105938
rect 545714 105618 545746 105854
rect 545982 105618 546066 105854
rect 546302 105618 546334 105854
rect 545714 69174 546334 105618
rect 545714 68938 545746 69174
rect 545982 68938 546066 69174
rect 546302 68938 546334 69174
rect 545714 68854 546334 68938
rect 545714 68618 545746 68854
rect 545982 68618 546066 68854
rect 546302 68618 546334 68854
rect 545714 32174 546334 68618
rect 545714 31938 545746 32174
rect 545982 31938 546066 32174
rect 546302 31938 546334 32174
rect 545714 31854 546334 31938
rect 545714 31618 545746 31854
rect 545982 31618 546066 31854
rect 546302 31618 546334 31854
rect 545714 -346 546334 31618
rect 545714 -582 545746 -346
rect 545982 -582 546066 -346
rect 546302 -582 546334 -346
rect 545714 -666 546334 -582
rect 545714 -902 545746 -666
rect 545982 -902 546066 -666
rect 546302 -902 546334 -666
rect 545714 -7654 546334 -902
rect 569994 705798 570614 711590
rect 569994 705562 570026 705798
rect 570262 705562 570346 705798
rect 570582 705562 570614 705798
rect 569994 705478 570614 705562
rect 569994 705242 570026 705478
rect 570262 705242 570346 705478
rect 570582 705242 570614 705478
rect 569994 694454 570614 705242
rect 569994 694218 570026 694454
rect 570262 694218 570346 694454
rect 570582 694218 570614 694454
rect 569994 694134 570614 694218
rect 569994 693898 570026 694134
rect 570262 693898 570346 694134
rect 570582 693898 570614 694134
rect 569994 657454 570614 693898
rect 569994 657218 570026 657454
rect 570262 657218 570346 657454
rect 570582 657218 570614 657454
rect 569994 657134 570614 657218
rect 569994 656898 570026 657134
rect 570262 656898 570346 657134
rect 570582 656898 570614 657134
rect 569994 620454 570614 656898
rect 569994 620218 570026 620454
rect 570262 620218 570346 620454
rect 570582 620218 570614 620454
rect 569994 620134 570614 620218
rect 569994 619898 570026 620134
rect 570262 619898 570346 620134
rect 570582 619898 570614 620134
rect 569994 583454 570614 619898
rect 569994 583218 570026 583454
rect 570262 583218 570346 583454
rect 570582 583218 570614 583454
rect 569994 583134 570614 583218
rect 569994 582898 570026 583134
rect 570262 582898 570346 583134
rect 570582 582898 570614 583134
rect 569994 546454 570614 582898
rect 569994 546218 570026 546454
rect 570262 546218 570346 546454
rect 570582 546218 570614 546454
rect 569994 546134 570614 546218
rect 569994 545898 570026 546134
rect 570262 545898 570346 546134
rect 570582 545898 570614 546134
rect 569994 509454 570614 545898
rect 569994 509218 570026 509454
rect 570262 509218 570346 509454
rect 570582 509218 570614 509454
rect 569994 509134 570614 509218
rect 569994 508898 570026 509134
rect 570262 508898 570346 509134
rect 570582 508898 570614 509134
rect 569994 472454 570614 508898
rect 569994 472218 570026 472454
rect 570262 472218 570346 472454
rect 570582 472218 570614 472454
rect 569994 472134 570614 472218
rect 569994 471898 570026 472134
rect 570262 471898 570346 472134
rect 570582 471898 570614 472134
rect 569994 435454 570614 471898
rect 569994 435218 570026 435454
rect 570262 435218 570346 435454
rect 570582 435218 570614 435454
rect 569994 435134 570614 435218
rect 569994 434898 570026 435134
rect 570262 434898 570346 435134
rect 570582 434898 570614 435134
rect 569994 398454 570614 434898
rect 569994 398218 570026 398454
rect 570262 398218 570346 398454
rect 570582 398218 570614 398454
rect 569994 398134 570614 398218
rect 569994 397898 570026 398134
rect 570262 397898 570346 398134
rect 570582 397898 570614 398134
rect 569994 361454 570614 397898
rect 569994 361218 570026 361454
rect 570262 361218 570346 361454
rect 570582 361218 570614 361454
rect 569994 361134 570614 361218
rect 569994 360898 570026 361134
rect 570262 360898 570346 361134
rect 570582 360898 570614 361134
rect 569994 324454 570614 360898
rect 569994 324218 570026 324454
rect 570262 324218 570346 324454
rect 570582 324218 570614 324454
rect 569994 324134 570614 324218
rect 569994 323898 570026 324134
rect 570262 323898 570346 324134
rect 570582 323898 570614 324134
rect 569994 287454 570614 323898
rect 569994 287218 570026 287454
rect 570262 287218 570346 287454
rect 570582 287218 570614 287454
rect 569994 287134 570614 287218
rect 569994 286898 570026 287134
rect 570262 286898 570346 287134
rect 570582 286898 570614 287134
rect 569994 250454 570614 286898
rect 569994 250218 570026 250454
rect 570262 250218 570346 250454
rect 570582 250218 570614 250454
rect 569994 250134 570614 250218
rect 569994 249898 570026 250134
rect 570262 249898 570346 250134
rect 570582 249898 570614 250134
rect 569994 213454 570614 249898
rect 569994 213218 570026 213454
rect 570262 213218 570346 213454
rect 570582 213218 570614 213454
rect 569994 213134 570614 213218
rect 569994 212898 570026 213134
rect 570262 212898 570346 213134
rect 570582 212898 570614 213134
rect 569994 176454 570614 212898
rect 569994 176218 570026 176454
rect 570262 176218 570346 176454
rect 570582 176218 570614 176454
rect 569994 176134 570614 176218
rect 569994 175898 570026 176134
rect 570262 175898 570346 176134
rect 570582 175898 570614 176134
rect 569994 139454 570614 175898
rect 569994 139218 570026 139454
rect 570262 139218 570346 139454
rect 570582 139218 570614 139454
rect 569994 139134 570614 139218
rect 569994 138898 570026 139134
rect 570262 138898 570346 139134
rect 570582 138898 570614 139134
rect 569994 102454 570614 138898
rect 569994 102218 570026 102454
rect 570262 102218 570346 102454
rect 570582 102218 570614 102454
rect 569994 102134 570614 102218
rect 569994 101898 570026 102134
rect 570262 101898 570346 102134
rect 570582 101898 570614 102134
rect 569994 65454 570614 101898
rect 569994 65218 570026 65454
rect 570262 65218 570346 65454
rect 570582 65218 570614 65454
rect 569994 65134 570614 65218
rect 569994 64898 570026 65134
rect 570262 64898 570346 65134
rect 570582 64898 570614 65134
rect 569994 28454 570614 64898
rect 569994 28218 570026 28454
rect 570262 28218 570346 28454
rect 570582 28218 570614 28454
rect 569994 28134 570614 28218
rect 569994 27898 570026 28134
rect 570262 27898 570346 28134
rect 570582 27898 570614 28134
rect 569994 -1306 570614 27898
rect 569994 -1542 570026 -1306
rect 570262 -1542 570346 -1306
rect 570582 -1542 570614 -1306
rect 569994 -1626 570614 -1542
rect 569994 -1862 570026 -1626
rect 570262 -1862 570346 -1626
rect 570582 -1862 570614 -1626
rect 569994 -7654 570614 -1862
rect 573714 704838 574334 711590
rect 592030 711558 592650 711590
rect 592030 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect 592030 711238 592650 711322
rect 592030 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect 591070 710598 591690 710630
rect 591070 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect 591070 710278 591690 710362
rect 591070 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect 590110 709638 590730 709670
rect 590110 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect 590110 709318 590730 709402
rect 590110 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect 589150 708678 589770 708710
rect 589150 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect 589150 708358 589770 708442
rect 589150 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect 588190 707718 588810 707750
rect 588190 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect 588190 707398 588810 707482
rect 588190 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect 587230 706758 587850 706790
rect 587230 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect 587230 706438 587850 706522
rect 587230 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect 586270 705798 586890 705830
rect 586270 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect 586270 705478 586890 705562
rect 586270 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect 573714 704602 573746 704838
rect 573982 704602 574066 704838
rect 574302 704602 574334 704838
rect 573714 704518 574334 704602
rect 573714 704282 573746 704518
rect 573982 704282 574066 704518
rect 574302 704282 574334 704518
rect 573714 698174 574334 704282
rect 573714 697938 573746 698174
rect 573982 697938 574066 698174
rect 574302 697938 574334 698174
rect 573714 697854 574334 697938
rect 573714 697618 573746 697854
rect 573982 697618 574066 697854
rect 574302 697618 574334 697854
rect 573714 661174 574334 697618
rect 573714 660938 573746 661174
rect 573982 660938 574066 661174
rect 574302 660938 574334 661174
rect 573714 660854 574334 660938
rect 573714 660618 573746 660854
rect 573982 660618 574066 660854
rect 574302 660618 574334 660854
rect 573714 624174 574334 660618
rect 573714 623938 573746 624174
rect 573982 623938 574066 624174
rect 574302 623938 574334 624174
rect 573714 623854 574334 623938
rect 573714 623618 573746 623854
rect 573982 623618 574066 623854
rect 574302 623618 574334 623854
rect 573714 587174 574334 623618
rect 573714 586938 573746 587174
rect 573982 586938 574066 587174
rect 574302 586938 574334 587174
rect 573714 586854 574334 586938
rect 573714 586618 573746 586854
rect 573982 586618 574066 586854
rect 574302 586618 574334 586854
rect 573714 550174 574334 586618
rect 573714 549938 573746 550174
rect 573982 549938 574066 550174
rect 574302 549938 574334 550174
rect 573714 549854 574334 549938
rect 573714 549618 573746 549854
rect 573982 549618 574066 549854
rect 574302 549618 574334 549854
rect 573714 513174 574334 549618
rect 573714 512938 573746 513174
rect 573982 512938 574066 513174
rect 574302 512938 574334 513174
rect 573714 512854 574334 512938
rect 573714 512618 573746 512854
rect 573982 512618 574066 512854
rect 574302 512618 574334 512854
rect 573714 476174 574334 512618
rect 573714 475938 573746 476174
rect 573982 475938 574066 476174
rect 574302 475938 574334 476174
rect 573714 475854 574334 475938
rect 573714 475618 573746 475854
rect 573982 475618 574066 475854
rect 574302 475618 574334 475854
rect 573714 439174 574334 475618
rect 573714 438938 573746 439174
rect 573982 438938 574066 439174
rect 574302 438938 574334 439174
rect 573714 438854 574334 438938
rect 573714 438618 573746 438854
rect 573982 438618 574066 438854
rect 574302 438618 574334 438854
rect 573714 402174 574334 438618
rect 573714 401938 573746 402174
rect 573982 401938 574066 402174
rect 574302 401938 574334 402174
rect 573714 401854 574334 401938
rect 573714 401618 573746 401854
rect 573982 401618 574066 401854
rect 574302 401618 574334 401854
rect 573714 365174 574334 401618
rect 573714 364938 573746 365174
rect 573982 364938 574066 365174
rect 574302 364938 574334 365174
rect 573714 364854 574334 364938
rect 573714 364618 573746 364854
rect 573982 364618 574066 364854
rect 574302 364618 574334 364854
rect 573714 328174 574334 364618
rect 573714 327938 573746 328174
rect 573982 327938 574066 328174
rect 574302 327938 574334 328174
rect 573714 327854 574334 327938
rect 573714 327618 573746 327854
rect 573982 327618 574066 327854
rect 574302 327618 574334 327854
rect 573714 291174 574334 327618
rect 573714 290938 573746 291174
rect 573982 290938 574066 291174
rect 574302 290938 574334 291174
rect 573714 290854 574334 290938
rect 573714 290618 573746 290854
rect 573982 290618 574066 290854
rect 574302 290618 574334 290854
rect 573714 254174 574334 290618
rect 573714 253938 573746 254174
rect 573982 253938 574066 254174
rect 574302 253938 574334 254174
rect 573714 253854 574334 253938
rect 573714 253618 573746 253854
rect 573982 253618 574066 253854
rect 574302 253618 574334 253854
rect 573714 217174 574334 253618
rect 573714 216938 573746 217174
rect 573982 216938 574066 217174
rect 574302 216938 574334 217174
rect 573714 216854 574334 216938
rect 573714 216618 573746 216854
rect 573982 216618 574066 216854
rect 574302 216618 574334 216854
rect 573714 180174 574334 216618
rect 573714 179938 573746 180174
rect 573982 179938 574066 180174
rect 574302 179938 574334 180174
rect 573714 179854 574334 179938
rect 573714 179618 573746 179854
rect 573982 179618 574066 179854
rect 574302 179618 574334 179854
rect 573714 143174 574334 179618
rect 573714 142938 573746 143174
rect 573982 142938 574066 143174
rect 574302 142938 574334 143174
rect 573714 142854 574334 142938
rect 573714 142618 573746 142854
rect 573982 142618 574066 142854
rect 574302 142618 574334 142854
rect 573714 106174 574334 142618
rect 573714 105938 573746 106174
rect 573982 105938 574066 106174
rect 574302 105938 574334 106174
rect 573714 105854 574334 105938
rect 573714 105618 573746 105854
rect 573982 105618 574066 105854
rect 574302 105618 574334 105854
rect 573714 69174 574334 105618
rect 573714 68938 573746 69174
rect 573982 68938 574066 69174
rect 574302 68938 574334 69174
rect 573714 68854 574334 68938
rect 573714 68618 573746 68854
rect 573982 68618 574066 68854
rect 574302 68618 574334 68854
rect 573714 32174 574334 68618
rect 573714 31938 573746 32174
rect 573982 31938 574066 32174
rect 574302 31938 574334 32174
rect 573714 31854 574334 31938
rect 573714 31618 573746 31854
rect 573982 31618 574066 31854
rect 574302 31618 574334 31854
rect 573714 -346 574334 31618
rect 573714 -582 573746 -346
rect 573982 -582 574066 -346
rect 574302 -582 574334 -346
rect 573714 -666 574334 -582
rect 573714 -902 573746 -666
rect 573982 -902 574066 -666
rect 574302 -902 574334 -666
rect 573714 -7654 574334 -902
rect 585310 704838 585930 704870
rect 585310 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect 585310 704518 585930 704602
rect 585310 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect 585310 698174 585930 704282
rect 585310 697938 585342 698174
rect 585578 697938 585662 698174
rect 585898 697938 585930 698174
rect 585310 697854 585930 697938
rect 585310 697618 585342 697854
rect 585578 697618 585662 697854
rect 585898 697618 585930 697854
rect 585310 661174 585930 697618
rect 585310 660938 585342 661174
rect 585578 660938 585662 661174
rect 585898 660938 585930 661174
rect 585310 660854 585930 660938
rect 585310 660618 585342 660854
rect 585578 660618 585662 660854
rect 585898 660618 585930 660854
rect 585310 624174 585930 660618
rect 585310 623938 585342 624174
rect 585578 623938 585662 624174
rect 585898 623938 585930 624174
rect 585310 623854 585930 623938
rect 585310 623618 585342 623854
rect 585578 623618 585662 623854
rect 585898 623618 585930 623854
rect 585310 587174 585930 623618
rect 585310 586938 585342 587174
rect 585578 586938 585662 587174
rect 585898 586938 585930 587174
rect 585310 586854 585930 586938
rect 585310 586618 585342 586854
rect 585578 586618 585662 586854
rect 585898 586618 585930 586854
rect 585310 550174 585930 586618
rect 585310 549938 585342 550174
rect 585578 549938 585662 550174
rect 585898 549938 585930 550174
rect 585310 549854 585930 549938
rect 585310 549618 585342 549854
rect 585578 549618 585662 549854
rect 585898 549618 585930 549854
rect 585310 513174 585930 549618
rect 585310 512938 585342 513174
rect 585578 512938 585662 513174
rect 585898 512938 585930 513174
rect 585310 512854 585930 512938
rect 585310 512618 585342 512854
rect 585578 512618 585662 512854
rect 585898 512618 585930 512854
rect 585310 476174 585930 512618
rect 585310 475938 585342 476174
rect 585578 475938 585662 476174
rect 585898 475938 585930 476174
rect 585310 475854 585930 475938
rect 585310 475618 585342 475854
rect 585578 475618 585662 475854
rect 585898 475618 585930 475854
rect 585310 439174 585930 475618
rect 585310 438938 585342 439174
rect 585578 438938 585662 439174
rect 585898 438938 585930 439174
rect 585310 438854 585930 438938
rect 585310 438618 585342 438854
rect 585578 438618 585662 438854
rect 585898 438618 585930 438854
rect 585310 402174 585930 438618
rect 585310 401938 585342 402174
rect 585578 401938 585662 402174
rect 585898 401938 585930 402174
rect 585310 401854 585930 401938
rect 585310 401618 585342 401854
rect 585578 401618 585662 401854
rect 585898 401618 585930 401854
rect 585310 365174 585930 401618
rect 585310 364938 585342 365174
rect 585578 364938 585662 365174
rect 585898 364938 585930 365174
rect 585310 364854 585930 364938
rect 585310 364618 585342 364854
rect 585578 364618 585662 364854
rect 585898 364618 585930 364854
rect 585310 328174 585930 364618
rect 585310 327938 585342 328174
rect 585578 327938 585662 328174
rect 585898 327938 585930 328174
rect 585310 327854 585930 327938
rect 585310 327618 585342 327854
rect 585578 327618 585662 327854
rect 585898 327618 585930 327854
rect 585310 291174 585930 327618
rect 585310 290938 585342 291174
rect 585578 290938 585662 291174
rect 585898 290938 585930 291174
rect 585310 290854 585930 290938
rect 585310 290618 585342 290854
rect 585578 290618 585662 290854
rect 585898 290618 585930 290854
rect 585310 254174 585930 290618
rect 585310 253938 585342 254174
rect 585578 253938 585662 254174
rect 585898 253938 585930 254174
rect 585310 253854 585930 253938
rect 585310 253618 585342 253854
rect 585578 253618 585662 253854
rect 585898 253618 585930 253854
rect 585310 217174 585930 253618
rect 585310 216938 585342 217174
rect 585578 216938 585662 217174
rect 585898 216938 585930 217174
rect 585310 216854 585930 216938
rect 585310 216618 585342 216854
rect 585578 216618 585662 216854
rect 585898 216618 585930 216854
rect 585310 180174 585930 216618
rect 585310 179938 585342 180174
rect 585578 179938 585662 180174
rect 585898 179938 585930 180174
rect 585310 179854 585930 179938
rect 585310 179618 585342 179854
rect 585578 179618 585662 179854
rect 585898 179618 585930 179854
rect 585310 143174 585930 179618
rect 585310 142938 585342 143174
rect 585578 142938 585662 143174
rect 585898 142938 585930 143174
rect 585310 142854 585930 142938
rect 585310 142618 585342 142854
rect 585578 142618 585662 142854
rect 585898 142618 585930 142854
rect 585310 106174 585930 142618
rect 585310 105938 585342 106174
rect 585578 105938 585662 106174
rect 585898 105938 585930 106174
rect 585310 105854 585930 105938
rect 585310 105618 585342 105854
rect 585578 105618 585662 105854
rect 585898 105618 585930 105854
rect 585310 69174 585930 105618
rect 585310 68938 585342 69174
rect 585578 68938 585662 69174
rect 585898 68938 585930 69174
rect 585310 68854 585930 68938
rect 585310 68618 585342 68854
rect 585578 68618 585662 68854
rect 585898 68618 585930 68854
rect 585310 32174 585930 68618
rect 585310 31938 585342 32174
rect 585578 31938 585662 32174
rect 585898 31938 585930 32174
rect 585310 31854 585930 31938
rect 585310 31618 585342 31854
rect 585578 31618 585662 31854
rect 585898 31618 585930 31854
rect 585310 -346 585930 31618
rect 585310 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect 585310 -666 585930 -582
rect 585310 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect 585310 -934 585930 -902
rect 586270 694454 586890 705242
rect 586270 694218 586302 694454
rect 586538 694218 586622 694454
rect 586858 694218 586890 694454
rect 586270 694134 586890 694218
rect 586270 693898 586302 694134
rect 586538 693898 586622 694134
rect 586858 693898 586890 694134
rect 586270 657454 586890 693898
rect 586270 657218 586302 657454
rect 586538 657218 586622 657454
rect 586858 657218 586890 657454
rect 586270 657134 586890 657218
rect 586270 656898 586302 657134
rect 586538 656898 586622 657134
rect 586858 656898 586890 657134
rect 586270 620454 586890 656898
rect 586270 620218 586302 620454
rect 586538 620218 586622 620454
rect 586858 620218 586890 620454
rect 586270 620134 586890 620218
rect 586270 619898 586302 620134
rect 586538 619898 586622 620134
rect 586858 619898 586890 620134
rect 586270 583454 586890 619898
rect 586270 583218 586302 583454
rect 586538 583218 586622 583454
rect 586858 583218 586890 583454
rect 586270 583134 586890 583218
rect 586270 582898 586302 583134
rect 586538 582898 586622 583134
rect 586858 582898 586890 583134
rect 586270 546454 586890 582898
rect 586270 546218 586302 546454
rect 586538 546218 586622 546454
rect 586858 546218 586890 546454
rect 586270 546134 586890 546218
rect 586270 545898 586302 546134
rect 586538 545898 586622 546134
rect 586858 545898 586890 546134
rect 586270 509454 586890 545898
rect 586270 509218 586302 509454
rect 586538 509218 586622 509454
rect 586858 509218 586890 509454
rect 586270 509134 586890 509218
rect 586270 508898 586302 509134
rect 586538 508898 586622 509134
rect 586858 508898 586890 509134
rect 586270 472454 586890 508898
rect 586270 472218 586302 472454
rect 586538 472218 586622 472454
rect 586858 472218 586890 472454
rect 586270 472134 586890 472218
rect 586270 471898 586302 472134
rect 586538 471898 586622 472134
rect 586858 471898 586890 472134
rect 586270 435454 586890 471898
rect 586270 435218 586302 435454
rect 586538 435218 586622 435454
rect 586858 435218 586890 435454
rect 586270 435134 586890 435218
rect 586270 434898 586302 435134
rect 586538 434898 586622 435134
rect 586858 434898 586890 435134
rect 586270 398454 586890 434898
rect 586270 398218 586302 398454
rect 586538 398218 586622 398454
rect 586858 398218 586890 398454
rect 586270 398134 586890 398218
rect 586270 397898 586302 398134
rect 586538 397898 586622 398134
rect 586858 397898 586890 398134
rect 586270 361454 586890 397898
rect 586270 361218 586302 361454
rect 586538 361218 586622 361454
rect 586858 361218 586890 361454
rect 586270 361134 586890 361218
rect 586270 360898 586302 361134
rect 586538 360898 586622 361134
rect 586858 360898 586890 361134
rect 586270 324454 586890 360898
rect 586270 324218 586302 324454
rect 586538 324218 586622 324454
rect 586858 324218 586890 324454
rect 586270 324134 586890 324218
rect 586270 323898 586302 324134
rect 586538 323898 586622 324134
rect 586858 323898 586890 324134
rect 586270 287454 586890 323898
rect 586270 287218 586302 287454
rect 586538 287218 586622 287454
rect 586858 287218 586890 287454
rect 586270 287134 586890 287218
rect 586270 286898 586302 287134
rect 586538 286898 586622 287134
rect 586858 286898 586890 287134
rect 586270 250454 586890 286898
rect 586270 250218 586302 250454
rect 586538 250218 586622 250454
rect 586858 250218 586890 250454
rect 586270 250134 586890 250218
rect 586270 249898 586302 250134
rect 586538 249898 586622 250134
rect 586858 249898 586890 250134
rect 586270 213454 586890 249898
rect 586270 213218 586302 213454
rect 586538 213218 586622 213454
rect 586858 213218 586890 213454
rect 586270 213134 586890 213218
rect 586270 212898 586302 213134
rect 586538 212898 586622 213134
rect 586858 212898 586890 213134
rect 586270 176454 586890 212898
rect 586270 176218 586302 176454
rect 586538 176218 586622 176454
rect 586858 176218 586890 176454
rect 586270 176134 586890 176218
rect 586270 175898 586302 176134
rect 586538 175898 586622 176134
rect 586858 175898 586890 176134
rect 586270 139454 586890 175898
rect 586270 139218 586302 139454
rect 586538 139218 586622 139454
rect 586858 139218 586890 139454
rect 586270 139134 586890 139218
rect 586270 138898 586302 139134
rect 586538 138898 586622 139134
rect 586858 138898 586890 139134
rect 586270 102454 586890 138898
rect 586270 102218 586302 102454
rect 586538 102218 586622 102454
rect 586858 102218 586890 102454
rect 586270 102134 586890 102218
rect 586270 101898 586302 102134
rect 586538 101898 586622 102134
rect 586858 101898 586890 102134
rect 586270 65454 586890 101898
rect 586270 65218 586302 65454
rect 586538 65218 586622 65454
rect 586858 65218 586890 65454
rect 586270 65134 586890 65218
rect 586270 64898 586302 65134
rect 586538 64898 586622 65134
rect 586858 64898 586890 65134
rect 586270 28454 586890 64898
rect 586270 28218 586302 28454
rect 586538 28218 586622 28454
rect 586858 28218 586890 28454
rect 586270 28134 586890 28218
rect 586270 27898 586302 28134
rect 586538 27898 586622 28134
rect 586858 27898 586890 28134
rect 586270 -1306 586890 27898
rect 586270 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect 586270 -1626 586890 -1542
rect 586270 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect 586270 -1894 586890 -1862
rect 587230 -2266 587850 706202
rect 587230 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect 587230 -2586 587850 -2502
rect 587230 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect 587230 -2854 587850 -2822
rect 588190 -3226 588810 707162
rect 588190 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect 588190 -3546 588810 -3462
rect 588190 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect 588190 -3814 588810 -3782
rect 589150 -4186 589770 708122
rect 589150 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect 589150 -4506 589770 -4422
rect 589150 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect 589150 -4774 589770 -4742
rect 590110 -5146 590730 709082
rect 590110 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect 590110 -5466 590730 -5382
rect 590110 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect 590110 -5734 590730 -5702
rect 591070 -6106 591690 710042
rect 591070 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect 591070 -6426 591690 -6342
rect 591070 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect 591070 -6694 591690 -6662
rect 592030 -7066 592650 711002
rect 592030 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect 592030 -7386 592650 -7302
rect 592030 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect 592030 -7654 592650 -7622
<< via4 >>
rect -8694 711322 -8458 711558
rect -8374 711322 -8138 711558
rect -8694 711002 -8458 711238
rect -8374 711002 -8138 711238
rect -7734 710362 -7498 710598
rect -7414 710362 -7178 710598
rect -7734 710042 -7498 710278
rect -7414 710042 -7178 710278
rect -6774 709402 -6538 709638
rect -6454 709402 -6218 709638
rect -6774 709082 -6538 709318
rect -6454 709082 -6218 709318
rect -5814 708442 -5578 708678
rect -5494 708442 -5258 708678
rect -5814 708122 -5578 708358
rect -5494 708122 -5258 708358
rect -4854 707482 -4618 707718
rect -4534 707482 -4298 707718
rect -4854 707162 -4618 707398
rect -4534 707162 -4298 707398
rect -3894 706522 -3658 706758
rect -3574 706522 -3338 706758
rect -3894 706202 -3658 706438
rect -3574 706202 -3338 706438
rect -2934 705562 -2698 705798
rect -2614 705562 -2378 705798
rect -2934 705242 -2698 705478
rect -2614 705242 -2378 705478
rect 38026 705562 38262 705798
rect 38346 705562 38582 705798
rect 38026 705242 38262 705478
rect 38346 705242 38582 705478
rect -2934 694218 -2698 694454
rect -2614 694218 -2378 694454
rect -2934 693898 -2698 694134
rect -2614 693898 -2378 694134
rect -2934 657218 -2698 657454
rect -2614 657218 -2378 657454
rect -2934 656898 -2698 657134
rect -2614 656898 -2378 657134
rect -2934 620218 -2698 620454
rect -2614 620218 -2378 620454
rect -2934 619898 -2698 620134
rect -2614 619898 -2378 620134
rect -2934 583218 -2698 583454
rect -2614 583218 -2378 583454
rect -2934 582898 -2698 583134
rect -2614 582898 -2378 583134
rect -2934 546218 -2698 546454
rect -2614 546218 -2378 546454
rect -2934 545898 -2698 546134
rect -2614 545898 -2378 546134
rect -2934 509218 -2698 509454
rect -2614 509218 -2378 509454
rect -2934 508898 -2698 509134
rect -2614 508898 -2378 509134
rect -2934 472218 -2698 472454
rect -2614 472218 -2378 472454
rect -2934 471898 -2698 472134
rect -2614 471898 -2378 472134
rect -2934 435218 -2698 435454
rect -2614 435218 -2378 435454
rect -2934 434898 -2698 435134
rect -2614 434898 -2378 435134
rect -2934 398218 -2698 398454
rect -2614 398218 -2378 398454
rect -2934 397898 -2698 398134
rect -2614 397898 -2378 398134
rect -2934 361218 -2698 361454
rect -2614 361218 -2378 361454
rect -2934 360898 -2698 361134
rect -2614 360898 -2378 361134
rect -2934 324218 -2698 324454
rect -2614 324218 -2378 324454
rect -2934 323898 -2698 324134
rect -2614 323898 -2378 324134
rect -2934 287218 -2698 287454
rect -2614 287218 -2378 287454
rect -2934 286898 -2698 287134
rect -2614 286898 -2378 287134
rect -2934 250218 -2698 250454
rect -2614 250218 -2378 250454
rect -2934 249898 -2698 250134
rect -2614 249898 -2378 250134
rect -2934 213218 -2698 213454
rect -2614 213218 -2378 213454
rect -2934 212898 -2698 213134
rect -2614 212898 -2378 213134
rect -2934 176218 -2698 176454
rect -2614 176218 -2378 176454
rect -2934 175898 -2698 176134
rect -2614 175898 -2378 176134
rect -2934 139218 -2698 139454
rect -2614 139218 -2378 139454
rect -2934 138898 -2698 139134
rect -2614 138898 -2378 139134
rect -2934 102218 -2698 102454
rect -2614 102218 -2378 102454
rect -2934 101898 -2698 102134
rect -2614 101898 -2378 102134
rect -2934 65218 -2698 65454
rect -2614 65218 -2378 65454
rect -2934 64898 -2698 65134
rect -2614 64898 -2378 65134
rect -2934 28218 -2698 28454
rect -2614 28218 -2378 28454
rect -2934 27898 -2698 28134
rect -2614 27898 -2378 28134
rect -1974 704602 -1738 704838
rect -1654 704602 -1418 704838
rect -1974 704282 -1738 704518
rect -1654 704282 -1418 704518
rect -1974 697938 -1738 698174
rect -1654 697938 -1418 698174
rect -1974 697618 -1738 697854
rect -1654 697618 -1418 697854
rect -1974 660938 -1738 661174
rect -1654 660938 -1418 661174
rect -1974 660618 -1738 660854
rect -1654 660618 -1418 660854
rect -1974 623938 -1738 624174
rect -1654 623938 -1418 624174
rect -1974 623618 -1738 623854
rect -1654 623618 -1418 623854
rect 38026 694218 38262 694454
rect 38346 694218 38582 694454
rect 38026 693898 38262 694134
rect 38346 693898 38582 694134
rect 38026 657218 38262 657454
rect 38346 657218 38582 657454
rect 38026 656898 38262 657134
rect 38346 656898 38582 657134
rect 38026 620218 38262 620454
rect 38346 620218 38582 620454
rect 38026 619898 38262 620134
rect 38346 619898 38582 620134
rect -1974 586938 -1738 587174
rect -1654 586938 -1418 587174
rect -1974 586618 -1738 586854
rect -1654 586618 -1418 586854
rect -1974 549938 -1738 550174
rect -1654 549938 -1418 550174
rect -1974 549618 -1738 549854
rect -1654 549618 -1418 549854
rect -1974 512938 -1738 513174
rect -1654 512938 -1418 513174
rect -1974 512618 -1738 512854
rect -1654 512618 -1418 512854
rect -1974 475938 -1738 476174
rect -1654 475938 -1418 476174
rect -1974 475618 -1738 475854
rect -1654 475618 -1418 475854
rect -1974 438938 -1738 439174
rect -1654 438938 -1418 439174
rect -1974 438618 -1738 438854
rect -1654 438618 -1418 438854
rect -1974 401938 -1738 402174
rect -1654 401938 -1418 402174
rect -1974 401618 -1738 401854
rect -1654 401618 -1418 401854
rect -1974 364938 -1738 365174
rect -1654 364938 -1418 365174
rect -1974 364618 -1738 364854
rect -1654 364618 -1418 364854
rect -1974 327938 -1738 328174
rect -1654 327938 -1418 328174
rect -1974 327618 -1738 327854
rect -1654 327618 -1418 327854
rect -1974 290938 -1738 291174
rect -1654 290938 -1418 291174
rect -1974 290618 -1738 290854
rect -1654 290618 -1418 290854
rect -1974 253938 -1738 254174
rect -1654 253938 -1418 254174
rect -1974 253618 -1738 253854
rect -1654 253618 -1418 253854
rect -1974 216938 -1738 217174
rect -1654 216938 -1418 217174
rect -1974 216618 -1738 216854
rect -1654 216618 -1418 216854
rect -1974 179938 -1738 180174
rect -1654 179938 -1418 180174
rect -1974 179618 -1738 179854
rect -1654 179618 -1418 179854
rect -1974 142938 -1738 143174
rect -1654 142938 -1418 143174
rect -1974 142618 -1738 142854
rect -1654 142618 -1418 142854
rect -1974 105938 -1738 106174
rect -1654 105938 -1418 106174
rect -1974 105618 -1738 105854
rect -1654 105618 -1418 105854
rect -1974 68938 -1738 69174
rect -1654 68938 -1418 69174
rect -1974 68618 -1738 68854
rect -1654 68618 -1418 68854
rect -1974 31938 -1738 32174
rect -1654 31938 -1418 32174
rect -1974 31618 -1738 31854
rect -1654 31618 -1418 31854
rect 38026 583218 38262 583454
rect 38346 583218 38582 583454
rect 38026 582898 38262 583134
rect 38346 582898 38582 583134
rect 38026 546218 38262 546454
rect 38346 546218 38582 546454
rect 38026 545898 38262 546134
rect 38346 545898 38582 546134
rect 38026 509218 38262 509454
rect 38346 509218 38582 509454
rect 38026 508898 38262 509134
rect 38346 508898 38582 509134
rect 38026 472218 38262 472454
rect 38346 472218 38582 472454
rect 38026 471898 38262 472134
rect 38346 471898 38582 472134
rect 38026 435218 38262 435454
rect 38346 435218 38582 435454
rect 38026 434898 38262 435134
rect 38346 434898 38582 435134
rect 38026 398218 38262 398454
rect 38346 398218 38582 398454
rect 38026 397898 38262 398134
rect 38346 397898 38582 398134
rect 38026 361218 38262 361454
rect 38346 361218 38582 361454
rect 38026 360898 38262 361134
rect 38346 360898 38582 361134
rect 38026 324218 38262 324454
rect 38346 324218 38582 324454
rect 38026 323898 38262 324134
rect 38346 323898 38582 324134
rect 38026 287218 38262 287454
rect 38346 287218 38582 287454
rect 38026 286898 38262 287134
rect 38346 286898 38582 287134
rect 38026 250218 38262 250454
rect 38346 250218 38582 250454
rect 38026 249898 38262 250134
rect 38346 249898 38582 250134
rect 38026 213218 38262 213454
rect 38346 213218 38582 213454
rect 38026 212898 38262 213134
rect 38346 212898 38582 213134
rect 38026 176218 38262 176454
rect 38346 176218 38582 176454
rect 38026 175898 38262 176134
rect 38346 175898 38582 176134
rect 38026 139218 38262 139454
rect 38346 139218 38582 139454
rect 38026 138898 38262 139134
rect 38346 138898 38582 139134
rect 38026 102218 38262 102454
rect 38346 102218 38582 102454
rect 38026 101898 38262 102134
rect 38346 101898 38582 102134
rect 38026 65218 38262 65454
rect 38346 65218 38582 65454
rect 38026 64898 38262 65134
rect 38346 64898 38582 65134
rect 26460 31938 26696 32174
rect 26460 31618 26696 31854
rect 37408 31938 37644 32174
rect 37408 31618 37644 31854
rect 31934 28218 32170 28454
rect 31934 27898 32170 28134
rect 38026 28218 38262 28454
rect 38346 28218 38582 28454
rect 38026 27898 38262 28134
rect 38346 27898 38582 28134
rect -1974 -582 -1738 -346
rect -1654 -582 -1418 -346
rect -1974 -902 -1738 -666
rect -1654 -902 -1418 -666
rect -2934 -1542 -2698 -1306
rect -2614 -1542 -2378 -1306
rect -2934 -1862 -2698 -1626
rect -2614 -1862 -2378 -1626
rect 38026 -1542 38262 -1306
rect 38346 -1542 38582 -1306
rect 38026 -1862 38262 -1626
rect 38346 -1862 38582 -1626
rect -3894 -2502 -3658 -2266
rect -3574 -2502 -3338 -2266
rect -3894 -2822 -3658 -2586
rect -3574 -2822 -3338 -2586
rect -4854 -3462 -4618 -3226
rect -4534 -3462 -4298 -3226
rect -4854 -3782 -4618 -3546
rect -4534 -3782 -4298 -3546
rect -5814 -4422 -5578 -4186
rect -5494 -4422 -5258 -4186
rect -5814 -4742 -5578 -4506
rect -5494 -4742 -5258 -4506
rect -6774 -5382 -6538 -5146
rect -6454 -5382 -6218 -5146
rect -6774 -5702 -6538 -5466
rect -6454 -5702 -6218 -5466
rect -7734 -6342 -7498 -6106
rect -7414 -6342 -7178 -6106
rect -7734 -6662 -7498 -6426
rect -7414 -6662 -7178 -6426
rect -8694 -7302 -8458 -7066
rect -8374 -7302 -8138 -7066
rect -8694 -7622 -8458 -7386
rect -8374 -7622 -8138 -7386
rect 41746 704602 41982 704838
rect 42066 704602 42302 704838
rect 41746 704282 41982 704518
rect 42066 704282 42302 704518
rect 41746 697938 41982 698174
rect 42066 697938 42302 698174
rect 41746 697618 41982 697854
rect 42066 697618 42302 697854
rect 41746 660938 41982 661174
rect 42066 660938 42302 661174
rect 41746 660618 41982 660854
rect 42066 660618 42302 660854
rect 41746 623938 41982 624174
rect 42066 623938 42302 624174
rect 41746 623618 41982 623854
rect 42066 623618 42302 623854
rect 41746 586938 41982 587174
rect 42066 586938 42302 587174
rect 41746 586618 41982 586854
rect 42066 586618 42302 586854
rect 41746 549938 41982 550174
rect 42066 549938 42302 550174
rect 41746 549618 41982 549854
rect 42066 549618 42302 549854
rect 41746 512938 41982 513174
rect 42066 512938 42302 513174
rect 41746 512618 41982 512854
rect 42066 512618 42302 512854
rect 41746 475938 41982 476174
rect 42066 475938 42302 476174
rect 41746 475618 41982 475854
rect 42066 475618 42302 475854
rect 41746 438938 41982 439174
rect 42066 438938 42302 439174
rect 41746 438618 41982 438854
rect 42066 438618 42302 438854
rect 41746 401938 41982 402174
rect 42066 401938 42302 402174
rect 41746 401618 41982 401854
rect 42066 401618 42302 401854
rect 41746 364938 41982 365174
rect 42066 364938 42302 365174
rect 41746 364618 41982 364854
rect 42066 364618 42302 364854
rect 41746 327938 41982 328174
rect 42066 327938 42302 328174
rect 41746 327618 41982 327854
rect 42066 327618 42302 327854
rect 41746 290938 41982 291174
rect 42066 290938 42302 291174
rect 41746 290618 41982 290854
rect 42066 290618 42302 290854
rect 41746 253938 41982 254174
rect 42066 253938 42302 254174
rect 41746 253618 41982 253854
rect 42066 253618 42302 253854
rect 41746 216938 41982 217174
rect 42066 216938 42302 217174
rect 41746 216618 41982 216854
rect 42066 216618 42302 216854
rect 41746 179938 41982 180174
rect 42066 179938 42302 180174
rect 41746 179618 41982 179854
rect 42066 179618 42302 179854
rect 41746 142938 41982 143174
rect 42066 142938 42302 143174
rect 41746 142618 41982 142854
rect 42066 142618 42302 142854
rect 41746 105938 41982 106174
rect 42066 105938 42302 106174
rect 41746 105618 41982 105854
rect 42066 105618 42302 105854
rect 41746 68938 41982 69174
rect 42066 68938 42302 69174
rect 41746 68618 41982 68854
rect 42066 68618 42302 68854
rect 66026 705562 66262 705798
rect 66346 705562 66582 705798
rect 66026 705242 66262 705478
rect 66346 705242 66582 705478
rect 66026 694218 66262 694454
rect 66346 694218 66582 694454
rect 66026 693898 66262 694134
rect 66346 693898 66582 694134
rect 66026 657218 66262 657454
rect 66346 657218 66582 657454
rect 66026 656898 66262 657134
rect 66346 656898 66582 657134
rect 66026 620218 66262 620454
rect 66346 620218 66582 620454
rect 66026 619898 66262 620134
rect 66346 619898 66582 620134
rect 66026 583218 66262 583454
rect 66346 583218 66582 583454
rect 66026 582898 66262 583134
rect 66346 582898 66582 583134
rect 66026 546218 66262 546454
rect 66346 546218 66582 546454
rect 66026 545898 66262 546134
rect 66346 545898 66582 546134
rect 66026 509218 66262 509454
rect 66346 509218 66582 509454
rect 66026 508898 66262 509134
rect 66346 508898 66582 509134
rect 66026 472218 66262 472454
rect 66346 472218 66582 472454
rect 66026 471898 66262 472134
rect 66346 471898 66582 472134
rect 66026 435218 66262 435454
rect 66346 435218 66582 435454
rect 66026 434898 66262 435134
rect 66346 434898 66582 435134
rect 66026 398218 66262 398454
rect 66346 398218 66582 398454
rect 66026 397898 66262 398134
rect 66346 397898 66582 398134
rect 66026 361218 66262 361454
rect 66346 361218 66582 361454
rect 66026 360898 66262 361134
rect 66346 360898 66582 361134
rect 66026 324218 66262 324454
rect 66346 324218 66582 324454
rect 66026 323898 66262 324134
rect 66346 323898 66582 324134
rect 66026 287218 66262 287454
rect 66346 287218 66582 287454
rect 66026 286898 66262 287134
rect 66346 286898 66582 287134
rect 66026 250218 66262 250454
rect 66346 250218 66582 250454
rect 66026 249898 66262 250134
rect 66346 249898 66582 250134
rect 66026 213218 66262 213454
rect 66346 213218 66582 213454
rect 66026 212898 66262 213134
rect 66346 212898 66582 213134
rect 66026 176218 66262 176454
rect 66346 176218 66582 176454
rect 66026 175898 66262 176134
rect 66346 175898 66582 176134
rect 66026 139218 66262 139454
rect 66346 139218 66582 139454
rect 66026 138898 66262 139134
rect 66346 138898 66582 139134
rect 66026 102218 66262 102454
rect 66346 102218 66582 102454
rect 66026 101898 66262 102134
rect 66346 101898 66582 102134
rect 66026 65218 66262 65454
rect 66346 65218 66582 65454
rect 66026 64898 66262 65134
rect 66346 64898 66582 65134
rect 41746 31938 41982 32174
rect 42066 31938 42302 32174
rect 41746 31618 41982 31854
rect 42066 31618 42302 31854
rect 42882 28218 43118 28454
rect 42882 27898 43118 28134
rect 48356 31938 48592 32174
rect 48356 31618 48592 31854
rect 53830 28218 54066 28454
rect 53830 27898 54066 28134
rect 59304 31938 59540 32174
rect 59304 31618 59540 31854
rect 64778 28218 65014 28454
rect 64778 27898 65014 28134
rect 66026 28218 66262 28454
rect 66346 28218 66582 28454
rect 66026 27898 66262 28134
rect 66346 27898 66582 28134
rect 41746 -582 41982 -346
rect 42066 -582 42302 -346
rect 41746 -902 41982 -666
rect 42066 -902 42302 -666
rect 66026 -1542 66262 -1306
rect 66346 -1542 66582 -1306
rect 66026 -1862 66262 -1626
rect 66346 -1862 66582 -1626
rect 69746 704602 69982 704838
rect 70066 704602 70302 704838
rect 69746 704282 69982 704518
rect 70066 704282 70302 704518
rect 69746 697938 69982 698174
rect 70066 697938 70302 698174
rect 69746 697618 69982 697854
rect 70066 697618 70302 697854
rect 69746 660938 69982 661174
rect 70066 660938 70302 661174
rect 69746 660618 69982 660854
rect 70066 660618 70302 660854
rect 69746 623938 69982 624174
rect 70066 623938 70302 624174
rect 69746 623618 69982 623854
rect 70066 623618 70302 623854
rect 69746 586938 69982 587174
rect 70066 586938 70302 587174
rect 69746 586618 69982 586854
rect 70066 586618 70302 586854
rect 69746 549938 69982 550174
rect 70066 549938 70302 550174
rect 69746 549618 69982 549854
rect 70066 549618 70302 549854
rect 69746 512938 69982 513174
rect 70066 512938 70302 513174
rect 69746 512618 69982 512854
rect 70066 512618 70302 512854
rect 69746 475938 69982 476174
rect 70066 475938 70302 476174
rect 69746 475618 69982 475854
rect 70066 475618 70302 475854
rect 69746 438938 69982 439174
rect 70066 438938 70302 439174
rect 69746 438618 69982 438854
rect 70066 438618 70302 438854
rect 69746 401938 69982 402174
rect 70066 401938 70302 402174
rect 69746 401618 69982 401854
rect 70066 401618 70302 401854
rect 69746 364938 69982 365174
rect 70066 364938 70302 365174
rect 69746 364618 69982 364854
rect 70066 364618 70302 364854
rect 69746 327938 69982 328174
rect 70066 327938 70302 328174
rect 69746 327618 69982 327854
rect 70066 327618 70302 327854
rect 69746 290938 69982 291174
rect 70066 290938 70302 291174
rect 69746 290618 69982 290854
rect 70066 290618 70302 290854
rect 69746 253938 69982 254174
rect 70066 253938 70302 254174
rect 69746 253618 69982 253854
rect 70066 253618 70302 253854
rect 69746 216938 69982 217174
rect 70066 216938 70302 217174
rect 69746 216618 69982 216854
rect 70066 216618 70302 216854
rect 69746 179938 69982 180174
rect 70066 179938 70302 180174
rect 69746 179618 69982 179854
rect 70066 179618 70302 179854
rect 69746 142938 69982 143174
rect 70066 142938 70302 143174
rect 69746 142618 69982 142854
rect 70066 142618 70302 142854
rect 69746 105938 69982 106174
rect 70066 105938 70302 106174
rect 69746 105618 69982 105854
rect 70066 105618 70302 105854
rect 69746 68938 69982 69174
rect 70066 68938 70302 69174
rect 69746 68618 69982 68854
rect 70066 68618 70302 68854
rect 94026 705562 94262 705798
rect 94346 705562 94582 705798
rect 94026 705242 94262 705478
rect 94346 705242 94582 705478
rect 94026 694218 94262 694454
rect 94346 694218 94582 694454
rect 94026 693898 94262 694134
rect 94346 693898 94582 694134
rect 94026 657218 94262 657454
rect 94346 657218 94582 657454
rect 94026 656898 94262 657134
rect 94346 656898 94582 657134
rect 94026 620218 94262 620454
rect 94346 620218 94582 620454
rect 94026 619898 94262 620134
rect 94346 619898 94582 620134
rect 94026 583218 94262 583454
rect 94346 583218 94582 583454
rect 94026 582898 94262 583134
rect 94346 582898 94582 583134
rect 94026 546218 94262 546454
rect 94346 546218 94582 546454
rect 94026 545898 94262 546134
rect 94346 545898 94582 546134
rect 94026 509218 94262 509454
rect 94346 509218 94582 509454
rect 94026 508898 94262 509134
rect 94346 508898 94582 509134
rect 94026 472218 94262 472454
rect 94346 472218 94582 472454
rect 94026 471898 94262 472134
rect 94346 471898 94582 472134
rect 94026 435218 94262 435454
rect 94346 435218 94582 435454
rect 94026 434898 94262 435134
rect 94346 434898 94582 435134
rect 94026 398218 94262 398454
rect 94346 398218 94582 398454
rect 94026 397898 94262 398134
rect 94346 397898 94582 398134
rect 94026 361218 94262 361454
rect 94346 361218 94582 361454
rect 94026 360898 94262 361134
rect 94346 360898 94582 361134
rect 94026 324218 94262 324454
rect 94346 324218 94582 324454
rect 94026 323898 94262 324134
rect 94346 323898 94582 324134
rect 94026 287218 94262 287454
rect 94346 287218 94582 287454
rect 94026 286898 94262 287134
rect 94346 286898 94582 287134
rect 94026 250218 94262 250454
rect 94346 250218 94582 250454
rect 94026 249898 94262 250134
rect 94346 249898 94582 250134
rect 94026 213218 94262 213454
rect 94346 213218 94582 213454
rect 94026 212898 94262 213134
rect 94346 212898 94582 213134
rect 94026 176218 94262 176454
rect 94346 176218 94582 176454
rect 94026 175898 94262 176134
rect 94346 175898 94582 176134
rect 94026 139218 94262 139454
rect 94346 139218 94582 139454
rect 94026 138898 94262 139134
rect 94346 138898 94582 139134
rect 94026 102218 94262 102454
rect 94346 102218 94582 102454
rect 94026 101898 94262 102134
rect 94346 101898 94582 102134
rect 94026 65218 94262 65454
rect 94346 65218 94582 65454
rect 94026 64898 94262 65134
rect 94346 64898 94582 65134
rect 97746 704602 97982 704838
rect 98066 704602 98302 704838
rect 97746 704282 97982 704518
rect 98066 704282 98302 704518
rect 97746 697938 97982 698174
rect 98066 697938 98302 698174
rect 97746 697618 97982 697854
rect 98066 697618 98302 697854
rect 97746 660938 97982 661174
rect 98066 660938 98302 661174
rect 97746 660618 97982 660854
rect 98066 660618 98302 660854
rect 97746 623938 97982 624174
rect 98066 623938 98302 624174
rect 97746 623618 97982 623854
rect 98066 623618 98302 623854
rect 97746 586938 97982 587174
rect 98066 586938 98302 587174
rect 97746 586618 97982 586854
rect 98066 586618 98302 586854
rect 97746 549938 97982 550174
rect 98066 549938 98302 550174
rect 97746 549618 97982 549854
rect 98066 549618 98302 549854
rect 97746 512938 97982 513174
rect 98066 512938 98302 513174
rect 97746 512618 97982 512854
rect 98066 512618 98302 512854
rect 97746 475938 97982 476174
rect 98066 475938 98302 476174
rect 97746 475618 97982 475854
rect 98066 475618 98302 475854
rect 97746 438938 97982 439174
rect 98066 438938 98302 439174
rect 97746 438618 97982 438854
rect 98066 438618 98302 438854
rect 97746 401938 97982 402174
rect 98066 401938 98302 402174
rect 97746 401618 97982 401854
rect 98066 401618 98302 401854
rect 97746 364938 97982 365174
rect 98066 364938 98302 365174
rect 97746 364618 97982 364854
rect 98066 364618 98302 364854
rect 97746 327938 97982 328174
rect 98066 327938 98302 328174
rect 97746 327618 97982 327854
rect 98066 327618 98302 327854
rect 97746 290938 97982 291174
rect 98066 290938 98302 291174
rect 97746 290618 97982 290854
rect 98066 290618 98302 290854
rect 97746 253938 97982 254174
rect 98066 253938 98302 254174
rect 97746 253618 97982 253854
rect 98066 253618 98302 253854
rect 97746 216938 97982 217174
rect 98066 216938 98302 217174
rect 97746 216618 97982 216854
rect 98066 216618 98302 216854
rect 97746 179938 97982 180174
rect 98066 179938 98302 180174
rect 97746 179618 97982 179854
rect 98066 179618 98302 179854
rect 97746 142938 97982 143174
rect 98066 142938 98302 143174
rect 97746 142618 97982 142854
rect 98066 142618 98302 142854
rect 97746 105938 97982 106174
rect 98066 105938 98302 106174
rect 97746 105618 97982 105854
rect 98066 105618 98302 105854
rect 97746 68938 97982 69174
rect 98066 68938 98302 69174
rect 97746 68618 97982 68854
rect 98066 68618 98302 68854
rect 69746 31938 69982 32174
rect 70066 31938 70302 32174
rect 69746 31618 69982 31854
rect 70066 31618 70302 31854
rect 91860 31938 92096 32174
rect 91860 31618 92096 31854
rect 92808 31938 93044 32174
rect 92808 31618 93044 31854
rect 93756 31938 93992 32174
rect 93756 31618 93992 31854
rect 94704 31938 94940 32174
rect 94704 31618 94940 31854
rect 122026 705562 122262 705798
rect 122346 705562 122582 705798
rect 122026 705242 122262 705478
rect 122346 705242 122582 705478
rect 122026 694218 122262 694454
rect 122346 694218 122582 694454
rect 122026 693898 122262 694134
rect 122346 693898 122582 694134
rect 122026 657218 122262 657454
rect 122346 657218 122582 657454
rect 122026 656898 122262 657134
rect 122346 656898 122582 657134
rect 122026 620218 122262 620454
rect 122346 620218 122582 620454
rect 122026 619898 122262 620134
rect 122346 619898 122582 620134
rect 122026 583218 122262 583454
rect 122346 583218 122582 583454
rect 122026 582898 122262 583134
rect 122346 582898 122582 583134
rect 122026 546218 122262 546454
rect 122346 546218 122582 546454
rect 122026 545898 122262 546134
rect 122346 545898 122582 546134
rect 122026 509218 122262 509454
rect 122346 509218 122582 509454
rect 122026 508898 122262 509134
rect 122346 508898 122582 509134
rect 122026 472218 122262 472454
rect 122346 472218 122582 472454
rect 122026 471898 122262 472134
rect 122346 471898 122582 472134
rect 122026 435218 122262 435454
rect 122346 435218 122582 435454
rect 122026 434898 122262 435134
rect 122346 434898 122582 435134
rect 122026 398218 122262 398454
rect 122346 398218 122582 398454
rect 122026 397898 122262 398134
rect 122346 397898 122582 398134
rect 122026 361218 122262 361454
rect 122346 361218 122582 361454
rect 122026 360898 122262 361134
rect 122346 360898 122582 361134
rect 122026 324218 122262 324454
rect 122346 324218 122582 324454
rect 122026 323898 122262 324134
rect 122346 323898 122582 324134
rect 122026 287218 122262 287454
rect 122346 287218 122582 287454
rect 122026 286898 122262 287134
rect 122346 286898 122582 287134
rect 122026 250218 122262 250454
rect 122346 250218 122582 250454
rect 122026 249898 122262 250134
rect 122346 249898 122582 250134
rect 122026 213218 122262 213454
rect 122346 213218 122582 213454
rect 122026 212898 122262 213134
rect 122346 212898 122582 213134
rect 122026 176218 122262 176454
rect 122346 176218 122582 176454
rect 122026 175898 122262 176134
rect 122346 175898 122582 176134
rect 122026 139218 122262 139454
rect 122346 139218 122582 139454
rect 122026 138898 122262 139134
rect 122346 138898 122582 139134
rect 122026 102218 122262 102454
rect 122346 102218 122582 102454
rect 122026 101898 122262 102134
rect 122346 101898 122582 102134
rect 122026 65218 122262 65454
rect 122346 65218 122582 65454
rect 122026 64898 122262 65134
rect 122346 64898 122582 65134
rect 97746 31938 97982 32174
rect 98066 31938 98302 32174
rect 97746 31618 97982 31854
rect 98066 31618 98302 31854
rect 92334 28218 92570 28454
rect 92334 27898 92570 28134
rect 93282 28218 93518 28454
rect 93282 27898 93518 28134
rect 94230 28218 94466 28454
rect 94230 27898 94466 28134
rect 69746 -582 69982 -346
rect 70066 -582 70302 -346
rect 69746 -902 69982 -666
rect 70066 -902 70302 -666
rect 102059 31938 102295 32174
rect 102059 31618 102295 31854
rect 109005 31938 109241 32174
rect 109005 31618 109241 31854
rect 115951 31938 116187 32174
rect 115951 31618 116187 31854
rect 105532 28218 105768 28454
rect 105532 27898 105768 28134
rect 112478 28218 112714 28454
rect 112478 27898 112714 28134
rect 119424 28218 119660 28454
rect 119424 27898 119660 28134
rect 125746 704602 125982 704838
rect 126066 704602 126302 704838
rect 125746 704282 125982 704518
rect 126066 704282 126302 704518
rect 125746 697938 125982 698174
rect 126066 697938 126302 698174
rect 125746 697618 125982 697854
rect 126066 697618 126302 697854
rect 125746 660938 125982 661174
rect 126066 660938 126302 661174
rect 125746 660618 125982 660854
rect 126066 660618 126302 660854
rect 125746 623938 125982 624174
rect 126066 623938 126302 624174
rect 125746 623618 125982 623854
rect 126066 623618 126302 623854
rect 125746 586938 125982 587174
rect 126066 586938 126302 587174
rect 125746 586618 125982 586854
rect 126066 586618 126302 586854
rect 125746 549938 125982 550174
rect 126066 549938 126302 550174
rect 125746 549618 125982 549854
rect 126066 549618 126302 549854
rect 125746 512938 125982 513174
rect 126066 512938 126302 513174
rect 125746 512618 125982 512854
rect 126066 512618 126302 512854
rect 125746 475938 125982 476174
rect 126066 475938 126302 476174
rect 125746 475618 125982 475854
rect 126066 475618 126302 475854
rect 125746 438938 125982 439174
rect 126066 438938 126302 439174
rect 125746 438618 125982 438854
rect 126066 438618 126302 438854
rect 125746 401938 125982 402174
rect 126066 401938 126302 402174
rect 125746 401618 125982 401854
rect 126066 401618 126302 401854
rect 125746 364938 125982 365174
rect 126066 364938 126302 365174
rect 125746 364618 125982 364854
rect 126066 364618 126302 364854
rect 125746 327938 125982 328174
rect 126066 327938 126302 328174
rect 125746 327618 125982 327854
rect 126066 327618 126302 327854
rect 125746 290938 125982 291174
rect 126066 290938 126302 291174
rect 125746 290618 125982 290854
rect 126066 290618 126302 290854
rect 125746 253938 125982 254174
rect 126066 253938 126302 254174
rect 125746 253618 125982 253854
rect 126066 253618 126302 253854
rect 125746 216938 125982 217174
rect 126066 216938 126302 217174
rect 125746 216618 125982 216854
rect 126066 216618 126302 216854
rect 125746 179938 125982 180174
rect 126066 179938 126302 180174
rect 125746 179618 125982 179854
rect 126066 179618 126302 179854
rect 125746 142938 125982 143174
rect 126066 142938 126302 143174
rect 125746 142618 125982 142854
rect 126066 142618 126302 142854
rect 125746 105938 125982 106174
rect 126066 105938 126302 106174
rect 125746 105618 125982 105854
rect 126066 105618 126302 105854
rect 125746 68938 125982 69174
rect 126066 68938 126302 69174
rect 125746 68618 125982 68854
rect 126066 68618 126302 68854
rect 150026 705562 150262 705798
rect 150346 705562 150582 705798
rect 150026 705242 150262 705478
rect 150346 705242 150582 705478
rect 150026 694218 150262 694454
rect 150346 694218 150582 694454
rect 150026 693898 150262 694134
rect 150346 693898 150582 694134
rect 150026 657218 150262 657454
rect 150346 657218 150582 657454
rect 150026 656898 150262 657134
rect 150346 656898 150582 657134
rect 150026 620218 150262 620454
rect 150346 620218 150582 620454
rect 150026 619898 150262 620134
rect 150346 619898 150582 620134
rect 150026 583218 150262 583454
rect 150346 583218 150582 583454
rect 150026 582898 150262 583134
rect 150346 582898 150582 583134
rect 150026 546218 150262 546454
rect 150346 546218 150582 546454
rect 150026 545898 150262 546134
rect 150346 545898 150582 546134
rect 150026 509218 150262 509454
rect 150346 509218 150582 509454
rect 150026 508898 150262 509134
rect 150346 508898 150582 509134
rect 150026 472218 150262 472454
rect 150346 472218 150582 472454
rect 150026 471898 150262 472134
rect 150346 471898 150582 472134
rect 150026 435218 150262 435454
rect 150346 435218 150582 435454
rect 150026 434898 150262 435134
rect 150346 434898 150582 435134
rect 150026 398218 150262 398454
rect 150346 398218 150582 398454
rect 150026 397898 150262 398134
rect 150346 397898 150582 398134
rect 150026 361218 150262 361454
rect 150346 361218 150582 361454
rect 150026 360898 150262 361134
rect 150346 360898 150582 361134
rect 150026 324218 150262 324454
rect 150346 324218 150582 324454
rect 150026 323898 150262 324134
rect 150346 323898 150582 324134
rect 150026 287218 150262 287454
rect 150346 287218 150582 287454
rect 150026 286898 150262 287134
rect 150346 286898 150582 287134
rect 150026 250218 150262 250454
rect 150346 250218 150582 250454
rect 150026 249898 150262 250134
rect 150346 249898 150582 250134
rect 150026 213218 150262 213454
rect 150346 213218 150582 213454
rect 150026 212898 150262 213134
rect 150346 212898 150582 213134
rect 150026 176218 150262 176454
rect 150346 176218 150582 176454
rect 150026 175898 150262 176134
rect 150346 175898 150582 176134
rect 150026 139218 150262 139454
rect 150346 139218 150582 139454
rect 150026 138898 150262 139134
rect 150346 138898 150582 139134
rect 150026 102218 150262 102454
rect 150346 102218 150582 102454
rect 150026 101898 150262 102134
rect 150346 101898 150582 102134
rect 150026 65218 150262 65454
rect 150346 65218 150582 65454
rect 150026 64898 150262 65134
rect 150346 64898 150582 65134
rect 122897 31938 123133 32174
rect 122897 31618 123133 31854
rect 132060 31938 132296 32174
rect 132060 31618 132296 31854
rect 133008 31938 133244 32174
rect 133008 31618 133244 31854
rect 133956 31938 134192 32174
rect 133956 31618 134192 31854
rect 134904 31938 135140 32174
rect 134904 31618 135140 31854
rect 142259 31938 142495 32174
rect 142259 31618 142495 31854
rect 149205 31938 149441 32174
rect 149205 31618 149441 31854
rect 122026 28218 122262 28454
rect 122346 28218 122582 28454
rect 122026 27898 122262 28134
rect 122346 27898 122582 28134
rect 97746 -582 97982 -346
rect 98066 -582 98302 -346
rect 97746 -902 97982 -666
rect 98066 -902 98302 -666
rect 126370 28218 126606 28454
rect 126370 27898 126606 28134
rect 132534 28218 132770 28454
rect 132534 27898 132770 28134
rect 133482 28218 133718 28454
rect 133482 27898 133718 28134
rect 134430 28218 134666 28454
rect 134430 27898 134666 28134
rect 145732 28218 145968 28454
rect 145732 27898 145968 28134
rect 153746 704602 153982 704838
rect 154066 704602 154302 704838
rect 153746 704282 153982 704518
rect 154066 704282 154302 704518
rect 153746 697938 153982 698174
rect 154066 697938 154302 698174
rect 153746 697618 153982 697854
rect 154066 697618 154302 697854
rect 153746 660938 153982 661174
rect 154066 660938 154302 661174
rect 153746 660618 153982 660854
rect 154066 660618 154302 660854
rect 153746 623938 153982 624174
rect 154066 623938 154302 624174
rect 153746 623618 153982 623854
rect 154066 623618 154302 623854
rect 153746 586938 153982 587174
rect 154066 586938 154302 587174
rect 153746 586618 153982 586854
rect 154066 586618 154302 586854
rect 153746 549938 153982 550174
rect 154066 549938 154302 550174
rect 153746 549618 153982 549854
rect 154066 549618 154302 549854
rect 153746 512938 153982 513174
rect 154066 512938 154302 513174
rect 153746 512618 153982 512854
rect 154066 512618 154302 512854
rect 153746 475938 153982 476174
rect 154066 475938 154302 476174
rect 153746 475618 153982 475854
rect 154066 475618 154302 475854
rect 153746 438938 153982 439174
rect 154066 438938 154302 439174
rect 153746 438618 153982 438854
rect 154066 438618 154302 438854
rect 153746 401938 153982 402174
rect 154066 401938 154302 402174
rect 153746 401618 153982 401854
rect 154066 401618 154302 401854
rect 153746 364938 153982 365174
rect 154066 364938 154302 365174
rect 153746 364618 153982 364854
rect 154066 364618 154302 364854
rect 153746 327938 153982 328174
rect 154066 327938 154302 328174
rect 153746 327618 153982 327854
rect 154066 327618 154302 327854
rect 153746 290938 153982 291174
rect 154066 290938 154302 291174
rect 153746 290618 153982 290854
rect 154066 290618 154302 290854
rect 153746 253938 153982 254174
rect 154066 253938 154302 254174
rect 153746 253618 153982 253854
rect 154066 253618 154302 253854
rect 153746 216938 153982 217174
rect 154066 216938 154302 217174
rect 153746 216618 153982 216854
rect 154066 216618 154302 216854
rect 153746 179938 153982 180174
rect 154066 179938 154302 180174
rect 153746 179618 153982 179854
rect 154066 179618 154302 179854
rect 153746 142938 153982 143174
rect 154066 142938 154302 143174
rect 153746 142618 153982 142854
rect 154066 142618 154302 142854
rect 153746 105938 153982 106174
rect 154066 105938 154302 106174
rect 153746 105618 153982 105854
rect 154066 105618 154302 105854
rect 153746 68938 153982 69174
rect 154066 68938 154302 69174
rect 153746 68618 153982 68854
rect 154066 68618 154302 68854
rect 178026 705562 178262 705798
rect 178346 705562 178582 705798
rect 178026 705242 178262 705478
rect 178346 705242 178582 705478
rect 178026 694218 178262 694454
rect 178346 694218 178582 694454
rect 178026 693898 178262 694134
rect 178346 693898 178582 694134
rect 178026 657218 178262 657454
rect 178346 657218 178582 657454
rect 178026 656898 178262 657134
rect 178346 656898 178582 657134
rect 178026 620218 178262 620454
rect 178346 620218 178582 620454
rect 178026 619898 178262 620134
rect 178346 619898 178582 620134
rect 178026 583218 178262 583454
rect 178346 583218 178582 583454
rect 178026 582898 178262 583134
rect 178346 582898 178582 583134
rect 178026 546218 178262 546454
rect 178346 546218 178582 546454
rect 178026 545898 178262 546134
rect 178346 545898 178582 546134
rect 178026 509218 178262 509454
rect 178346 509218 178582 509454
rect 178026 508898 178262 509134
rect 178346 508898 178582 509134
rect 178026 472218 178262 472454
rect 178346 472218 178582 472454
rect 178026 471898 178262 472134
rect 178346 471898 178582 472134
rect 178026 435218 178262 435454
rect 178346 435218 178582 435454
rect 178026 434898 178262 435134
rect 178346 434898 178582 435134
rect 178026 398218 178262 398454
rect 178346 398218 178582 398454
rect 178026 397898 178262 398134
rect 178346 397898 178582 398134
rect 178026 361218 178262 361454
rect 178346 361218 178582 361454
rect 178026 360898 178262 361134
rect 178346 360898 178582 361134
rect 178026 324218 178262 324454
rect 178346 324218 178582 324454
rect 178026 323898 178262 324134
rect 178346 323898 178582 324134
rect 178026 287218 178262 287454
rect 178346 287218 178582 287454
rect 178026 286898 178262 287134
rect 178346 286898 178582 287134
rect 178026 250218 178262 250454
rect 178346 250218 178582 250454
rect 178026 249898 178262 250134
rect 178346 249898 178582 250134
rect 178026 213218 178262 213454
rect 178346 213218 178582 213454
rect 178026 212898 178262 213134
rect 178346 212898 178582 213134
rect 178026 176218 178262 176454
rect 178346 176218 178582 176454
rect 178026 175898 178262 176134
rect 178346 175898 178582 176134
rect 178026 139218 178262 139454
rect 178346 139218 178582 139454
rect 178026 138898 178262 139134
rect 178346 138898 178582 139134
rect 178026 102218 178262 102454
rect 178346 102218 178582 102454
rect 178026 101898 178262 102134
rect 178346 101898 178582 102134
rect 178026 65218 178262 65454
rect 178346 65218 178582 65454
rect 178026 64898 178262 65134
rect 178346 64898 178582 65134
rect 153746 31938 153982 32174
rect 154066 31938 154302 32174
rect 153746 31618 153982 31854
rect 154066 31618 154302 31854
rect 150026 28218 150262 28454
rect 150346 28218 150582 28454
rect 150026 27898 150262 28134
rect 150346 27898 150582 28134
rect 122026 -1542 122262 -1306
rect 122346 -1542 122582 -1306
rect 122026 -1862 122262 -1626
rect 122346 -1862 122582 -1626
rect 152678 28218 152914 28454
rect 152678 27898 152914 28134
rect 150026 -1542 150262 -1306
rect 150346 -1542 150582 -1306
rect 150026 -1862 150262 -1626
rect 150346 -1862 150582 -1626
rect 156151 31938 156387 32174
rect 156151 31618 156387 31854
rect 163097 31938 163333 32174
rect 163097 31618 163333 31854
rect 172260 31938 172496 32174
rect 172260 31618 172496 31854
rect 173208 31938 173444 32174
rect 173208 31618 173444 31854
rect 174156 31938 174392 32174
rect 174156 31618 174392 31854
rect 175104 31938 175340 32174
rect 175104 31618 175340 31854
rect 159624 28218 159860 28454
rect 159624 27898 159860 28134
rect 166570 28218 166806 28454
rect 166570 27898 166806 28134
rect 172734 28218 172970 28454
rect 172734 27898 172970 28134
rect 173682 28218 173918 28454
rect 173682 27898 173918 28134
rect 174630 28218 174866 28454
rect 174630 27898 174866 28134
rect 178026 28218 178262 28454
rect 178346 28218 178582 28454
rect 178026 27898 178262 28134
rect 178346 27898 178582 28134
rect 153746 -582 153982 -346
rect 154066 -582 154302 -346
rect 153746 -902 153982 -666
rect 154066 -902 154302 -666
rect 178026 -1542 178262 -1306
rect 178346 -1542 178582 -1306
rect 178026 -1862 178262 -1626
rect 178346 -1862 178582 -1626
rect 181746 704602 181982 704838
rect 182066 704602 182302 704838
rect 181746 704282 181982 704518
rect 182066 704282 182302 704518
rect 181746 697938 181982 698174
rect 182066 697938 182302 698174
rect 181746 697618 181982 697854
rect 182066 697618 182302 697854
rect 181746 660938 181982 661174
rect 182066 660938 182302 661174
rect 181746 660618 181982 660854
rect 182066 660618 182302 660854
rect 181746 623938 181982 624174
rect 182066 623938 182302 624174
rect 181746 623618 181982 623854
rect 182066 623618 182302 623854
rect 181746 586938 181982 587174
rect 182066 586938 182302 587174
rect 181746 586618 181982 586854
rect 182066 586618 182302 586854
rect 181746 549938 181982 550174
rect 182066 549938 182302 550174
rect 181746 549618 181982 549854
rect 182066 549618 182302 549854
rect 181746 512938 181982 513174
rect 182066 512938 182302 513174
rect 181746 512618 181982 512854
rect 182066 512618 182302 512854
rect 181746 475938 181982 476174
rect 182066 475938 182302 476174
rect 181746 475618 181982 475854
rect 182066 475618 182302 475854
rect 181746 438938 181982 439174
rect 182066 438938 182302 439174
rect 181746 438618 181982 438854
rect 182066 438618 182302 438854
rect 181746 401938 181982 402174
rect 182066 401938 182302 402174
rect 181746 401618 181982 401854
rect 182066 401618 182302 401854
rect 181746 364938 181982 365174
rect 182066 364938 182302 365174
rect 181746 364618 181982 364854
rect 182066 364618 182302 364854
rect 181746 327938 181982 328174
rect 182066 327938 182302 328174
rect 181746 327618 181982 327854
rect 182066 327618 182302 327854
rect 181746 290938 181982 291174
rect 182066 290938 182302 291174
rect 181746 290618 181982 290854
rect 182066 290618 182302 290854
rect 181746 253938 181982 254174
rect 182066 253938 182302 254174
rect 181746 253618 181982 253854
rect 182066 253618 182302 253854
rect 181746 216938 181982 217174
rect 182066 216938 182302 217174
rect 181746 216618 181982 216854
rect 182066 216618 182302 216854
rect 181746 179938 181982 180174
rect 182066 179938 182302 180174
rect 181746 179618 181982 179854
rect 182066 179618 182302 179854
rect 181746 142938 181982 143174
rect 182066 142938 182302 143174
rect 181746 142618 181982 142854
rect 182066 142618 182302 142854
rect 181746 105938 181982 106174
rect 182066 105938 182302 106174
rect 181746 105618 181982 105854
rect 182066 105618 182302 105854
rect 181746 68938 181982 69174
rect 182066 68938 182302 69174
rect 181746 68618 181982 68854
rect 182066 68618 182302 68854
rect 206026 705562 206262 705798
rect 206346 705562 206582 705798
rect 206026 705242 206262 705478
rect 206346 705242 206582 705478
rect 206026 694218 206262 694454
rect 206346 694218 206582 694454
rect 206026 693898 206262 694134
rect 206346 693898 206582 694134
rect 206026 657218 206262 657454
rect 206346 657218 206582 657454
rect 206026 656898 206262 657134
rect 206346 656898 206582 657134
rect 206026 620218 206262 620454
rect 206346 620218 206582 620454
rect 206026 619898 206262 620134
rect 206346 619898 206582 620134
rect 206026 583218 206262 583454
rect 206346 583218 206582 583454
rect 206026 582898 206262 583134
rect 206346 582898 206582 583134
rect 206026 546218 206262 546454
rect 206346 546218 206582 546454
rect 206026 545898 206262 546134
rect 206346 545898 206582 546134
rect 206026 509218 206262 509454
rect 206346 509218 206582 509454
rect 206026 508898 206262 509134
rect 206346 508898 206582 509134
rect 206026 472218 206262 472454
rect 206346 472218 206582 472454
rect 206026 471898 206262 472134
rect 206346 471898 206582 472134
rect 206026 435218 206262 435454
rect 206346 435218 206582 435454
rect 206026 434898 206262 435134
rect 206346 434898 206582 435134
rect 206026 398218 206262 398454
rect 206346 398218 206582 398454
rect 206026 397898 206262 398134
rect 206346 397898 206582 398134
rect 206026 361218 206262 361454
rect 206346 361218 206582 361454
rect 206026 360898 206262 361134
rect 206346 360898 206582 361134
rect 206026 324218 206262 324454
rect 206346 324218 206582 324454
rect 206026 323898 206262 324134
rect 206346 323898 206582 324134
rect 206026 287218 206262 287454
rect 206346 287218 206582 287454
rect 206026 286898 206262 287134
rect 206346 286898 206582 287134
rect 206026 250218 206262 250454
rect 206346 250218 206582 250454
rect 206026 249898 206262 250134
rect 206346 249898 206582 250134
rect 206026 213218 206262 213454
rect 206346 213218 206582 213454
rect 206026 212898 206262 213134
rect 206346 212898 206582 213134
rect 206026 176218 206262 176454
rect 206346 176218 206582 176454
rect 206026 175898 206262 176134
rect 206346 175898 206582 176134
rect 206026 139218 206262 139454
rect 206346 139218 206582 139454
rect 206026 138898 206262 139134
rect 206346 138898 206582 139134
rect 206026 102218 206262 102454
rect 206346 102218 206582 102454
rect 206026 101898 206262 102134
rect 206346 101898 206582 102134
rect 206026 65218 206262 65454
rect 206346 65218 206582 65454
rect 206026 64898 206262 65134
rect 206346 64898 206582 65134
rect 181746 31938 181982 32174
rect 182066 31938 182302 32174
rect 181746 31618 181982 31854
rect 182066 31618 182302 31854
rect 182459 31938 182695 32174
rect 182459 31618 182695 31854
rect 189405 31938 189641 32174
rect 189405 31618 189641 31854
rect 196351 31938 196587 32174
rect 196351 31618 196587 31854
rect 203297 31938 203533 32174
rect 203297 31618 203533 31854
rect 185932 28218 186168 28454
rect 185932 27898 186168 28134
rect 192878 28218 193114 28454
rect 192878 27898 193114 28134
rect 199824 28218 200060 28454
rect 199824 27898 200060 28134
rect 209746 704602 209982 704838
rect 210066 704602 210302 704838
rect 209746 704282 209982 704518
rect 210066 704282 210302 704518
rect 209746 697938 209982 698174
rect 210066 697938 210302 698174
rect 209746 697618 209982 697854
rect 210066 697618 210302 697854
rect 209746 660938 209982 661174
rect 210066 660938 210302 661174
rect 209746 660618 209982 660854
rect 210066 660618 210302 660854
rect 209746 623938 209982 624174
rect 210066 623938 210302 624174
rect 209746 623618 209982 623854
rect 210066 623618 210302 623854
rect 209746 586938 209982 587174
rect 210066 586938 210302 587174
rect 209746 586618 209982 586854
rect 210066 586618 210302 586854
rect 209746 549938 209982 550174
rect 210066 549938 210302 550174
rect 209746 549618 209982 549854
rect 210066 549618 210302 549854
rect 209746 512938 209982 513174
rect 210066 512938 210302 513174
rect 209746 512618 209982 512854
rect 210066 512618 210302 512854
rect 209746 475938 209982 476174
rect 210066 475938 210302 476174
rect 209746 475618 209982 475854
rect 210066 475618 210302 475854
rect 209746 438938 209982 439174
rect 210066 438938 210302 439174
rect 209746 438618 209982 438854
rect 210066 438618 210302 438854
rect 209746 401938 209982 402174
rect 210066 401938 210302 402174
rect 209746 401618 209982 401854
rect 210066 401618 210302 401854
rect 209746 364938 209982 365174
rect 210066 364938 210302 365174
rect 209746 364618 209982 364854
rect 210066 364618 210302 364854
rect 209746 327938 209982 328174
rect 210066 327938 210302 328174
rect 209746 327618 209982 327854
rect 210066 327618 210302 327854
rect 209746 290938 209982 291174
rect 210066 290938 210302 291174
rect 209746 290618 209982 290854
rect 210066 290618 210302 290854
rect 209746 253938 209982 254174
rect 210066 253938 210302 254174
rect 209746 253618 209982 253854
rect 210066 253618 210302 253854
rect 209746 216938 209982 217174
rect 210066 216938 210302 217174
rect 209746 216618 209982 216854
rect 210066 216618 210302 216854
rect 209746 179938 209982 180174
rect 210066 179938 210302 180174
rect 209746 179618 209982 179854
rect 210066 179618 210302 179854
rect 209746 142938 209982 143174
rect 210066 142938 210302 143174
rect 209746 142618 209982 142854
rect 210066 142618 210302 142854
rect 209746 105938 209982 106174
rect 210066 105938 210302 106174
rect 209746 105618 209982 105854
rect 210066 105618 210302 105854
rect 209746 68938 209982 69174
rect 210066 68938 210302 69174
rect 209746 68618 209982 68854
rect 210066 68618 210302 68854
rect 234026 705562 234262 705798
rect 234346 705562 234582 705798
rect 234026 705242 234262 705478
rect 234346 705242 234582 705478
rect 234026 694218 234262 694454
rect 234346 694218 234582 694454
rect 234026 693898 234262 694134
rect 234346 693898 234582 694134
rect 234026 657218 234262 657454
rect 234346 657218 234582 657454
rect 234026 656898 234262 657134
rect 234346 656898 234582 657134
rect 234026 620218 234262 620454
rect 234346 620218 234582 620454
rect 234026 619898 234262 620134
rect 234346 619898 234582 620134
rect 234026 583218 234262 583454
rect 234346 583218 234582 583454
rect 234026 582898 234262 583134
rect 234346 582898 234582 583134
rect 234026 546218 234262 546454
rect 234346 546218 234582 546454
rect 234026 545898 234262 546134
rect 234346 545898 234582 546134
rect 234026 509218 234262 509454
rect 234346 509218 234582 509454
rect 234026 508898 234262 509134
rect 234346 508898 234582 509134
rect 234026 472218 234262 472454
rect 234346 472218 234582 472454
rect 234026 471898 234262 472134
rect 234346 471898 234582 472134
rect 234026 435218 234262 435454
rect 234346 435218 234582 435454
rect 234026 434898 234262 435134
rect 234346 434898 234582 435134
rect 234026 398218 234262 398454
rect 234346 398218 234582 398454
rect 234026 397898 234262 398134
rect 234346 397898 234582 398134
rect 234026 361218 234262 361454
rect 234346 361218 234582 361454
rect 234026 360898 234262 361134
rect 234346 360898 234582 361134
rect 234026 324218 234262 324454
rect 234346 324218 234582 324454
rect 234026 323898 234262 324134
rect 234346 323898 234582 324134
rect 234026 287218 234262 287454
rect 234346 287218 234582 287454
rect 234026 286898 234262 287134
rect 234346 286898 234582 287134
rect 234026 250218 234262 250454
rect 234346 250218 234582 250454
rect 234026 249898 234262 250134
rect 234346 249898 234582 250134
rect 234026 213218 234262 213454
rect 234346 213218 234582 213454
rect 234026 212898 234262 213134
rect 234346 212898 234582 213134
rect 234026 176218 234262 176454
rect 234346 176218 234582 176454
rect 234026 175898 234262 176134
rect 234346 175898 234582 176134
rect 234026 139218 234262 139454
rect 234346 139218 234582 139454
rect 234026 138898 234262 139134
rect 234346 138898 234582 139134
rect 234026 102218 234262 102454
rect 234346 102218 234582 102454
rect 234026 101898 234262 102134
rect 234346 101898 234582 102134
rect 234026 65218 234262 65454
rect 234346 65218 234582 65454
rect 234026 64898 234262 65134
rect 234346 64898 234582 65134
rect 237746 704602 237982 704838
rect 238066 704602 238302 704838
rect 237746 704282 237982 704518
rect 238066 704282 238302 704518
rect 237746 697938 237982 698174
rect 238066 697938 238302 698174
rect 237746 697618 237982 697854
rect 238066 697618 238302 697854
rect 237746 660938 237982 661174
rect 238066 660938 238302 661174
rect 237746 660618 237982 660854
rect 238066 660618 238302 660854
rect 237746 623938 237982 624174
rect 238066 623938 238302 624174
rect 237746 623618 237982 623854
rect 238066 623618 238302 623854
rect 237746 586938 237982 587174
rect 238066 586938 238302 587174
rect 237746 586618 237982 586854
rect 238066 586618 238302 586854
rect 237746 549938 237982 550174
rect 238066 549938 238302 550174
rect 237746 549618 237982 549854
rect 238066 549618 238302 549854
rect 237746 512938 237982 513174
rect 238066 512938 238302 513174
rect 237746 512618 237982 512854
rect 238066 512618 238302 512854
rect 237746 475938 237982 476174
rect 238066 475938 238302 476174
rect 237746 475618 237982 475854
rect 238066 475618 238302 475854
rect 237746 438938 237982 439174
rect 238066 438938 238302 439174
rect 237746 438618 237982 438854
rect 238066 438618 238302 438854
rect 237746 401938 237982 402174
rect 238066 401938 238302 402174
rect 237746 401618 237982 401854
rect 238066 401618 238302 401854
rect 237746 364938 237982 365174
rect 238066 364938 238302 365174
rect 237746 364618 237982 364854
rect 238066 364618 238302 364854
rect 237746 327938 237982 328174
rect 238066 327938 238302 328174
rect 237746 327618 237982 327854
rect 238066 327618 238302 327854
rect 237746 290938 237982 291174
rect 238066 290938 238302 291174
rect 237746 290618 237982 290854
rect 238066 290618 238302 290854
rect 237746 253938 237982 254174
rect 238066 253938 238302 254174
rect 237746 253618 237982 253854
rect 238066 253618 238302 253854
rect 237746 216938 237982 217174
rect 238066 216938 238302 217174
rect 237746 216618 237982 216854
rect 238066 216618 238302 216854
rect 237746 179938 237982 180174
rect 238066 179938 238302 180174
rect 237746 179618 237982 179854
rect 238066 179618 238302 179854
rect 237746 142938 237982 143174
rect 238066 142938 238302 143174
rect 237746 142618 237982 142854
rect 238066 142618 238302 142854
rect 237746 105938 237982 106174
rect 238066 105938 238302 106174
rect 237746 105618 237982 105854
rect 238066 105618 238302 105854
rect 237746 68938 237982 69174
rect 238066 68938 238302 69174
rect 237746 68618 237982 68854
rect 238066 68618 238302 68854
rect 262026 705562 262262 705798
rect 262346 705562 262582 705798
rect 262026 705242 262262 705478
rect 262346 705242 262582 705478
rect 262026 694218 262262 694454
rect 262346 694218 262582 694454
rect 262026 693898 262262 694134
rect 262346 693898 262582 694134
rect 262026 657218 262262 657454
rect 262346 657218 262582 657454
rect 262026 656898 262262 657134
rect 262346 656898 262582 657134
rect 262026 620218 262262 620454
rect 262346 620218 262582 620454
rect 262026 619898 262262 620134
rect 262346 619898 262582 620134
rect 262026 583218 262262 583454
rect 262346 583218 262582 583454
rect 262026 582898 262262 583134
rect 262346 582898 262582 583134
rect 262026 546218 262262 546454
rect 262346 546218 262582 546454
rect 262026 545898 262262 546134
rect 262346 545898 262582 546134
rect 262026 509218 262262 509454
rect 262346 509218 262582 509454
rect 262026 508898 262262 509134
rect 262346 508898 262582 509134
rect 262026 472218 262262 472454
rect 262346 472218 262582 472454
rect 262026 471898 262262 472134
rect 262346 471898 262582 472134
rect 262026 435218 262262 435454
rect 262346 435218 262582 435454
rect 262026 434898 262262 435134
rect 262346 434898 262582 435134
rect 262026 398218 262262 398454
rect 262346 398218 262582 398454
rect 262026 397898 262262 398134
rect 262346 397898 262582 398134
rect 262026 361218 262262 361454
rect 262346 361218 262582 361454
rect 262026 360898 262262 361134
rect 262346 360898 262582 361134
rect 262026 324218 262262 324454
rect 262346 324218 262582 324454
rect 262026 323898 262262 324134
rect 262346 323898 262582 324134
rect 262026 287218 262262 287454
rect 262346 287218 262582 287454
rect 262026 286898 262262 287134
rect 262346 286898 262582 287134
rect 262026 250218 262262 250454
rect 262346 250218 262582 250454
rect 262026 249898 262262 250134
rect 262346 249898 262582 250134
rect 262026 213218 262262 213454
rect 262346 213218 262582 213454
rect 262026 212898 262262 213134
rect 262346 212898 262582 213134
rect 262026 176218 262262 176454
rect 262346 176218 262582 176454
rect 262026 175898 262262 176134
rect 262346 175898 262582 176134
rect 262026 139218 262262 139454
rect 262346 139218 262582 139454
rect 262026 138898 262262 139134
rect 262346 138898 262582 139134
rect 262026 102218 262262 102454
rect 262346 102218 262582 102454
rect 262026 101898 262262 102134
rect 262346 101898 262582 102134
rect 262026 65218 262262 65454
rect 262346 65218 262582 65454
rect 262026 64898 262262 65134
rect 262346 64898 262582 65134
rect 265746 704602 265982 704838
rect 266066 704602 266302 704838
rect 265746 704282 265982 704518
rect 266066 704282 266302 704518
rect 265746 697938 265982 698174
rect 266066 697938 266302 698174
rect 265746 697618 265982 697854
rect 266066 697618 266302 697854
rect 265746 660938 265982 661174
rect 266066 660938 266302 661174
rect 265746 660618 265982 660854
rect 266066 660618 266302 660854
rect 265746 623938 265982 624174
rect 266066 623938 266302 624174
rect 265746 623618 265982 623854
rect 266066 623618 266302 623854
rect 265746 586938 265982 587174
rect 266066 586938 266302 587174
rect 265746 586618 265982 586854
rect 266066 586618 266302 586854
rect 265746 549938 265982 550174
rect 266066 549938 266302 550174
rect 265746 549618 265982 549854
rect 266066 549618 266302 549854
rect 265746 512938 265982 513174
rect 266066 512938 266302 513174
rect 265746 512618 265982 512854
rect 266066 512618 266302 512854
rect 265746 475938 265982 476174
rect 266066 475938 266302 476174
rect 265746 475618 265982 475854
rect 266066 475618 266302 475854
rect 265746 438938 265982 439174
rect 266066 438938 266302 439174
rect 265746 438618 265982 438854
rect 266066 438618 266302 438854
rect 265746 401938 265982 402174
rect 266066 401938 266302 402174
rect 265746 401618 265982 401854
rect 266066 401618 266302 401854
rect 265746 364938 265982 365174
rect 266066 364938 266302 365174
rect 265746 364618 265982 364854
rect 266066 364618 266302 364854
rect 265746 327938 265982 328174
rect 266066 327938 266302 328174
rect 265746 327618 265982 327854
rect 266066 327618 266302 327854
rect 265746 290938 265982 291174
rect 266066 290938 266302 291174
rect 265746 290618 265982 290854
rect 266066 290618 266302 290854
rect 265746 253938 265982 254174
rect 266066 253938 266302 254174
rect 265746 253618 265982 253854
rect 266066 253618 266302 253854
rect 265746 216938 265982 217174
rect 266066 216938 266302 217174
rect 265746 216618 265982 216854
rect 266066 216618 266302 216854
rect 265746 179938 265982 180174
rect 266066 179938 266302 180174
rect 265746 179618 265982 179854
rect 266066 179618 266302 179854
rect 265746 142938 265982 143174
rect 266066 142938 266302 143174
rect 265746 142618 265982 142854
rect 266066 142618 266302 142854
rect 265746 105938 265982 106174
rect 266066 105938 266302 106174
rect 265746 105618 265982 105854
rect 266066 105618 266302 105854
rect 265746 68938 265982 69174
rect 266066 68938 266302 69174
rect 265746 68618 265982 68854
rect 266066 68618 266302 68854
rect 290026 705562 290262 705798
rect 290346 705562 290582 705798
rect 290026 705242 290262 705478
rect 290346 705242 290582 705478
rect 290026 694218 290262 694454
rect 290346 694218 290582 694454
rect 290026 693898 290262 694134
rect 290346 693898 290582 694134
rect 290026 657218 290262 657454
rect 290346 657218 290582 657454
rect 290026 656898 290262 657134
rect 290346 656898 290582 657134
rect 290026 620218 290262 620454
rect 290346 620218 290582 620454
rect 290026 619898 290262 620134
rect 290346 619898 290582 620134
rect 290026 583218 290262 583454
rect 290346 583218 290582 583454
rect 290026 582898 290262 583134
rect 290346 582898 290582 583134
rect 290026 546218 290262 546454
rect 290346 546218 290582 546454
rect 290026 545898 290262 546134
rect 290346 545898 290582 546134
rect 290026 509218 290262 509454
rect 290346 509218 290582 509454
rect 290026 508898 290262 509134
rect 290346 508898 290582 509134
rect 290026 472218 290262 472454
rect 290346 472218 290582 472454
rect 290026 471898 290262 472134
rect 290346 471898 290582 472134
rect 290026 435218 290262 435454
rect 290346 435218 290582 435454
rect 290026 434898 290262 435134
rect 290346 434898 290582 435134
rect 290026 398218 290262 398454
rect 290346 398218 290582 398454
rect 290026 397898 290262 398134
rect 290346 397898 290582 398134
rect 290026 361218 290262 361454
rect 290346 361218 290582 361454
rect 290026 360898 290262 361134
rect 290346 360898 290582 361134
rect 290026 324218 290262 324454
rect 290346 324218 290582 324454
rect 290026 323898 290262 324134
rect 290346 323898 290582 324134
rect 290026 287218 290262 287454
rect 290346 287218 290582 287454
rect 290026 286898 290262 287134
rect 290346 286898 290582 287134
rect 290026 250218 290262 250454
rect 290346 250218 290582 250454
rect 290026 249898 290262 250134
rect 290346 249898 290582 250134
rect 290026 213218 290262 213454
rect 290346 213218 290582 213454
rect 290026 212898 290262 213134
rect 290346 212898 290582 213134
rect 290026 176218 290262 176454
rect 290346 176218 290582 176454
rect 290026 175898 290262 176134
rect 290346 175898 290582 176134
rect 290026 139218 290262 139454
rect 290346 139218 290582 139454
rect 290026 138898 290262 139134
rect 290346 138898 290582 139134
rect 290026 102218 290262 102454
rect 290346 102218 290582 102454
rect 290026 101898 290262 102134
rect 290346 101898 290582 102134
rect 290026 65218 290262 65454
rect 290346 65218 290582 65454
rect 290026 64898 290262 65134
rect 290346 64898 290582 65134
rect 209746 31938 209982 32174
rect 210066 31938 210302 32174
rect 209746 31618 209982 31854
rect 210066 31618 210302 31854
rect 206026 28218 206262 28454
rect 206346 28218 206582 28454
rect 206026 27898 206262 28134
rect 206346 27898 206582 28134
rect 181746 -582 181982 -346
rect 182066 -582 182302 -346
rect 181746 -902 181982 -666
rect 182066 -902 182302 -666
rect 206770 28218 207006 28454
rect 206770 27898 207006 28134
rect 206026 -1542 206262 -1306
rect 206346 -1542 206582 -1306
rect 206026 -1862 206262 -1626
rect 206346 -1862 206582 -1626
rect 212460 31938 212696 32174
rect 212460 31618 212696 31854
rect 213408 31938 213644 32174
rect 213408 31618 213644 31854
rect 214356 31938 214592 32174
rect 214356 31618 214592 31854
rect 215304 31938 215540 32174
rect 215304 31618 215540 31854
rect 222659 31938 222895 32174
rect 222659 31618 222895 31854
rect 229605 31938 229841 32174
rect 229605 31618 229841 31854
rect 236551 31938 236787 32174
rect 236551 31618 236787 31854
rect 243497 31938 243733 32174
rect 243497 31618 243733 31854
rect 252660 31938 252896 32174
rect 252660 31618 252896 31854
rect 253608 31938 253844 32174
rect 253608 31618 253844 31854
rect 254556 31938 254792 32174
rect 254556 31618 254792 31854
rect 255504 31938 255740 32174
rect 255504 31618 255740 31854
rect 262859 31938 263095 32174
rect 262859 31618 263095 31854
rect 269805 31938 270041 32174
rect 269805 31618 270041 31854
rect 276751 31938 276987 32174
rect 276751 31618 276987 31854
rect 283697 31938 283933 32174
rect 283697 31618 283933 31854
rect 212934 28218 213170 28454
rect 212934 27898 213170 28134
rect 213882 28218 214118 28454
rect 213882 27898 214118 28134
rect 214830 28218 215066 28454
rect 214830 27898 215066 28134
rect 226132 28218 226368 28454
rect 226132 27898 226368 28134
rect 233078 28218 233314 28454
rect 233078 27898 233314 28134
rect 240024 28218 240260 28454
rect 240024 27898 240260 28134
rect 246970 28218 247206 28454
rect 246970 27898 247206 28134
rect 253134 28218 253370 28454
rect 253134 27898 253370 28134
rect 254082 28218 254318 28454
rect 254082 27898 254318 28134
rect 255030 28218 255266 28454
rect 255030 27898 255266 28134
rect 266332 28218 266568 28454
rect 266332 27898 266568 28134
rect 273278 28218 273514 28454
rect 273278 27898 273514 28134
rect 280224 28218 280460 28454
rect 280224 27898 280460 28134
rect 287170 28218 287406 28454
rect 287170 27898 287406 28134
rect 290026 28218 290262 28454
rect 290346 28218 290582 28454
rect 290026 27898 290262 28134
rect 290346 27898 290582 28134
rect 209746 -582 209982 -346
rect 210066 -582 210302 -346
rect 209746 -902 209982 -666
rect 210066 -902 210302 -666
rect 290026 -1542 290262 -1306
rect 290346 -1542 290582 -1306
rect 290026 -1862 290262 -1626
rect 290346 -1862 290582 -1626
rect 293746 704602 293982 704838
rect 294066 704602 294302 704838
rect 293746 704282 293982 704518
rect 294066 704282 294302 704518
rect 293746 697938 293982 698174
rect 294066 697938 294302 698174
rect 293746 697618 293982 697854
rect 294066 697618 294302 697854
rect 293746 660938 293982 661174
rect 294066 660938 294302 661174
rect 293746 660618 293982 660854
rect 294066 660618 294302 660854
rect 293746 623938 293982 624174
rect 294066 623938 294302 624174
rect 293746 623618 293982 623854
rect 294066 623618 294302 623854
rect 293746 586938 293982 587174
rect 294066 586938 294302 587174
rect 293746 586618 293982 586854
rect 294066 586618 294302 586854
rect 293746 549938 293982 550174
rect 294066 549938 294302 550174
rect 293746 549618 293982 549854
rect 294066 549618 294302 549854
rect 293746 512938 293982 513174
rect 294066 512938 294302 513174
rect 293746 512618 293982 512854
rect 294066 512618 294302 512854
rect 293746 475938 293982 476174
rect 294066 475938 294302 476174
rect 293746 475618 293982 475854
rect 294066 475618 294302 475854
rect 293746 438938 293982 439174
rect 294066 438938 294302 439174
rect 293746 438618 293982 438854
rect 294066 438618 294302 438854
rect 293746 401938 293982 402174
rect 294066 401938 294302 402174
rect 293746 401618 293982 401854
rect 294066 401618 294302 401854
rect 293746 364938 293982 365174
rect 294066 364938 294302 365174
rect 293746 364618 293982 364854
rect 294066 364618 294302 364854
rect 293746 327938 293982 328174
rect 294066 327938 294302 328174
rect 293746 327618 293982 327854
rect 294066 327618 294302 327854
rect 293746 290938 293982 291174
rect 294066 290938 294302 291174
rect 293746 290618 293982 290854
rect 294066 290618 294302 290854
rect 293746 253938 293982 254174
rect 294066 253938 294302 254174
rect 293746 253618 293982 253854
rect 294066 253618 294302 253854
rect 293746 216938 293982 217174
rect 294066 216938 294302 217174
rect 293746 216618 293982 216854
rect 294066 216618 294302 216854
rect 293746 179938 293982 180174
rect 294066 179938 294302 180174
rect 293746 179618 293982 179854
rect 294066 179618 294302 179854
rect 293746 142938 293982 143174
rect 294066 142938 294302 143174
rect 293746 142618 293982 142854
rect 294066 142618 294302 142854
rect 293746 105938 293982 106174
rect 294066 105938 294302 106174
rect 293746 105618 293982 105854
rect 294066 105618 294302 105854
rect 293746 68938 293982 69174
rect 294066 68938 294302 69174
rect 293746 68618 293982 68854
rect 294066 68618 294302 68854
rect 293746 31938 293982 32174
rect 294066 31938 294302 32174
rect 293746 31618 293982 31854
rect 294066 31618 294302 31854
rect 293746 -582 293982 -346
rect 294066 -582 294302 -346
rect 293746 -902 293982 -666
rect 294066 -902 294302 -666
rect 318026 705562 318262 705798
rect 318346 705562 318582 705798
rect 318026 705242 318262 705478
rect 318346 705242 318582 705478
rect 318026 694218 318262 694454
rect 318346 694218 318582 694454
rect 318026 693898 318262 694134
rect 318346 693898 318582 694134
rect 318026 657218 318262 657454
rect 318346 657218 318582 657454
rect 318026 656898 318262 657134
rect 318346 656898 318582 657134
rect 318026 620218 318262 620454
rect 318346 620218 318582 620454
rect 318026 619898 318262 620134
rect 318346 619898 318582 620134
rect 318026 583218 318262 583454
rect 318346 583218 318582 583454
rect 318026 582898 318262 583134
rect 318346 582898 318582 583134
rect 318026 546218 318262 546454
rect 318346 546218 318582 546454
rect 318026 545898 318262 546134
rect 318346 545898 318582 546134
rect 318026 509218 318262 509454
rect 318346 509218 318582 509454
rect 318026 508898 318262 509134
rect 318346 508898 318582 509134
rect 318026 472218 318262 472454
rect 318346 472218 318582 472454
rect 318026 471898 318262 472134
rect 318346 471898 318582 472134
rect 318026 435218 318262 435454
rect 318346 435218 318582 435454
rect 318026 434898 318262 435134
rect 318346 434898 318582 435134
rect 318026 398218 318262 398454
rect 318346 398218 318582 398454
rect 318026 397898 318262 398134
rect 318346 397898 318582 398134
rect 318026 361218 318262 361454
rect 318346 361218 318582 361454
rect 318026 360898 318262 361134
rect 318346 360898 318582 361134
rect 318026 324218 318262 324454
rect 318346 324218 318582 324454
rect 318026 323898 318262 324134
rect 318346 323898 318582 324134
rect 318026 287218 318262 287454
rect 318346 287218 318582 287454
rect 318026 286898 318262 287134
rect 318346 286898 318582 287134
rect 318026 250218 318262 250454
rect 318346 250218 318582 250454
rect 318026 249898 318262 250134
rect 318346 249898 318582 250134
rect 318026 213218 318262 213454
rect 318346 213218 318582 213454
rect 318026 212898 318262 213134
rect 318346 212898 318582 213134
rect 318026 176218 318262 176454
rect 318346 176218 318582 176454
rect 318026 175898 318262 176134
rect 318346 175898 318582 176134
rect 318026 139218 318262 139454
rect 318346 139218 318582 139454
rect 318026 138898 318262 139134
rect 318346 138898 318582 139134
rect 318026 102218 318262 102454
rect 318346 102218 318582 102454
rect 318026 101898 318262 102134
rect 318346 101898 318582 102134
rect 318026 65218 318262 65454
rect 318346 65218 318582 65454
rect 318026 64898 318262 65134
rect 318346 64898 318582 65134
rect 318026 28218 318262 28454
rect 318346 28218 318582 28454
rect 318026 27898 318262 28134
rect 318346 27898 318582 28134
rect 318026 -1542 318262 -1306
rect 318346 -1542 318582 -1306
rect 318026 -1862 318262 -1626
rect 318346 -1862 318582 -1626
rect 321746 704602 321982 704838
rect 322066 704602 322302 704838
rect 321746 704282 321982 704518
rect 322066 704282 322302 704518
rect 321746 697938 321982 698174
rect 322066 697938 322302 698174
rect 321746 697618 321982 697854
rect 322066 697618 322302 697854
rect 321746 660938 321982 661174
rect 322066 660938 322302 661174
rect 321746 660618 321982 660854
rect 322066 660618 322302 660854
rect 321746 623938 321982 624174
rect 322066 623938 322302 624174
rect 321746 623618 321982 623854
rect 322066 623618 322302 623854
rect 321746 586938 321982 587174
rect 322066 586938 322302 587174
rect 321746 586618 321982 586854
rect 322066 586618 322302 586854
rect 321746 549938 321982 550174
rect 322066 549938 322302 550174
rect 321746 549618 321982 549854
rect 322066 549618 322302 549854
rect 321746 512938 321982 513174
rect 322066 512938 322302 513174
rect 321746 512618 321982 512854
rect 322066 512618 322302 512854
rect 321746 475938 321982 476174
rect 322066 475938 322302 476174
rect 321746 475618 321982 475854
rect 322066 475618 322302 475854
rect 321746 438938 321982 439174
rect 322066 438938 322302 439174
rect 321746 438618 321982 438854
rect 322066 438618 322302 438854
rect 321746 401938 321982 402174
rect 322066 401938 322302 402174
rect 321746 401618 321982 401854
rect 322066 401618 322302 401854
rect 321746 364938 321982 365174
rect 322066 364938 322302 365174
rect 321746 364618 321982 364854
rect 322066 364618 322302 364854
rect 321746 327938 321982 328174
rect 322066 327938 322302 328174
rect 321746 327618 321982 327854
rect 322066 327618 322302 327854
rect 321746 290938 321982 291174
rect 322066 290938 322302 291174
rect 321746 290618 321982 290854
rect 322066 290618 322302 290854
rect 321746 253938 321982 254174
rect 322066 253938 322302 254174
rect 321746 253618 321982 253854
rect 322066 253618 322302 253854
rect 321746 216938 321982 217174
rect 322066 216938 322302 217174
rect 321746 216618 321982 216854
rect 322066 216618 322302 216854
rect 321746 179938 321982 180174
rect 322066 179938 322302 180174
rect 321746 179618 321982 179854
rect 322066 179618 322302 179854
rect 321746 142938 321982 143174
rect 322066 142938 322302 143174
rect 321746 142618 321982 142854
rect 322066 142618 322302 142854
rect 321746 105938 321982 106174
rect 322066 105938 322302 106174
rect 321746 105618 321982 105854
rect 322066 105618 322302 105854
rect 321746 68938 321982 69174
rect 322066 68938 322302 69174
rect 321746 68618 321982 68854
rect 322066 68618 322302 68854
rect 321746 31938 321982 32174
rect 322066 31938 322302 32174
rect 321746 31618 321982 31854
rect 322066 31618 322302 31854
rect 321746 -582 321982 -346
rect 322066 -582 322302 -346
rect 321746 -902 321982 -666
rect 322066 -902 322302 -666
rect 346026 705562 346262 705798
rect 346346 705562 346582 705798
rect 346026 705242 346262 705478
rect 346346 705242 346582 705478
rect 346026 694218 346262 694454
rect 346346 694218 346582 694454
rect 346026 693898 346262 694134
rect 346346 693898 346582 694134
rect 346026 657218 346262 657454
rect 346346 657218 346582 657454
rect 346026 656898 346262 657134
rect 346346 656898 346582 657134
rect 346026 620218 346262 620454
rect 346346 620218 346582 620454
rect 346026 619898 346262 620134
rect 346346 619898 346582 620134
rect 346026 583218 346262 583454
rect 346346 583218 346582 583454
rect 346026 582898 346262 583134
rect 346346 582898 346582 583134
rect 346026 546218 346262 546454
rect 346346 546218 346582 546454
rect 346026 545898 346262 546134
rect 346346 545898 346582 546134
rect 346026 509218 346262 509454
rect 346346 509218 346582 509454
rect 346026 508898 346262 509134
rect 346346 508898 346582 509134
rect 346026 472218 346262 472454
rect 346346 472218 346582 472454
rect 346026 471898 346262 472134
rect 346346 471898 346582 472134
rect 346026 435218 346262 435454
rect 346346 435218 346582 435454
rect 346026 434898 346262 435134
rect 346346 434898 346582 435134
rect 346026 398218 346262 398454
rect 346346 398218 346582 398454
rect 346026 397898 346262 398134
rect 346346 397898 346582 398134
rect 346026 361218 346262 361454
rect 346346 361218 346582 361454
rect 346026 360898 346262 361134
rect 346346 360898 346582 361134
rect 346026 324218 346262 324454
rect 346346 324218 346582 324454
rect 346026 323898 346262 324134
rect 346346 323898 346582 324134
rect 346026 287218 346262 287454
rect 346346 287218 346582 287454
rect 346026 286898 346262 287134
rect 346346 286898 346582 287134
rect 346026 250218 346262 250454
rect 346346 250218 346582 250454
rect 346026 249898 346262 250134
rect 346346 249898 346582 250134
rect 346026 213218 346262 213454
rect 346346 213218 346582 213454
rect 346026 212898 346262 213134
rect 346346 212898 346582 213134
rect 346026 176218 346262 176454
rect 346346 176218 346582 176454
rect 346026 175898 346262 176134
rect 346346 175898 346582 176134
rect 346026 139218 346262 139454
rect 346346 139218 346582 139454
rect 346026 138898 346262 139134
rect 346346 138898 346582 139134
rect 346026 102218 346262 102454
rect 346346 102218 346582 102454
rect 346026 101898 346262 102134
rect 346346 101898 346582 102134
rect 346026 65218 346262 65454
rect 346346 65218 346582 65454
rect 346026 64898 346262 65134
rect 346346 64898 346582 65134
rect 346026 28218 346262 28454
rect 346346 28218 346582 28454
rect 346026 27898 346262 28134
rect 346346 27898 346582 28134
rect 346026 -1542 346262 -1306
rect 346346 -1542 346582 -1306
rect 346026 -1862 346262 -1626
rect 346346 -1862 346582 -1626
rect 349746 704602 349982 704838
rect 350066 704602 350302 704838
rect 349746 704282 349982 704518
rect 350066 704282 350302 704518
rect 349746 697938 349982 698174
rect 350066 697938 350302 698174
rect 349746 697618 349982 697854
rect 350066 697618 350302 697854
rect 349746 660938 349982 661174
rect 350066 660938 350302 661174
rect 349746 660618 349982 660854
rect 350066 660618 350302 660854
rect 349746 623938 349982 624174
rect 350066 623938 350302 624174
rect 349746 623618 349982 623854
rect 350066 623618 350302 623854
rect 349746 586938 349982 587174
rect 350066 586938 350302 587174
rect 349746 586618 349982 586854
rect 350066 586618 350302 586854
rect 349746 549938 349982 550174
rect 350066 549938 350302 550174
rect 349746 549618 349982 549854
rect 350066 549618 350302 549854
rect 349746 512938 349982 513174
rect 350066 512938 350302 513174
rect 349746 512618 349982 512854
rect 350066 512618 350302 512854
rect 349746 475938 349982 476174
rect 350066 475938 350302 476174
rect 349746 475618 349982 475854
rect 350066 475618 350302 475854
rect 349746 438938 349982 439174
rect 350066 438938 350302 439174
rect 349746 438618 349982 438854
rect 350066 438618 350302 438854
rect 349746 401938 349982 402174
rect 350066 401938 350302 402174
rect 349746 401618 349982 401854
rect 350066 401618 350302 401854
rect 349746 364938 349982 365174
rect 350066 364938 350302 365174
rect 349746 364618 349982 364854
rect 350066 364618 350302 364854
rect 349746 327938 349982 328174
rect 350066 327938 350302 328174
rect 349746 327618 349982 327854
rect 350066 327618 350302 327854
rect 349746 290938 349982 291174
rect 350066 290938 350302 291174
rect 349746 290618 349982 290854
rect 350066 290618 350302 290854
rect 349746 253938 349982 254174
rect 350066 253938 350302 254174
rect 349746 253618 349982 253854
rect 350066 253618 350302 253854
rect 349746 216938 349982 217174
rect 350066 216938 350302 217174
rect 349746 216618 349982 216854
rect 350066 216618 350302 216854
rect 349746 179938 349982 180174
rect 350066 179938 350302 180174
rect 349746 179618 349982 179854
rect 350066 179618 350302 179854
rect 349746 142938 349982 143174
rect 350066 142938 350302 143174
rect 349746 142618 349982 142854
rect 350066 142618 350302 142854
rect 349746 105938 349982 106174
rect 350066 105938 350302 106174
rect 349746 105618 349982 105854
rect 350066 105618 350302 105854
rect 349746 68938 349982 69174
rect 350066 68938 350302 69174
rect 349746 68618 349982 68854
rect 350066 68618 350302 68854
rect 349746 31938 349982 32174
rect 350066 31938 350302 32174
rect 349746 31618 349982 31854
rect 350066 31618 350302 31854
rect 349746 -582 349982 -346
rect 350066 -582 350302 -346
rect 349746 -902 349982 -666
rect 350066 -902 350302 -666
rect 374026 705562 374262 705798
rect 374346 705562 374582 705798
rect 374026 705242 374262 705478
rect 374346 705242 374582 705478
rect 374026 694218 374262 694454
rect 374346 694218 374582 694454
rect 374026 693898 374262 694134
rect 374346 693898 374582 694134
rect 374026 657218 374262 657454
rect 374346 657218 374582 657454
rect 374026 656898 374262 657134
rect 374346 656898 374582 657134
rect 374026 620218 374262 620454
rect 374346 620218 374582 620454
rect 374026 619898 374262 620134
rect 374346 619898 374582 620134
rect 374026 583218 374262 583454
rect 374346 583218 374582 583454
rect 374026 582898 374262 583134
rect 374346 582898 374582 583134
rect 374026 546218 374262 546454
rect 374346 546218 374582 546454
rect 374026 545898 374262 546134
rect 374346 545898 374582 546134
rect 374026 509218 374262 509454
rect 374346 509218 374582 509454
rect 374026 508898 374262 509134
rect 374346 508898 374582 509134
rect 374026 472218 374262 472454
rect 374346 472218 374582 472454
rect 374026 471898 374262 472134
rect 374346 471898 374582 472134
rect 374026 435218 374262 435454
rect 374346 435218 374582 435454
rect 374026 434898 374262 435134
rect 374346 434898 374582 435134
rect 374026 398218 374262 398454
rect 374346 398218 374582 398454
rect 374026 397898 374262 398134
rect 374346 397898 374582 398134
rect 374026 361218 374262 361454
rect 374346 361218 374582 361454
rect 374026 360898 374262 361134
rect 374346 360898 374582 361134
rect 374026 324218 374262 324454
rect 374346 324218 374582 324454
rect 374026 323898 374262 324134
rect 374346 323898 374582 324134
rect 374026 287218 374262 287454
rect 374346 287218 374582 287454
rect 374026 286898 374262 287134
rect 374346 286898 374582 287134
rect 374026 250218 374262 250454
rect 374346 250218 374582 250454
rect 374026 249898 374262 250134
rect 374346 249898 374582 250134
rect 374026 213218 374262 213454
rect 374346 213218 374582 213454
rect 374026 212898 374262 213134
rect 374346 212898 374582 213134
rect 374026 176218 374262 176454
rect 374346 176218 374582 176454
rect 374026 175898 374262 176134
rect 374346 175898 374582 176134
rect 374026 139218 374262 139454
rect 374346 139218 374582 139454
rect 374026 138898 374262 139134
rect 374346 138898 374582 139134
rect 374026 102218 374262 102454
rect 374346 102218 374582 102454
rect 374026 101898 374262 102134
rect 374346 101898 374582 102134
rect 374026 65218 374262 65454
rect 374346 65218 374582 65454
rect 374026 64898 374262 65134
rect 374346 64898 374582 65134
rect 374026 28218 374262 28454
rect 374346 28218 374582 28454
rect 374026 27898 374262 28134
rect 374346 27898 374582 28134
rect 374026 -1542 374262 -1306
rect 374346 -1542 374582 -1306
rect 374026 -1862 374262 -1626
rect 374346 -1862 374582 -1626
rect 377746 704602 377982 704838
rect 378066 704602 378302 704838
rect 377746 704282 377982 704518
rect 378066 704282 378302 704518
rect 377746 697938 377982 698174
rect 378066 697938 378302 698174
rect 377746 697618 377982 697854
rect 378066 697618 378302 697854
rect 377746 660938 377982 661174
rect 378066 660938 378302 661174
rect 377746 660618 377982 660854
rect 378066 660618 378302 660854
rect 377746 623938 377982 624174
rect 378066 623938 378302 624174
rect 377746 623618 377982 623854
rect 378066 623618 378302 623854
rect 377746 586938 377982 587174
rect 378066 586938 378302 587174
rect 377746 586618 377982 586854
rect 378066 586618 378302 586854
rect 377746 549938 377982 550174
rect 378066 549938 378302 550174
rect 377746 549618 377982 549854
rect 378066 549618 378302 549854
rect 377746 512938 377982 513174
rect 378066 512938 378302 513174
rect 377746 512618 377982 512854
rect 378066 512618 378302 512854
rect 377746 475938 377982 476174
rect 378066 475938 378302 476174
rect 377746 475618 377982 475854
rect 378066 475618 378302 475854
rect 377746 438938 377982 439174
rect 378066 438938 378302 439174
rect 377746 438618 377982 438854
rect 378066 438618 378302 438854
rect 377746 401938 377982 402174
rect 378066 401938 378302 402174
rect 377746 401618 377982 401854
rect 378066 401618 378302 401854
rect 377746 364938 377982 365174
rect 378066 364938 378302 365174
rect 377746 364618 377982 364854
rect 378066 364618 378302 364854
rect 377746 327938 377982 328174
rect 378066 327938 378302 328174
rect 377746 327618 377982 327854
rect 378066 327618 378302 327854
rect 377746 290938 377982 291174
rect 378066 290938 378302 291174
rect 377746 290618 377982 290854
rect 378066 290618 378302 290854
rect 377746 253938 377982 254174
rect 378066 253938 378302 254174
rect 377746 253618 377982 253854
rect 378066 253618 378302 253854
rect 377746 216938 377982 217174
rect 378066 216938 378302 217174
rect 377746 216618 377982 216854
rect 378066 216618 378302 216854
rect 377746 179938 377982 180174
rect 378066 179938 378302 180174
rect 377746 179618 377982 179854
rect 378066 179618 378302 179854
rect 377746 142938 377982 143174
rect 378066 142938 378302 143174
rect 377746 142618 377982 142854
rect 378066 142618 378302 142854
rect 377746 105938 377982 106174
rect 378066 105938 378302 106174
rect 377746 105618 377982 105854
rect 378066 105618 378302 105854
rect 377746 68938 377982 69174
rect 378066 68938 378302 69174
rect 377746 68618 377982 68854
rect 378066 68618 378302 68854
rect 377746 31938 377982 32174
rect 378066 31938 378302 32174
rect 377746 31618 377982 31854
rect 378066 31618 378302 31854
rect 377746 -582 377982 -346
rect 378066 -582 378302 -346
rect 377746 -902 377982 -666
rect 378066 -902 378302 -666
rect 402026 705562 402262 705798
rect 402346 705562 402582 705798
rect 402026 705242 402262 705478
rect 402346 705242 402582 705478
rect 402026 694218 402262 694454
rect 402346 694218 402582 694454
rect 402026 693898 402262 694134
rect 402346 693898 402582 694134
rect 402026 657218 402262 657454
rect 402346 657218 402582 657454
rect 402026 656898 402262 657134
rect 402346 656898 402582 657134
rect 402026 620218 402262 620454
rect 402346 620218 402582 620454
rect 402026 619898 402262 620134
rect 402346 619898 402582 620134
rect 402026 583218 402262 583454
rect 402346 583218 402582 583454
rect 402026 582898 402262 583134
rect 402346 582898 402582 583134
rect 402026 546218 402262 546454
rect 402346 546218 402582 546454
rect 402026 545898 402262 546134
rect 402346 545898 402582 546134
rect 402026 509218 402262 509454
rect 402346 509218 402582 509454
rect 402026 508898 402262 509134
rect 402346 508898 402582 509134
rect 402026 472218 402262 472454
rect 402346 472218 402582 472454
rect 402026 471898 402262 472134
rect 402346 471898 402582 472134
rect 402026 435218 402262 435454
rect 402346 435218 402582 435454
rect 402026 434898 402262 435134
rect 402346 434898 402582 435134
rect 402026 398218 402262 398454
rect 402346 398218 402582 398454
rect 402026 397898 402262 398134
rect 402346 397898 402582 398134
rect 402026 361218 402262 361454
rect 402346 361218 402582 361454
rect 402026 360898 402262 361134
rect 402346 360898 402582 361134
rect 402026 324218 402262 324454
rect 402346 324218 402582 324454
rect 402026 323898 402262 324134
rect 402346 323898 402582 324134
rect 402026 287218 402262 287454
rect 402346 287218 402582 287454
rect 402026 286898 402262 287134
rect 402346 286898 402582 287134
rect 402026 250218 402262 250454
rect 402346 250218 402582 250454
rect 402026 249898 402262 250134
rect 402346 249898 402582 250134
rect 402026 213218 402262 213454
rect 402346 213218 402582 213454
rect 402026 212898 402262 213134
rect 402346 212898 402582 213134
rect 402026 176218 402262 176454
rect 402346 176218 402582 176454
rect 402026 175898 402262 176134
rect 402346 175898 402582 176134
rect 402026 139218 402262 139454
rect 402346 139218 402582 139454
rect 402026 138898 402262 139134
rect 402346 138898 402582 139134
rect 402026 102218 402262 102454
rect 402346 102218 402582 102454
rect 402026 101898 402262 102134
rect 402346 101898 402582 102134
rect 402026 65218 402262 65454
rect 402346 65218 402582 65454
rect 402026 64898 402262 65134
rect 402346 64898 402582 65134
rect 402026 28218 402262 28454
rect 402346 28218 402582 28454
rect 402026 27898 402262 28134
rect 402346 27898 402582 28134
rect 402026 -1542 402262 -1306
rect 402346 -1542 402582 -1306
rect 402026 -1862 402262 -1626
rect 402346 -1862 402582 -1626
rect 405746 704602 405982 704838
rect 406066 704602 406302 704838
rect 405746 704282 405982 704518
rect 406066 704282 406302 704518
rect 405746 697938 405982 698174
rect 406066 697938 406302 698174
rect 405746 697618 405982 697854
rect 406066 697618 406302 697854
rect 405746 660938 405982 661174
rect 406066 660938 406302 661174
rect 405746 660618 405982 660854
rect 406066 660618 406302 660854
rect 405746 623938 405982 624174
rect 406066 623938 406302 624174
rect 405746 623618 405982 623854
rect 406066 623618 406302 623854
rect 405746 586938 405982 587174
rect 406066 586938 406302 587174
rect 405746 586618 405982 586854
rect 406066 586618 406302 586854
rect 405746 549938 405982 550174
rect 406066 549938 406302 550174
rect 405746 549618 405982 549854
rect 406066 549618 406302 549854
rect 405746 512938 405982 513174
rect 406066 512938 406302 513174
rect 405746 512618 405982 512854
rect 406066 512618 406302 512854
rect 405746 475938 405982 476174
rect 406066 475938 406302 476174
rect 405746 475618 405982 475854
rect 406066 475618 406302 475854
rect 405746 438938 405982 439174
rect 406066 438938 406302 439174
rect 405746 438618 405982 438854
rect 406066 438618 406302 438854
rect 405746 401938 405982 402174
rect 406066 401938 406302 402174
rect 405746 401618 405982 401854
rect 406066 401618 406302 401854
rect 405746 364938 405982 365174
rect 406066 364938 406302 365174
rect 405746 364618 405982 364854
rect 406066 364618 406302 364854
rect 405746 327938 405982 328174
rect 406066 327938 406302 328174
rect 405746 327618 405982 327854
rect 406066 327618 406302 327854
rect 405746 290938 405982 291174
rect 406066 290938 406302 291174
rect 405746 290618 405982 290854
rect 406066 290618 406302 290854
rect 405746 253938 405982 254174
rect 406066 253938 406302 254174
rect 405746 253618 405982 253854
rect 406066 253618 406302 253854
rect 405746 216938 405982 217174
rect 406066 216938 406302 217174
rect 405746 216618 405982 216854
rect 406066 216618 406302 216854
rect 405746 179938 405982 180174
rect 406066 179938 406302 180174
rect 405746 179618 405982 179854
rect 406066 179618 406302 179854
rect 405746 142938 405982 143174
rect 406066 142938 406302 143174
rect 405746 142618 405982 142854
rect 406066 142618 406302 142854
rect 405746 105938 405982 106174
rect 406066 105938 406302 106174
rect 405746 105618 405982 105854
rect 406066 105618 406302 105854
rect 405746 68938 405982 69174
rect 406066 68938 406302 69174
rect 405746 68618 405982 68854
rect 406066 68618 406302 68854
rect 405746 31938 405982 32174
rect 406066 31938 406302 32174
rect 405746 31618 405982 31854
rect 406066 31618 406302 31854
rect 405746 -582 405982 -346
rect 406066 -582 406302 -346
rect 405746 -902 405982 -666
rect 406066 -902 406302 -666
rect 430026 705562 430262 705798
rect 430346 705562 430582 705798
rect 430026 705242 430262 705478
rect 430346 705242 430582 705478
rect 430026 694218 430262 694454
rect 430346 694218 430582 694454
rect 430026 693898 430262 694134
rect 430346 693898 430582 694134
rect 430026 657218 430262 657454
rect 430346 657218 430582 657454
rect 430026 656898 430262 657134
rect 430346 656898 430582 657134
rect 430026 620218 430262 620454
rect 430346 620218 430582 620454
rect 430026 619898 430262 620134
rect 430346 619898 430582 620134
rect 430026 583218 430262 583454
rect 430346 583218 430582 583454
rect 430026 582898 430262 583134
rect 430346 582898 430582 583134
rect 430026 546218 430262 546454
rect 430346 546218 430582 546454
rect 430026 545898 430262 546134
rect 430346 545898 430582 546134
rect 430026 509218 430262 509454
rect 430346 509218 430582 509454
rect 430026 508898 430262 509134
rect 430346 508898 430582 509134
rect 430026 472218 430262 472454
rect 430346 472218 430582 472454
rect 430026 471898 430262 472134
rect 430346 471898 430582 472134
rect 430026 435218 430262 435454
rect 430346 435218 430582 435454
rect 430026 434898 430262 435134
rect 430346 434898 430582 435134
rect 430026 398218 430262 398454
rect 430346 398218 430582 398454
rect 430026 397898 430262 398134
rect 430346 397898 430582 398134
rect 430026 361218 430262 361454
rect 430346 361218 430582 361454
rect 430026 360898 430262 361134
rect 430346 360898 430582 361134
rect 430026 324218 430262 324454
rect 430346 324218 430582 324454
rect 430026 323898 430262 324134
rect 430346 323898 430582 324134
rect 430026 287218 430262 287454
rect 430346 287218 430582 287454
rect 430026 286898 430262 287134
rect 430346 286898 430582 287134
rect 430026 250218 430262 250454
rect 430346 250218 430582 250454
rect 430026 249898 430262 250134
rect 430346 249898 430582 250134
rect 430026 213218 430262 213454
rect 430346 213218 430582 213454
rect 430026 212898 430262 213134
rect 430346 212898 430582 213134
rect 430026 176218 430262 176454
rect 430346 176218 430582 176454
rect 430026 175898 430262 176134
rect 430346 175898 430582 176134
rect 430026 139218 430262 139454
rect 430346 139218 430582 139454
rect 430026 138898 430262 139134
rect 430346 138898 430582 139134
rect 430026 102218 430262 102454
rect 430346 102218 430582 102454
rect 430026 101898 430262 102134
rect 430346 101898 430582 102134
rect 430026 65218 430262 65454
rect 430346 65218 430582 65454
rect 430026 64898 430262 65134
rect 430346 64898 430582 65134
rect 430026 28218 430262 28454
rect 430346 28218 430582 28454
rect 430026 27898 430262 28134
rect 430346 27898 430582 28134
rect 430026 -1542 430262 -1306
rect 430346 -1542 430582 -1306
rect 430026 -1862 430262 -1626
rect 430346 -1862 430582 -1626
rect 433746 704602 433982 704838
rect 434066 704602 434302 704838
rect 433746 704282 433982 704518
rect 434066 704282 434302 704518
rect 433746 697938 433982 698174
rect 434066 697938 434302 698174
rect 433746 697618 433982 697854
rect 434066 697618 434302 697854
rect 433746 660938 433982 661174
rect 434066 660938 434302 661174
rect 433746 660618 433982 660854
rect 434066 660618 434302 660854
rect 433746 623938 433982 624174
rect 434066 623938 434302 624174
rect 433746 623618 433982 623854
rect 434066 623618 434302 623854
rect 433746 586938 433982 587174
rect 434066 586938 434302 587174
rect 433746 586618 433982 586854
rect 434066 586618 434302 586854
rect 433746 549938 433982 550174
rect 434066 549938 434302 550174
rect 433746 549618 433982 549854
rect 434066 549618 434302 549854
rect 433746 512938 433982 513174
rect 434066 512938 434302 513174
rect 433746 512618 433982 512854
rect 434066 512618 434302 512854
rect 433746 475938 433982 476174
rect 434066 475938 434302 476174
rect 433746 475618 433982 475854
rect 434066 475618 434302 475854
rect 433746 438938 433982 439174
rect 434066 438938 434302 439174
rect 433746 438618 433982 438854
rect 434066 438618 434302 438854
rect 433746 401938 433982 402174
rect 434066 401938 434302 402174
rect 433746 401618 433982 401854
rect 434066 401618 434302 401854
rect 433746 364938 433982 365174
rect 434066 364938 434302 365174
rect 433746 364618 433982 364854
rect 434066 364618 434302 364854
rect 433746 327938 433982 328174
rect 434066 327938 434302 328174
rect 433746 327618 433982 327854
rect 434066 327618 434302 327854
rect 433746 290938 433982 291174
rect 434066 290938 434302 291174
rect 433746 290618 433982 290854
rect 434066 290618 434302 290854
rect 433746 253938 433982 254174
rect 434066 253938 434302 254174
rect 433746 253618 433982 253854
rect 434066 253618 434302 253854
rect 433746 216938 433982 217174
rect 434066 216938 434302 217174
rect 433746 216618 433982 216854
rect 434066 216618 434302 216854
rect 433746 179938 433982 180174
rect 434066 179938 434302 180174
rect 433746 179618 433982 179854
rect 434066 179618 434302 179854
rect 433746 142938 433982 143174
rect 434066 142938 434302 143174
rect 433746 142618 433982 142854
rect 434066 142618 434302 142854
rect 433746 105938 433982 106174
rect 434066 105938 434302 106174
rect 433746 105618 433982 105854
rect 434066 105618 434302 105854
rect 433746 68938 433982 69174
rect 434066 68938 434302 69174
rect 433746 68618 433982 68854
rect 434066 68618 434302 68854
rect 433746 31938 433982 32174
rect 434066 31938 434302 32174
rect 433746 31618 433982 31854
rect 434066 31618 434302 31854
rect 433746 -582 433982 -346
rect 434066 -582 434302 -346
rect 433746 -902 433982 -666
rect 434066 -902 434302 -666
rect 458026 705562 458262 705798
rect 458346 705562 458582 705798
rect 458026 705242 458262 705478
rect 458346 705242 458582 705478
rect 458026 694218 458262 694454
rect 458346 694218 458582 694454
rect 458026 693898 458262 694134
rect 458346 693898 458582 694134
rect 458026 657218 458262 657454
rect 458346 657218 458582 657454
rect 458026 656898 458262 657134
rect 458346 656898 458582 657134
rect 458026 620218 458262 620454
rect 458346 620218 458582 620454
rect 458026 619898 458262 620134
rect 458346 619898 458582 620134
rect 458026 583218 458262 583454
rect 458346 583218 458582 583454
rect 458026 582898 458262 583134
rect 458346 582898 458582 583134
rect 458026 546218 458262 546454
rect 458346 546218 458582 546454
rect 458026 545898 458262 546134
rect 458346 545898 458582 546134
rect 458026 509218 458262 509454
rect 458346 509218 458582 509454
rect 458026 508898 458262 509134
rect 458346 508898 458582 509134
rect 458026 472218 458262 472454
rect 458346 472218 458582 472454
rect 458026 471898 458262 472134
rect 458346 471898 458582 472134
rect 458026 435218 458262 435454
rect 458346 435218 458582 435454
rect 458026 434898 458262 435134
rect 458346 434898 458582 435134
rect 458026 398218 458262 398454
rect 458346 398218 458582 398454
rect 458026 397898 458262 398134
rect 458346 397898 458582 398134
rect 458026 361218 458262 361454
rect 458346 361218 458582 361454
rect 458026 360898 458262 361134
rect 458346 360898 458582 361134
rect 458026 324218 458262 324454
rect 458346 324218 458582 324454
rect 458026 323898 458262 324134
rect 458346 323898 458582 324134
rect 458026 287218 458262 287454
rect 458346 287218 458582 287454
rect 458026 286898 458262 287134
rect 458346 286898 458582 287134
rect 458026 250218 458262 250454
rect 458346 250218 458582 250454
rect 458026 249898 458262 250134
rect 458346 249898 458582 250134
rect 458026 213218 458262 213454
rect 458346 213218 458582 213454
rect 458026 212898 458262 213134
rect 458346 212898 458582 213134
rect 458026 176218 458262 176454
rect 458346 176218 458582 176454
rect 458026 175898 458262 176134
rect 458346 175898 458582 176134
rect 458026 139218 458262 139454
rect 458346 139218 458582 139454
rect 458026 138898 458262 139134
rect 458346 138898 458582 139134
rect 458026 102218 458262 102454
rect 458346 102218 458582 102454
rect 458026 101898 458262 102134
rect 458346 101898 458582 102134
rect 458026 65218 458262 65454
rect 458346 65218 458582 65454
rect 458026 64898 458262 65134
rect 458346 64898 458582 65134
rect 458026 28218 458262 28454
rect 458346 28218 458582 28454
rect 458026 27898 458262 28134
rect 458346 27898 458582 28134
rect 458026 -1542 458262 -1306
rect 458346 -1542 458582 -1306
rect 458026 -1862 458262 -1626
rect 458346 -1862 458582 -1626
rect 461746 704602 461982 704838
rect 462066 704602 462302 704838
rect 461746 704282 461982 704518
rect 462066 704282 462302 704518
rect 461746 697938 461982 698174
rect 462066 697938 462302 698174
rect 461746 697618 461982 697854
rect 462066 697618 462302 697854
rect 461746 660938 461982 661174
rect 462066 660938 462302 661174
rect 461746 660618 461982 660854
rect 462066 660618 462302 660854
rect 461746 623938 461982 624174
rect 462066 623938 462302 624174
rect 461746 623618 461982 623854
rect 462066 623618 462302 623854
rect 461746 586938 461982 587174
rect 462066 586938 462302 587174
rect 461746 586618 461982 586854
rect 462066 586618 462302 586854
rect 461746 549938 461982 550174
rect 462066 549938 462302 550174
rect 461746 549618 461982 549854
rect 462066 549618 462302 549854
rect 461746 512938 461982 513174
rect 462066 512938 462302 513174
rect 461746 512618 461982 512854
rect 462066 512618 462302 512854
rect 461746 475938 461982 476174
rect 462066 475938 462302 476174
rect 461746 475618 461982 475854
rect 462066 475618 462302 475854
rect 461746 438938 461982 439174
rect 462066 438938 462302 439174
rect 461746 438618 461982 438854
rect 462066 438618 462302 438854
rect 461746 401938 461982 402174
rect 462066 401938 462302 402174
rect 461746 401618 461982 401854
rect 462066 401618 462302 401854
rect 461746 364938 461982 365174
rect 462066 364938 462302 365174
rect 461746 364618 461982 364854
rect 462066 364618 462302 364854
rect 461746 327938 461982 328174
rect 462066 327938 462302 328174
rect 461746 327618 461982 327854
rect 462066 327618 462302 327854
rect 461746 290938 461982 291174
rect 462066 290938 462302 291174
rect 461746 290618 461982 290854
rect 462066 290618 462302 290854
rect 461746 253938 461982 254174
rect 462066 253938 462302 254174
rect 461746 253618 461982 253854
rect 462066 253618 462302 253854
rect 461746 216938 461982 217174
rect 462066 216938 462302 217174
rect 461746 216618 461982 216854
rect 462066 216618 462302 216854
rect 461746 179938 461982 180174
rect 462066 179938 462302 180174
rect 461746 179618 461982 179854
rect 462066 179618 462302 179854
rect 461746 142938 461982 143174
rect 462066 142938 462302 143174
rect 461746 142618 461982 142854
rect 462066 142618 462302 142854
rect 461746 105938 461982 106174
rect 462066 105938 462302 106174
rect 461746 105618 461982 105854
rect 462066 105618 462302 105854
rect 461746 68938 461982 69174
rect 462066 68938 462302 69174
rect 461746 68618 461982 68854
rect 462066 68618 462302 68854
rect 461746 31938 461982 32174
rect 462066 31938 462302 32174
rect 461746 31618 461982 31854
rect 462066 31618 462302 31854
rect 461746 -582 461982 -346
rect 462066 -582 462302 -346
rect 461746 -902 461982 -666
rect 462066 -902 462302 -666
rect 486026 705562 486262 705798
rect 486346 705562 486582 705798
rect 486026 705242 486262 705478
rect 486346 705242 486582 705478
rect 486026 694218 486262 694454
rect 486346 694218 486582 694454
rect 486026 693898 486262 694134
rect 486346 693898 486582 694134
rect 486026 657218 486262 657454
rect 486346 657218 486582 657454
rect 486026 656898 486262 657134
rect 486346 656898 486582 657134
rect 486026 620218 486262 620454
rect 486346 620218 486582 620454
rect 486026 619898 486262 620134
rect 486346 619898 486582 620134
rect 486026 583218 486262 583454
rect 486346 583218 486582 583454
rect 486026 582898 486262 583134
rect 486346 582898 486582 583134
rect 486026 546218 486262 546454
rect 486346 546218 486582 546454
rect 486026 545898 486262 546134
rect 486346 545898 486582 546134
rect 486026 509218 486262 509454
rect 486346 509218 486582 509454
rect 486026 508898 486262 509134
rect 486346 508898 486582 509134
rect 486026 472218 486262 472454
rect 486346 472218 486582 472454
rect 486026 471898 486262 472134
rect 486346 471898 486582 472134
rect 486026 435218 486262 435454
rect 486346 435218 486582 435454
rect 486026 434898 486262 435134
rect 486346 434898 486582 435134
rect 486026 398218 486262 398454
rect 486346 398218 486582 398454
rect 486026 397898 486262 398134
rect 486346 397898 486582 398134
rect 486026 361218 486262 361454
rect 486346 361218 486582 361454
rect 486026 360898 486262 361134
rect 486346 360898 486582 361134
rect 486026 324218 486262 324454
rect 486346 324218 486582 324454
rect 486026 323898 486262 324134
rect 486346 323898 486582 324134
rect 486026 287218 486262 287454
rect 486346 287218 486582 287454
rect 486026 286898 486262 287134
rect 486346 286898 486582 287134
rect 486026 250218 486262 250454
rect 486346 250218 486582 250454
rect 486026 249898 486262 250134
rect 486346 249898 486582 250134
rect 486026 213218 486262 213454
rect 486346 213218 486582 213454
rect 486026 212898 486262 213134
rect 486346 212898 486582 213134
rect 486026 176218 486262 176454
rect 486346 176218 486582 176454
rect 486026 175898 486262 176134
rect 486346 175898 486582 176134
rect 486026 139218 486262 139454
rect 486346 139218 486582 139454
rect 486026 138898 486262 139134
rect 486346 138898 486582 139134
rect 486026 102218 486262 102454
rect 486346 102218 486582 102454
rect 486026 101898 486262 102134
rect 486346 101898 486582 102134
rect 486026 65218 486262 65454
rect 486346 65218 486582 65454
rect 486026 64898 486262 65134
rect 486346 64898 486582 65134
rect 486026 28218 486262 28454
rect 486346 28218 486582 28454
rect 486026 27898 486262 28134
rect 486346 27898 486582 28134
rect 486026 -1542 486262 -1306
rect 486346 -1542 486582 -1306
rect 486026 -1862 486262 -1626
rect 486346 -1862 486582 -1626
rect 489746 704602 489982 704838
rect 490066 704602 490302 704838
rect 489746 704282 489982 704518
rect 490066 704282 490302 704518
rect 489746 697938 489982 698174
rect 490066 697938 490302 698174
rect 489746 697618 489982 697854
rect 490066 697618 490302 697854
rect 489746 660938 489982 661174
rect 490066 660938 490302 661174
rect 489746 660618 489982 660854
rect 490066 660618 490302 660854
rect 489746 623938 489982 624174
rect 490066 623938 490302 624174
rect 489746 623618 489982 623854
rect 490066 623618 490302 623854
rect 489746 586938 489982 587174
rect 490066 586938 490302 587174
rect 489746 586618 489982 586854
rect 490066 586618 490302 586854
rect 489746 549938 489982 550174
rect 490066 549938 490302 550174
rect 489746 549618 489982 549854
rect 490066 549618 490302 549854
rect 489746 512938 489982 513174
rect 490066 512938 490302 513174
rect 489746 512618 489982 512854
rect 490066 512618 490302 512854
rect 489746 475938 489982 476174
rect 490066 475938 490302 476174
rect 489746 475618 489982 475854
rect 490066 475618 490302 475854
rect 489746 438938 489982 439174
rect 490066 438938 490302 439174
rect 489746 438618 489982 438854
rect 490066 438618 490302 438854
rect 489746 401938 489982 402174
rect 490066 401938 490302 402174
rect 489746 401618 489982 401854
rect 490066 401618 490302 401854
rect 489746 364938 489982 365174
rect 490066 364938 490302 365174
rect 489746 364618 489982 364854
rect 490066 364618 490302 364854
rect 489746 327938 489982 328174
rect 490066 327938 490302 328174
rect 489746 327618 489982 327854
rect 490066 327618 490302 327854
rect 489746 290938 489982 291174
rect 490066 290938 490302 291174
rect 489746 290618 489982 290854
rect 490066 290618 490302 290854
rect 489746 253938 489982 254174
rect 490066 253938 490302 254174
rect 489746 253618 489982 253854
rect 490066 253618 490302 253854
rect 489746 216938 489982 217174
rect 490066 216938 490302 217174
rect 489746 216618 489982 216854
rect 490066 216618 490302 216854
rect 489746 179938 489982 180174
rect 490066 179938 490302 180174
rect 489746 179618 489982 179854
rect 490066 179618 490302 179854
rect 489746 142938 489982 143174
rect 490066 142938 490302 143174
rect 489746 142618 489982 142854
rect 490066 142618 490302 142854
rect 489746 105938 489982 106174
rect 490066 105938 490302 106174
rect 489746 105618 489982 105854
rect 490066 105618 490302 105854
rect 489746 68938 489982 69174
rect 490066 68938 490302 69174
rect 489746 68618 489982 68854
rect 490066 68618 490302 68854
rect 489746 31938 489982 32174
rect 490066 31938 490302 32174
rect 489746 31618 489982 31854
rect 490066 31618 490302 31854
rect 489746 -582 489982 -346
rect 490066 -582 490302 -346
rect 489746 -902 489982 -666
rect 490066 -902 490302 -666
rect 514026 705562 514262 705798
rect 514346 705562 514582 705798
rect 514026 705242 514262 705478
rect 514346 705242 514582 705478
rect 514026 694218 514262 694454
rect 514346 694218 514582 694454
rect 514026 693898 514262 694134
rect 514346 693898 514582 694134
rect 514026 657218 514262 657454
rect 514346 657218 514582 657454
rect 514026 656898 514262 657134
rect 514346 656898 514582 657134
rect 514026 620218 514262 620454
rect 514346 620218 514582 620454
rect 514026 619898 514262 620134
rect 514346 619898 514582 620134
rect 514026 583218 514262 583454
rect 514346 583218 514582 583454
rect 514026 582898 514262 583134
rect 514346 582898 514582 583134
rect 514026 546218 514262 546454
rect 514346 546218 514582 546454
rect 514026 545898 514262 546134
rect 514346 545898 514582 546134
rect 514026 509218 514262 509454
rect 514346 509218 514582 509454
rect 514026 508898 514262 509134
rect 514346 508898 514582 509134
rect 514026 472218 514262 472454
rect 514346 472218 514582 472454
rect 514026 471898 514262 472134
rect 514346 471898 514582 472134
rect 514026 435218 514262 435454
rect 514346 435218 514582 435454
rect 514026 434898 514262 435134
rect 514346 434898 514582 435134
rect 514026 398218 514262 398454
rect 514346 398218 514582 398454
rect 514026 397898 514262 398134
rect 514346 397898 514582 398134
rect 514026 361218 514262 361454
rect 514346 361218 514582 361454
rect 514026 360898 514262 361134
rect 514346 360898 514582 361134
rect 514026 324218 514262 324454
rect 514346 324218 514582 324454
rect 514026 323898 514262 324134
rect 514346 323898 514582 324134
rect 514026 287218 514262 287454
rect 514346 287218 514582 287454
rect 514026 286898 514262 287134
rect 514346 286898 514582 287134
rect 514026 250218 514262 250454
rect 514346 250218 514582 250454
rect 514026 249898 514262 250134
rect 514346 249898 514582 250134
rect 514026 213218 514262 213454
rect 514346 213218 514582 213454
rect 514026 212898 514262 213134
rect 514346 212898 514582 213134
rect 514026 176218 514262 176454
rect 514346 176218 514582 176454
rect 514026 175898 514262 176134
rect 514346 175898 514582 176134
rect 514026 139218 514262 139454
rect 514346 139218 514582 139454
rect 514026 138898 514262 139134
rect 514346 138898 514582 139134
rect 514026 102218 514262 102454
rect 514346 102218 514582 102454
rect 514026 101898 514262 102134
rect 514346 101898 514582 102134
rect 514026 65218 514262 65454
rect 514346 65218 514582 65454
rect 514026 64898 514262 65134
rect 514346 64898 514582 65134
rect 514026 28218 514262 28454
rect 514346 28218 514582 28454
rect 514026 27898 514262 28134
rect 514346 27898 514582 28134
rect 514026 -1542 514262 -1306
rect 514346 -1542 514582 -1306
rect 514026 -1862 514262 -1626
rect 514346 -1862 514582 -1626
rect 517746 704602 517982 704838
rect 518066 704602 518302 704838
rect 517746 704282 517982 704518
rect 518066 704282 518302 704518
rect 517746 697938 517982 698174
rect 518066 697938 518302 698174
rect 517746 697618 517982 697854
rect 518066 697618 518302 697854
rect 517746 660938 517982 661174
rect 518066 660938 518302 661174
rect 517746 660618 517982 660854
rect 518066 660618 518302 660854
rect 517746 623938 517982 624174
rect 518066 623938 518302 624174
rect 517746 623618 517982 623854
rect 518066 623618 518302 623854
rect 517746 586938 517982 587174
rect 518066 586938 518302 587174
rect 517746 586618 517982 586854
rect 518066 586618 518302 586854
rect 517746 549938 517982 550174
rect 518066 549938 518302 550174
rect 517746 549618 517982 549854
rect 518066 549618 518302 549854
rect 517746 512938 517982 513174
rect 518066 512938 518302 513174
rect 517746 512618 517982 512854
rect 518066 512618 518302 512854
rect 517746 475938 517982 476174
rect 518066 475938 518302 476174
rect 517746 475618 517982 475854
rect 518066 475618 518302 475854
rect 517746 438938 517982 439174
rect 518066 438938 518302 439174
rect 517746 438618 517982 438854
rect 518066 438618 518302 438854
rect 517746 401938 517982 402174
rect 518066 401938 518302 402174
rect 517746 401618 517982 401854
rect 518066 401618 518302 401854
rect 517746 364938 517982 365174
rect 518066 364938 518302 365174
rect 517746 364618 517982 364854
rect 518066 364618 518302 364854
rect 517746 327938 517982 328174
rect 518066 327938 518302 328174
rect 517746 327618 517982 327854
rect 518066 327618 518302 327854
rect 517746 290938 517982 291174
rect 518066 290938 518302 291174
rect 517746 290618 517982 290854
rect 518066 290618 518302 290854
rect 517746 253938 517982 254174
rect 518066 253938 518302 254174
rect 517746 253618 517982 253854
rect 518066 253618 518302 253854
rect 517746 216938 517982 217174
rect 518066 216938 518302 217174
rect 517746 216618 517982 216854
rect 518066 216618 518302 216854
rect 517746 179938 517982 180174
rect 518066 179938 518302 180174
rect 517746 179618 517982 179854
rect 518066 179618 518302 179854
rect 517746 142938 517982 143174
rect 518066 142938 518302 143174
rect 517746 142618 517982 142854
rect 518066 142618 518302 142854
rect 517746 105938 517982 106174
rect 518066 105938 518302 106174
rect 517746 105618 517982 105854
rect 518066 105618 518302 105854
rect 517746 68938 517982 69174
rect 518066 68938 518302 69174
rect 517746 68618 517982 68854
rect 518066 68618 518302 68854
rect 517746 31938 517982 32174
rect 518066 31938 518302 32174
rect 517746 31618 517982 31854
rect 518066 31618 518302 31854
rect 517746 -582 517982 -346
rect 518066 -582 518302 -346
rect 517746 -902 517982 -666
rect 518066 -902 518302 -666
rect 542026 705562 542262 705798
rect 542346 705562 542582 705798
rect 542026 705242 542262 705478
rect 542346 705242 542582 705478
rect 542026 694218 542262 694454
rect 542346 694218 542582 694454
rect 542026 693898 542262 694134
rect 542346 693898 542582 694134
rect 542026 657218 542262 657454
rect 542346 657218 542582 657454
rect 542026 656898 542262 657134
rect 542346 656898 542582 657134
rect 542026 620218 542262 620454
rect 542346 620218 542582 620454
rect 542026 619898 542262 620134
rect 542346 619898 542582 620134
rect 542026 583218 542262 583454
rect 542346 583218 542582 583454
rect 542026 582898 542262 583134
rect 542346 582898 542582 583134
rect 542026 546218 542262 546454
rect 542346 546218 542582 546454
rect 542026 545898 542262 546134
rect 542346 545898 542582 546134
rect 542026 509218 542262 509454
rect 542346 509218 542582 509454
rect 542026 508898 542262 509134
rect 542346 508898 542582 509134
rect 542026 472218 542262 472454
rect 542346 472218 542582 472454
rect 542026 471898 542262 472134
rect 542346 471898 542582 472134
rect 542026 435218 542262 435454
rect 542346 435218 542582 435454
rect 542026 434898 542262 435134
rect 542346 434898 542582 435134
rect 542026 398218 542262 398454
rect 542346 398218 542582 398454
rect 542026 397898 542262 398134
rect 542346 397898 542582 398134
rect 542026 361218 542262 361454
rect 542346 361218 542582 361454
rect 542026 360898 542262 361134
rect 542346 360898 542582 361134
rect 542026 324218 542262 324454
rect 542346 324218 542582 324454
rect 542026 323898 542262 324134
rect 542346 323898 542582 324134
rect 542026 287218 542262 287454
rect 542346 287218 542582 287454
rect 542026 286898 542262 287134
rect 542346 286898 542582 287134
rect 542026 250218 542262 250454
rect 542346 250218 542582 250454
rect 542026 249898 542262 250134
rect 542346 249898 542582 250134
rect 542026 213218 542262 213454
rect 542346 213218 542582 213454
rect 542026 212898 542262 213134
rect 542346 212898 542582 213134
rect 542026 176218 542262 176454
rect 542346 176218 542582 176454
rect 542026 175898 542262 176134
rect 542346 175898 542582 176134
rect 542026 139218 542262 139454
rect 542346 139218 542582 139454
rect 542026 138898 542262 139134
rect 542346 138898 542582 139134
rect 542026 102218 542262 102454
rect 542346 102218 542582 102454
rect 542026 101898 542262 102134
rect 542346 101898 542582 102134
rect 542026 65218 542262 65454
rect 542346 65218 542582 65454
rect 542026 64898 542262 65134
rect 542346 64898 542582 65134
rect 542026 28218 542262 28454
rect 542346 28218 542582 28454
rect 542026 27898 542262 28134
rect 542346 27898 542582 28134
rect 542026 -1542 542262 -1306
rect 542346 -1542 542582 -1306
rect 542026 -1862 542262 -1626
rect 542346 -1862 542582 -1626
rect 545746 704602 545982 704838
rect 546066 704602 546302 704838
rect 545746 704282 545982 704518
rect 546066 704282 546302 704518
rect 545746 697938 545982 698174
rect 546066 697938 546302 698174
rect 545746 697618 545982 697854
rect 546066 697618 546302 697854
rect 545746 660938 545982 661174
rect 546066 660938 546302 661174
rect 545746 660618 545982 660854
rect 546066 660618 546302 660854
rect 545746 623938 545982 624174
rect 546066 623938 546302 624174
rect 545746 623618 545982 623854
rect 546066 623618 546302 623854
rect 545746 586938 545982 587174
rect 546066 586938 546302 587174
rect 545746 586618 545982 586854
rect 546066 586618 546302 586854
rect 545746 549938 545982 550174
rect 546066 549938 546302 550174
rect 545746 549618 545982 549854
rect 546066 549618 546302 549854
rect 545746 512938 545982 513174
rect 546066 512938 546302 513174
rect 545746 512618 545982 512854
rect 546066 512618 546302 512854
rect 545746 475938 545982 476174
rect 546066 475938 546302 476174
rect 545746 475618 545982 475854
rect 546066 475618 546302 475854
rect 545746 438938 545982 439174
rect 546066 438938 546302 439174
rect 545746 438618 545982 438854
rect 546066 438618 546302 438854
rect 545746 401938 545982 402174
rect 546066 401938 546302 402174
rect 545746 401618 545982 401854
rect 546066 401618 546302 401854
rect 545746 364938 545982 365174
rect 546066 364938 546302 365174
rect 545746 364618 545982 364854
rect 546066 364618 546302 364854
rect 545746 327938 545982 328174
rect 546066 327938 546302 328174
rect 545746 327618 545982 327854
rect 546066 327618 546302 327854
rect 545746 290938 545982 291174
rect 546066 290938 546302 291174
rect 545746 290618 545982 290854
rect 546066 290618 546302 290854
rect 545746 253938 545982 254174
rect 546066 253938 546302 254174
rect 545746 253618 545982 253854
rect 546066 253618 546302 253854
rect 545746 216938 545982 217174
rect 546066 216938 546302 217174
rect 545746 216618 545982 216854
rect 546066 216618 546302 216854
rect 545746 179938 545982 180174
rect 546066 179938 546302 180174
rect 545746 179618 545982 179854
rect 546066 179618 546302 179854
rect 545746 142938 545982 143174
rect 546066 142938 546302 143174
rect 545746 142618 545982 142854
rect 546066 142618 546302 142854
rect 545746 105938 545982 106174
rect 546066 105938 546302 106174
rect 545746 105618 545982 105854
rect 546066 105618 546302 105854
rect 545746 68938 545982 69174
rect 546066 68938 546302 69174
rect 545746 68618 545982 68854
rect 546066 68618 546302 68854
rect 545746 31938 545982 32174
rect 546066 31938 546302 32174
rect 545746 31618 545982 31854
rect 546066 31618 546302 31854
rect 545746 -582 545982 -346
rect 546066 -582 546302 -346
rect 545746 -902 545982 -666
rect 546066 -902 546302 -666
rect 570026 705562 570262 705798
rect 570346 705562 570582 705798
rect 570026 705242 570262 705478
rect 570346 705242 570582 705478
rect 570026 694218 570262 694454
rect 570346 694218 570582 694454
rect 570026 693898 570262 694134
rect 570346 693898 570582 694134
rect 570026 657218 570262 657454
rect 570346 657218 570582 657454
rect 570026 656898 570262 657134
rect 570346 656898 570582 657134
rect 570026 620218 570262 620454
rect 570346 620218 570582 620454
rect 570026 619898 570262 620134
rect 570346 619898 570582 620134
rect 570026 583218 570262 583454
rect 570346 583218 570582 583454
rect 570026 582898 570262 583134
rect 570346 582898 570582 583134
rect 570026 546218 570262 546454
rect 570346 546218 570582 546454
rect 570026 545898 570262 546134
rect 570346 545898 570582 546134
rect 570026 509218 570262 509454
rect 570346 509218 570582 509454
rect 570026 508898 570262 509134
rect 570346 508898 570582 509134
rect 570026 472218 570262 472454
rect 570346 472218 570582 472454
rect 570026 471898 570262 472134
rect 570346 471898 570582 472134
rect 570026 435218 570262 435454
rect 570346 435218 570582 435454
rect 570026 434898 570262 435134
rect 570346 434898 570582 435134
rect 570026 398218 570262 398454
rect 570346 398218 570582 398454
rect 570026 397898 570262 398134
rect 570346 397898 570582 398134
rect 570026 361218 570262 361454
rect 570346 361218 570582 361454
rect 570026 360898 570262 361134
rect 570346 360898 570582 361134
rect 570026 324218 570262 324454
rect 570346 324218 570582 324454
rect 570026 323898 570262 324134
rect 570346 323898 570582 324134
rect 570026 287218 570262 287454
rect 570346 287218 570582 287454
rect 570026 286898 570262 287134
rect 570346 286898 570582 287134
rect 570026 250218 570262 250454
rect 570346 250218 570582 250454
rect 570026 249898 570262 250134
rect 570346 249898 570582 250134
rect 570026 213218 570262 213454
rect 570346 213218 570582 213454
rect 570026 212898 570262 213134
rect 570346 212898 570582 213134
rect 570026 176218 570262 176454
rect 570346 176218 570582 176454
rect 570026 175898 570262 176134
rect 570346 175898 570582 176134
rect 570026 139218 570262 139454
rect 570346 139218 570582 139454
rect 570026 138898 570262 139134
rect 570346 138898 570582 139134
rect 570026 102218 570262 102454
rect 570346 102218 570582 102454
rect 570026 101898 570262 102134
rect 570346 101898 570582 102134
rect 570026 65218 570262 65454
rect 570346 65218 570582 65454
rect 570026 64898 570262 65134
rect 570346 64898 570582 65134
rect 570026 28218 570262 28454
rect 570346 28218 570582 28454
rect 570026 27898 570262 28134
rect 570346 27898 570582 28134
rect 570026 -1542 570262 -1306
rect 570346 -1542 570582 -1306
rect 570026 -1862 570262 -1626
rect 570346 -1862 570582 -1626
rect 592062 711322 592298 711558
rect 592382 711322 592618 711558
rect 592062 711002 592298 711238
rect 592382 711002 592618 711238
rect 591102 710362 591338 710598
rect 591422 710362 591658 710598
rect 591102 710042 591338 710278
rect 591422 710042 591658 710278
rect 590142 709402 590378 709638
rect 590462 709402 590698 709638
rect 590142 709082 590378 709318
rect 590462 709082 590698 709318
rect 589182 708442 589418 708678
rect 589502 708442 589738 708678
rect 589182 708122 589418 708358
rect 589502 708122 589738 708358
rect 588222 707482 588458 707718
rect 588542 707482 588778 707718
rect 588222 707162 588458 707398
rect 588542 707162 588778 707398
rect 587262 706522 587498 706758
rect 587582 706522 587818 706758
rect 587262 706202 587498 706438
rect 587582 706202 587818 706438
rect 586302 705562 586538 705798
rect 586622 705562 586858 705798
rect 586302 705242 586538 705478
rect 586622 705242 586858 705478
rect 573746 704602 573982 704838
rect 574066 704602 574302 704838
rect 573746 704282 573982 704518
rect 574066 704282 574302 704518
rect 573746 697938 573982 698174
rect 574066 697938 574302 698174
rect 573746 697618 573982 697854
rect 574066 697618 574302 697854
rect 573746 660938 573982 661174
rect 574066 660938 574302 661174
rect 573746 660618 573982 660854
rect 574066 660618 574302 660854
rect 573746 623938 573982 624174
rect 574066 623938 574302 624174
rect 573746 623618 573982 623854
rect 574066 623618 574302 623854
rect 573746 586938 573982 587174
rect 574066 586938 574302 587174
rect 573746 586618 573982 586854
rect 574066 586618 574302 586854
rect 573746 549938 573982 550174
rect 574066 549938 574302 550174
rect 573746 549618 573982 549854
rect 574066 549618 574302 549854
rect 573746 512938 573982 513174
rect 574066 512938 574302 513174
rect 573746 512618 573982 512854
rect 574066 512618 574302 512854
rect 573746 475938 573982 476174
rect 574066 475938 574302 476174
rect 573746 475618 573982 475854
rect 574066 475618 574302 475854
rect 573746 438938 573982 439174
rect 574066 438938 574302 439174
rect 573746 438618 573982 438854
rect 574066 438618 574302 438854
rect 573746 401938 573982 402174
rect 574066 401938 574302 402174
rect 573746 401618 573982 401854
rect 574066 401618 574302 401854
rect 573746 364938 573982 365174
rect 574066 364938 574302 365174
rect 573746 364618 573982 364854
rect 574066 364618 574302 364854
rect 573746 327938 573982 328174
rect 574066 327938 574302 328174
rect 573746 327618 573982 327854
rect 574066 327618 574302 327854
rect 573746 290938 573982 291174
rect 574066 290938 574302 291174
rect 573746 290618 573982 290854
rect 574066 290618 574302 290854
rect 573746 253938 573982 254174
rect 574066 253938 574302 254174
rect 573746 253618 573982 253854
rect 574066 253618 574302 253854
rect 573746 216938 573982 217174
rect 574066 216938 574302 217174
rect 573746 216618 573982 216854
rect 574066 216618 574302 216854
rect 573746 179938 573982 180174
rect 574066 179938 574302 180174
rect 573746 179618 573982 179854
rect 574066 179618 574302 179854
rect 573746 142938 573982 143174
rect 574066 142938 574302 143174
rect 573746 142618 573982 142854
rect 574066 142618 574302 142854
rect 573746 105938 573982 106174
rect 574066 105938 574302 106174
rect 573746 105618 573982 105854
rect 574066 105618 574302 105854
rect 573746 68938 573982 69174
rect 574066 68938 574302 69174
rect 573746 68618 573982 68854
rect 574066 68618 574302 68854
rect 573746 31938 573982 32174
rect 574066 31938 574302 32174
rect 573746 31618 573982 31854
rect 574066 31618 574302 31854
rect 573746 -582 573982 -346
rect 574066 -582 574302 -346
rect 573746 -902 573982 -666
rect 574066 -902 574302 -666
rect 585342 704602 585578 704838
rect 585662 704602 585898 704838
rect 585342 704282 585578 704518
rect 585662 704282 585898 704518
rect 585342 697938 585578 698174
rect 585662 697938 585898 698174
rect 585342 697618 585578 697854
rect 585662 697618 585898 697854
rect 585342 660938 585578 661174
rect 585662 660938 585898 661174
rect 585342 660618 585578 660854
rect 585662 660618 585898 660854
rect 585342 623938 585578 624174
rect 585662 623938 585898 624174
rect 585342 623618 585578 623854
rect 585662 623618 585898 623854
rect 585342 586938 585578 587174
rect 585662 586938 585898 587174
rect 585342 586618 585578 586854
rect 585662 586618 585898 586854
rect 585342 549938 585578 550174
rect 585662 549938 585898 550174
rect 585342 549618 585578 549854
rect 585662 549618 585898 549854
rect 585342 512938 585578 513174
rect 585662 512938 585898 513174
rect 585342 512618 585578 512854
rect 585662 512618 585898 512854
rect 585342 475938 585578 476174
rect 585662 475938 585898 476174
rect 585342 475618 585578 475854
rect 585662 475618 585898 475854
rect 585342 438938 585578 439174
rect 585662 438938 585898 439174
rect 585342 438618 585578 438854
rect 585662 438618 585898 438854
rect 585342 401938 585578 402174
rect 585662 401938 585898 402174
rect 585342 401618 585578 401854
rect 585662 401618 585898 401854
rect 585342 364938 585578 365174
rect 585662 364938 585898 365174
rect 585342 364618 585578 364854
rect 585662 364618 585898 364854
rect 585342 327938 585578 328174
rect 585662 327938 585898 328174
rect 585342 327618 585578 327854
rect 585662 327618 585898 327854
rect 585342 290938 585578 291174
rect 585662 290938 585898 291174
rect 585342 290618 585578 290854
rect 585662 290618 585898 290854
rect 585342 253938 585578 254174
rect 585662 253938 585898 254174
rect 585342 253618 585578 253854
rect 585662 253618 585898 253854
rect 585342 216938 585578 217174
rect 585662 216938 585898 217174
rect 585342 216618 585578 216854
rect 585662 216618 585898 216854
rect 585342 179938 585578 180174
rect 585662 179938 585898 180174
rect 585342 179618 585578 179854
rect 585662 179618 585898 179854
rect 585342 142938 585578 143174
rect 585662 142938 585898 143174
rect 585342 142618 585578 142854
rect 585662 142618 585898 142854
rect 585342 105938 585578 106174
rect 585662 105938 585898 106174
rect 585342 105618 585578 105854
rect 585662 105618 585898 105854
rect 585342 68938 585578 69174
rect 585662 68938 585898 69174
rect 585342 68618 585578 68854
rect 585662 68618 585898 68854
rect 585342 31938 585578 32174
rect 585662 31938 585898 32174
rect 585342 31618 585578 31854
rect 585662 31618 585898 31854
rect 585342 -582 585578 -346
rect 585662 -582 585898 -346
rect 585342 -902 585578 -666
rect 585662 -902 585898 -666
rect 586302 694218 586538 694454
rect 586622 694218 586858 694454
rect 586302 693898 586538 694134
rect 586622 693898 586858 694134
rect 586302 657218 586538 657454
rect 586622 657218 586858 657454
rect 586302 656898 586538 657134
rect 586622 656898 586858 657134
rect 586302 620218 586538 620454
rect 586622 620218 586858 620454
rect 586302 619898 586538 620134
rect 586622 619898 586858 620134
rect 586302 583218 586538 583454
rect 586622 583218 586858 583454
rect 586302 582898 586538 583134
rect 586622 582898 586858 583134
rect 586302 546218 586538 546454
rect 586622 546218 586858 546454
rect 586302 545898 586538 546134
rect 586622 545898 586858 546134
rect 586302 509218 586538 509454
rect 586622 509218 586858 509454
rect 586302 508898 586538 509134
rect 586622 508898 586858 509134
rect 586302 472218 586538 472454
rect 586622 472218 586858 472454
rect 586302 471898 586538 472134
rect 586622 471898 586858 472134
rect 586302 435218 586538 435454
rect 586622 435218 586858 435454
rect 586302 434898 586538 435134
rect 586622 434898 586858 435134
rect 586302 398218 586538 398454
rect 586622 398218 586858 398454
rect 586302 397898 586538 398134
rect 586622 397898 586858 398134
rect 586302 361218 586538 361454
rect 586622 361218 586858 361454
rect 586302 360898 586538 361134
rect 586622 360898 586858 361134
rect 586302 324218 586538 324454
rect 586622 324218 586858 324454
rect 586302 323898 586538 324134
rect 586622 323898 586858 324134
rect 586302 287218 586538 287454
rect 586622 287218 586858 287454
rect 586302 286898 586538 287134
rect 586622 286898 586858 287134
rect 586302 250218 586538 250454
rect 586622 250218 586858 250454
rect 586302 249898 586538 250134
rect 586622 249898 586858 250134
rect 586302 213218 586538 213454
rect 586622 213218 586858 213454
rect 586302 212898 586538 213134
rect 586622 212898 586858 213134
rect 586302 176218 586538 176454
rect 586622 176218 586858 176454
rect 586302 175898 586538 176134
rect 586622 175898 586858 176134
rect 586302 139218 586538 139454
rect 586622 139218 586858 139454
rect 586302 138898 586538 139134
rect 586622 138898 586858 139134
rect 586302 102218 586538 102454
rect 586622 102218 586858 102454
rect 586302 101898 586538 102134
rect 586622 101898 586858 102134
rect 586302 65218 586538 65454
rect 586622 65218 586858 65454
rect 586302 64898 586538 65134
rect 586622 64898 586858 65134
rect 586302 28218 586538 28454
rect 586622 28218 586858 28454
rect 586302 27898 586538 28134
rect 586622 27898 586858 28134
rect 586302 -1542 586538 -1306
rect 586622 -1542 586858 -1306
rect 586302 -1862 586538 -1626
rect 586622 -1862 586858 -1626
rect 587262 -2502 587498 -2266
rect 587582 -2502 587818 -2266
rect 587262 -2822 587498 -2586
rect 587582 -2822 587818 -2586
rect 588222 -3462 588458 -3226
rect 588542 -3462 588778 -3226
rect 588222 -3782 588458 -3546
rect 588542 -3782 588778 -3546
rect 589182 -4422 589418 -4186
rect 589502 -4422 589738 -4186
rect 589182 -4742 589418 -4506
rect 589502 -4742 589738 -4506
rect 590142 -5382 590378 -5146
rect 590462 -5382 590698 -5146
rect 590142 -5702 590378 -5466
rect 590462 -5702 590698 -5466
rect 591102 -6342 591338 -6106
rect 591422 -6342 591658 -6106
rect 591102 -6662 591338 -6426
rect 591422 -6662 591658 -6426
rect 592062 -7302 592298 -7066
rect 592382 -7302 592618 -7066
rect 592062 -7622 592298 -7386
rect 592382 -7622 592618 -7386
<< metal5 >>
rect -8726 711558 592650 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect -8726 711238 592650 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect -8726 710970 592650 711002
rect -7766 710598 591690 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect -7766 710278 591690 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect -7766 710010 591690 710042
rect -6806 709638 590730 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect -6806 709318 590730 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect -6806 709050 590730 709082
rect -5846 708678 589770 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect -5846 708358 589770 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect -5846 708090 589770 708122
rect -4886 707718 588810 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect -4886 707398 588810 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect -4886 707130 588810 707162
rect -3926 706758 587850 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect -3926 706438 587850 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect -3926 706170 587850 706202
rect -2966 705798 586890 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 38026 705798
rect 38262 705562 38346 705798
rect 38582 705562 66026 705798
rect 66262 705562 66346 705798
rect 66582 705562 94026 705798
rect 94262 705562 94346 705798
rect 94582 705562 122026 705798
rect 122262 705562 122346 705798
rect 122582 705562 150026 705798
rect 150262 705562 150346 705798
rect 150582 705562 178026 705798
rect 178262 705562 178346 705798
rect 178582 705562 206026 705798
rect 206262 705562 206346 705798
rect 206582 705562 234026 705798
rect 234262 705562 234346 705798
rect 234582 705562 262026 705798
rect 262262 705562 262346 705798
rect 262582 705562 290026 705798
rect 290262 705562 290346 705798
rect 290582 705562 318026 705798
rect 318262 705562 318346 705798
rect 318582 705562 346026 705798
rect 346262 705562 346346 705798
rect 346582 705562 374026 705798
rect 374262 705562 374346 705798
rect 374582 705562 402026 705798
rect 402262 705562 402346 705798
rect 402582 705562 430026 705798
rect 430262 705562 430346 705798
rect 430582 705562 458026 705798
rect 458262 705562 458346 705798
rect 458582 705562 486026 705798
rect 486262 705562 486346 705798
rect 486582 705562 514026 705798
rect 514262 705562 514346 705798
rect 514582 705562 542026 705798
rect 542262 705562 542346 705798
rect 542582 705562 570026 705798
rect 570262 705562 570346 705798
rect 570582 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect -2966 705478 586890 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 38026 705478
rect 38262 705242 38346 705478
rect 38582 705242 66026 705478
rect 66262 705242 66346 705478
rect 66582 705242 94026 705478
rect 94262 705242 94346 705478
rect 94582 705242 122026 705478
rect 122262 705242 122346 705478
rect 122582 705242 150026 705478
rect 150262 705242 150346 705478
rect 150582 705242 178026 705478
rect 178262 705242 178346 705478
rect 178582 705242 206026 705478
rect 206262 705242 206346 705478
rect 206582 705242 234026 705478
rect 234262 705242 234346 705478
rect 234582 705242 262026 705478
rect 262262 705242 262346 705478
rect 262582 705242 290026 705478
rect 290262 705242 290346 705478
rect 290582 705242 318026 705478
rect 318262 705242 318346 705478
rect 318582 705242 346026 705478
rect 346262 705242 346346 705478
rect 346582 705242 374026 705478
rect 374262 705242 374346 705478
rect 374582 705242 402026 705478
rect 402262 705242 402346 705478
rect 402582 705242 430026 705478
rect 430262 705242 430346 705478
rect 430582 705242 458026 705478
rect 458262 705242 458346 705478
rect 458582 705242 486026 705478
rect 486262 705242 486346 705478
rect 486582 705242 514026 705478
rect 514262 705242 514346 705478
rect 514582 705242 542026 705478
rect 542262 705242 542346 705478
rect 542582 705242 570026 705478
rect 570262 705242 570346 705478
rect 570582 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect -2966 705210 586890 705242
rect -2006 704838 585930 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 41746 704838
rect 41982 704602 42066 704838
rect 42302 704602 69746 704838
rect 69982 704602 70066 704838
rect 70302 704602 97746 704838
rect 97982 704602 98066 704838
rect 98302 704602 125746 704838
rect 125982 704602 126066 704838
rect 126302 704602 153746 704838
rect 153982 704602 154066 704838
rect 154302 704602 181746 704838
rect 181982 704602 182066 704838
rect 182302 704602 209746 704838
rect 209982 704602 210066 704838
rect 210302 704602 237746 704838
rect 237982 704602 238066 704838
rect 238302 704602 265746 704838
rect 265982 704602 266066 704838
rect 266302 704602 293746 704838
rect 293982 704602 294066 704838
rect 294302 704602 321746 704838
rect 321982 704602 322066 704838
rect 322302 704602 349746 704838
rect 349982 704602 350066 704838
rect 350302 704602 377746 704838
rect 377982 704602 378066 704838
rect 378302 704602 405746 704838
rect 405982 704602 406066 704838
rect 406302 704602 433746 704838
rect 433982 704602 434066 704838
rect 434302 704602 461746 704838
rect 461982 704602 462066 704838
rect 462302 704602 489746 704838
rect 489982 704602 490066 704838
rect 490302 704602 517746 704838
rect 517982 704602 518066 704838
rect 518302 704602 545746 704838
rect 545982 704602 546066 704838
rect 546302 704602 573746 704838
rect 573982 704602 574066 704838
rect 574302 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect -2006 704518 585930 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 41746 704518
rect 41982 704282 42066 704518
rect 42302 704282 69746 704518
rect 69982 704282 70066 704518
rect 70302 704282 97746 704518
rect 97982 704282 98066 704518
rect 98302 704282 125746 704518
rect 125982 704282 126066 704518
rect 126302 704282 153746 704518
rect 153982 704282 154066 704518
rect 154302 704282 181746 704518
rect 181982 704282 182066 704518
rect 182302 704282 209746 704518
rect 209982 704282 210066 704518
rect 210302 704282 237746 704518
rect 237982 704282 238066 704518
rect 238302 704282 265746 704518
rect 265982 704282 266066 704518
rect 266302 704282 293746 704518
rect 293982 704282 294066 704518
rect 294302 704282 321746 704518
rect 321982 704282 322066 704518
rect 322302 704282 349746 704518
rect 349982 704282 350066 704518
rect 350302 704282 377746 704518
rect 377982 704282 378066 704518
rect 378302 704282 405746 704518
rect 405982 704282 406066 704518
rect 406302 704282 433746 704518
rect 433982 704282 434066 704518
rect 434302 704282 461746 704518
rect 461982 704282 462066 704518
rect 462302 704282 489746 704518
rect 489982 704282 490066 704518
rect 490302 704282 517746 704518
rect 517982 704282 518066 704518
rect 518302 704282 545746 704518
rect 545982 704282 546066 704518
rect 546302 704282 573746 704518
rect 573982 704282 574066 704518
rect 574302 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect -2006 704250 585930 704282
rect -8726 698174 592650 698206
rect -8726 697938 -1974 698174
rect -1738 697938 -1654 698174
rect -1418 697938 41746 698174
rect 41982 697938 42066 698174
rect 42302 697938 69746 698174
rect 69982 697938 70066 698174
rect 70302 697938 97746 698174
rect 97982 697938 98066 698174
rect 98302 697938 125746 698174
rect 125982 697938 126066 698174
rect 126302 697938 153746 698174
rect 153982 697938 154066 698174
rect 154302 697938 181746 698174
rect 181982 697938 182066 698174
rect 182302 697938 209746 698174
rect 209982 697938 210066 698174
rect 210302 697938 237746 698174
rect 237982 697938 238066 698174
rect 238302 697938 265746 698174
rect 265982 697938 266066 698174
rect 266302 697938 293746 698174
rect 293982 697938 294066 698174
rect 294302 697938 321746 698174
rect 321982 697938 322066 698174
rect 322302 697938 349746 698174
rect 349982 697938 350066 698174
rect 350302 697938 377746 698174
rect 377982 697938 378066 698174
rect 378302 697938 405746 698174
rect 405982 697938 406066 698174
rect 406302 697938 433746 698174
rect 433982 697938 434066 698174
rect 434302 697938 461746 698174
rect 461982 697938 462066 698174
rect 462302 697938 489746 698174
rect 489982 697938 490066 698174
rect 490302 697938 517746 698174
rect 517982 697938 518066 698174
rect 518302 697938 545746 698174
rect 545982 697938 546066 698174
rect 546302 697938 573746 698174
rect 573982 697938 574066 698174
rect 574302 697938 585342 698174
rect 585578 697938 585662 698174
rect 585898 697938 592650 698174
rect -8726 697854 592650 697938
rect -8726 697618 -1974 697854
rect -1738 697618 -1654 697854
rect -1418 697618 41746 697854
rect 41982 697618 42066 697854
rect 42302 697618 69746 697854
rect 69982 697618 70066 697854
rect 70302 697618 97746 697854
rect 97982 697618 98066 697854
rect 98302 697618 125746 697854
rect 125982 697618 126066 697854
rect 126302 697618 153746 697854
rect 153982 697618 154066 697854
rect 154302 697618 181746 697854
rect 181982 697618 182066 697854
rect 182302 697618 209746 697854
rect 209982 697618 210066 697854
rect 210302 697618 237746 697854
rect 237982 697618 238066 697854
rect 238302 697618 265746 697854
rect 265982 697618 266066 697854
rect 266302 697618 293746 697854
rect 293982 697618 294066 697854
rect 294302 697618 321746 697854
rect 321982 697618 322066 697854
rect 322302 697618 349746 697854
rect 349982 697618 350066 697854
rect 350302 697618 377746 697854
rect 377982 697618 378066 697854
rect 378302 697618 405746 697854
rect 405982 697618 406066 697854
rect 406302 697618 433746 697854
rect 433982 697618 434066 697854
rect 434302 697618 461746 697854
rect 461982 697618 462066 697854
rect 462302 697618 489746 697854
rect 489982 697618 490066 697854
rect 490302 697618 517746 697854
rect 517982 697618 518066 697854
rect 518302 697618 545746 697854
rect 545982 697618 546066 697854
rect 546302 697618 573746 697854
rect 573982 697618 574066 697854
rect 574302 697618 585342 697854
rect 585578 697618 585662 697854
rect 585898 697618 592650 697854
rect -8726 697586 592650 697618
rect -8726 694454 592650 694486
rect -8726 694218 -2934 694454
rect -2698 694218 -2614 694454
rect -2378 694218 38026 694454
rect 38262 694218 38346 694454
rect 38582 694218 66026 694454
rect 66262 694218 66346 694454
rect 66582 694218 94026 694454
rect 94262 694218 94346 694454
rect 94582 694218 122026 694454
rect 122262 694218 122346 694454
rect 122582 694218 150026 694454
rect 150262 694218 150346 694454
rect 150582 694218 178026 694454
rect 178262 694218 178346 694454
rect 178582 694218 206026 694454
rect 206262 694218 206346 694454
rect 206582 694218 234026 694454
rect 234262 694218 234346 694454
rect 234582 694218 262026 694454
rect 262262 694218 262346 694454
rect 262582 694218 290026 694454
rect 290262 694218 290346 694454
rect 290582 694218 318026 694454
rect 318262 694218 318346 694454
rect 318582 694218 346026 694454
rect 346262 694218 346346 694454
rect 346582 694218 374026 694454
rect 374262 694218 374346 694454
rect 374582 694218 402026 694454
rect 402262 694218 402346 694454
rect 402582 694218 430026 694454
rect 430262 694218 430346 694454
rect 430582 694218 458026 694454
rect 458262 694218 458346 694454
rect 458582 694218 486026 694454
rect 486262 694218 486346 694454
rect 486582 694218 514026 694454
rect 514262 694218 514346 694454
rect 514582 694218 542026 694454
rect 542262 694218 542346 694454
rect 542582 694218 570026 694454
rect 570262 694218 570346 694454
rect 570582 694218 586302 694454
rect 586538 694218 586622 694454
rect 586858 694218 592650 694454
rect -8726 694134 592650 694218
rect -8726 693898 -2934 694134
rect -2698 693898 -2614 694134
rect -2378 693898 38026 694134
rect 38262 693898 38346 694134
rect 38582 693898 66026 694134
rect 66262 693898 66346 694134
rect 66582 693898 94026 694134
rect 94262 693898 94346 694134
rect 94582 693898 122026 694134
rect 122262 693898 122346 694134
rect 122582 693898 150026 694134
rect 150262 693898 150346 694134
rect 150582 693898 178026 694134
rect 178262 693898 178346 694134
rect 178582 693898 206026 694134
rect 206262 693898 206346 694134
rect 206582 693898 234026 694134
rect 234262 693898 234346 694134
rect 234582 693898 262026 694134
rect 262262 693898 262346 694134
rect 262582 693898 290026 694134
rect 290262 693898 290346 694134
rect 290582 693898 318026 694134
rect 318262 693898 318346 694134
rect 318582 693898 346026 694134
rect 346262 693898 346346 694134
rect 346582 693898 374026 694134
rect 374262 693898 374346 694134
rect 374582 693898 402026 694134
rect 402262 693898 402346 694134
rect 402582 693898 430026 694134
rect 430262 693898 430346 694134
rect 430582 693898 458026 694134
rect 458262 693898 458346 694134
rect 458582 693898 486026 694134
rect 486262 693898 486346 694134
rect 486582 693898 514026 694134
rect 514262 693898 514346 694134
rect 514582 693898 542026 694134
rect 542262 693898 542346 694134
rect 542582 693898 570026 694134
rect 570262 693898 570346 694134
rect 570582 693898 586302 694134
rect 586538 693898 586622 694134
rect 586858 693898 592650 694134
rect -8726 693866 592650 693898
rect -8726 661174 592650 661206
rect -8726 660938 -1974 661174
rect -1738 660938 -1654 661174
rect -1418 660938 41746 661174
rect 41982 660938 42066 661174
rect 42302 660938 69746 661174
rect 69982 660938 70066 661174
rect 70302 660938 97746 661174
rect 97982 660938 98066 661174
rect 98302 660938 125746 661174
rect 125982 660938 126066 661174
rect 126302 660938 153746 661174
rect 153982 660938 154066 661174
rect 154302 660938 181746 661174
rect 181982 660938 182066 661174
rect 182302 660938 209746 661174
rect 209982 660938 210066 661174
rect 210302 660938 237746 661174
rect 237982 660938 238066 661174
rect 238302 660938 265746 661174
rect 265982 660938 266066 661174
rect 266302 660938 293746 661174
rect 293982 660938 294066 661174
rect 294302 660938 321746 661174
rect 321982 660938 322066 661174
rect 322302 660938 349746 661174
rect 349982 660938 350066 661174
rect 350302 660938 377746 661174
rect 377982 660938 378066 661174
rect 378302 660938 405746 661174
rect 405982 660938 406066 661174
rect 406302 660938 433746 661174
rect 433982 660938 434066 661174
rect 434302 660938 461746 661174
rect 461982 660938 462066 661174
rect 462302 660938 489746 661174
rect 489982 660938 490066 661174
rect 490302 660938 517746 661174
rect 517982 660938 518066 661174
rect 518302 660938 545746 661174
rect 545982 660938 546066 661174
rect 546302 660938 573746 661174
rect 573982 660938 574066 661174
rect 574302 660938 585342 661174
rect 585578 660938 585662 661174
rect 585898 660938 592650 661174
rect -8726 660854 592650 660938
rect -8726 660618 -1974 660854
rect -1738 660618 -1654 660854
rect -1418 660618 41746 660854
rect 41982 660618 42066 660854
rect 42302 660618 69746 660854
rect 69982 660618 70066 660854
rect 70302 660618 97746 660854
rect 97982 660618 98066 660854
rect 98302 660618 125746 660854
rect 125982 660618 126066 660854
rect 126302 660618 153746 660854
rect 153982 660618 154066 660854
rect 154302 660618 181746 660854
rect 181982 660618 182066 660854
rect 182302 660618 209746 660854
rect 209982 660618 210066 660854
rect 210302 660618 237746 660854
rect 237982 660618 238066 660854
rect 238302 660618 265746 660854
rect 265982 660618 266066 660854
rect 266302 660618 293746 660854
rect 293982 660618 294066 660854
rect 294302 660618 321746 660854
rect 321982 660618 322066 660854
rect 322302 660618 349746 660854
rect 349982 660618 350066 660854
rect 350302 660618 377746 660854
rect 377982 660618 378066 660854
rect 378302 660618 405746 660854
rect 405982 660618 406066 660854
rect 406302 660618 433746 660854
rect 433982 660618 434066 660854
rect 434302 660618 461746 660854
rect 461982 660618 462066 660854
rect 462302 660618 489746 660854
rect 489982 660618 490066 660854
rect 490302 660618 517746 660854
rect 517982 660618 518066 660854
rect 518302 660618 545746 660854
rect 545982 660618 546066 660854
rect 546302 660618 573746 660854
rect 573982 660618 574066 660854
rect 574302 660618 585342 660854
rect 585578 660618 585662 660854
rect 585898 660618 592650 660854
rect -8726 660586 592650 660618
rect -8726 657454 592650 657486
rect -8726 657218 -2934 657454
rect -2698 657218 -2614 657454
rect -2378 657218 38026 657454
rect 38262 657218 38346 657454
rect 38582 657218 66026 657454
rect 66262 657218 66346 657454
rect 66582 657218 94026 657454
rect 94262 657218 94346 657454
rect 94582 657218 122026 657454
rect 122262 657218 122346 657454
rect 122582 657218 150026 657454
rect 150262 657218 150346 657454
rect 150582 657218 178026 657454
rect 178262 657218 178346 657454
rect 178582 657218 206026 657454
rect 206262 657218 206346 657454
rect 206582 657218 234026 657454
rect 234262 657218 234346 657454
rect 234582 657218 262026 657454
rect 262262 657218 262346 657454
rect 262582 657218 290026 657454
rect 290262 657218 290346 657454
rect 290582 657218 318026 657454
rect 318262 657218 318346 657454
rect 318582 657218 346026 657454
rect 346262 657218 346346 657454
rect 346582 657218 374026 657454
rect 374262 657218 374346 657454
rect 374582 657218 402026 657454
rect 402262 657218 402346 657454
rect 402582 657218 430026 657454
rect 430262 657218 430346 657454
rect 430582 657218 458026 657454
rect 458262 657218 458346 657454
rect 458582 657218 486026 657454
rect 486262 657218 486346 657454
rect 486582 657218 514026 657454
rect 514262 657218 514346 657454
rect 514582 657218 542026 657454
rect 542262 657218 542346 657454
rect 542582 657218 570026 657454
rect 570262 657218 570346 657454
rect 570582 657218 586302 657454
rect 586538 657218 586622 657454
rect 586858 657218 592650 657454
rect -8726 657134 592650 657218
rect -8726 656898 -2934 657134
rect -2698 656898 -2614 657134
rect -2378 656898 38026 657134
rect 38262 656898 38346 657134
rect 38582 656898 66026 657134
rect 66262 656898 66346 657134
rect 66582 656898 94026 657134
rect 94262 656898 94346 657134
rect 94582 656898 122026 657134
rect 122262 656898 122346 657134
rect 122582 656898 150026 657134
rect 150262 656898 150346 657134
rect 150582 656898 178026 657134
rect 178262 656898 178346 657134
rect 178582 656898 206026 657134
rect 206262 656898 206346 657134
rect 206582 656898 234026 657134
rect 234262 656898 234346 657134
rect 234582 656898 262026 657134
rect 262262 656898 262346 657134
rect 262582 656898 290026 657134
rect 290262 656898 290346 657134
rect 290582 656898 318026 657134
rect 318262 656898 318346 657134
rect 318582 656898 346026 657134
rect 346262 656898 346346 657134
rect 346582 656898 374026 657134
rect 374262 656898 374346 657134
rect 374582 656898 402026 657134
rect 402262 656898 402346 657134
rect 402582 656898 430026 657134
rect 430262 656898 430346 657134
rect 430582 656898 458026 657134
rect 458262 656898 458346 657134
rect 458582 656898 486026 657134
rect 486262 656898 486346 657134
rect 486582 656898 514026 657134
rect 514262 656898 514346 657134
rect 514582 656898 542026 657134
rect 542262 656898 542346 657134
rect 542582 656898 570026 657134
rect 570262 656898 570346 657134
rect 570582 656898 586302 657134
rect 586538 656898 586622 657134
rect 586858 656898 592650 657134
rect -8726 656866 592650 656898
rect -8726 624174 592650 624206
rect -8726 623938 -1974 624174
rect -1738 623938 -1654 624174
rect -1418 623938 41746 624174
rect 41982 623938 42066 624174
rect 42302 623938 69746 624174
rect 69982 623938 70066 624174
rect 70302 623938 97746 624174
rect 97982 623938 98066 624174
rect 98302 623938 125746 624174
rect 125982 623938 126066 624174
rect 126302 623938 153746 624174
rect 153982 623938 154066 624174
rect 154302 623938 181746 624174
rect 181982 623938 182066 624174
rect 182302 623938 209746 624174
rect 209982 623938 210066 624174
rect 210302 623938 237746 624174
rect 237982 623938 238066 624174
rect 238302 623938 265746 624174
rect 265982 623938 266066 624174
rect 266302 623938 293746 624174
rect 293982 623938 294066 624174
rect 294302 623938 321746 624174
rect 321982 623938 322066 624174
rect 322302 623938 349746 624174
rect 349982 623938 350066 624174
rect 350302 623938 377746 624174
rect 377982 623938 378066 624174
rect 378302 623938 405746 624174
rect 405982 623938 406066 624174
rect 406302 623938 433746 624174
rect 433982 623938 434066 624174
rect 434302 623938 461746 624174
rect 461982 623938 462066 624174
rect 462302 623938 489746 624174
rect 489982 623938 490066 624174
rect 490302 623938 517746 624174
rect 517982 623938 518066 624174
rect 518302 623938 545746 624174
rect 545982 623938 546066 624174
rect 546302 623938 573746 624174
rect 573982 623938 574066 624174
rect 574302 623938 585342 624174
rect 585578 623938 585662 624174
rect 585898 623938 592650 624174
rect -8726 623854 592650 623938
rect -8726 623618 -1974 623854
rect -1738 623618 -1654 623854
rect -1418 623618 41746 623854
rect 41982 623618 42066 623854
rect 42302 623618 69746 623854
rect 69982 623618 70066 623854
rect 70302 623618 97746 623854
rect 97982 623618 98066 623854
rect 98302 623618 125746 623854
rect 125982 623618 126066 623854
rect 126302 623618 153746 623854
rect 153982 623618 154066 623854
rect 154302 623618 181746 623854
rect 181982 623618 182066 623854
rect 182302 623618 209746 623854
rect 209982 623618 210066 623854
rect 210302 623618 237746 623854
rect 237982 623618 238066 623854
rect 238302 623618 265746 623854
rect 265982 623618 266066 623854
rect 266302 623618 293746 623854
rect 293982 623618 294066 623854
rect 294302 623618 321746 623854
rect 321982 623618 322066 623854
rect 322302 623618 349746 623854
rect 349982 623618 350066 623854
rect 350302 623618 377746 623854
rect 377982 623618 378066 623854
rect 378302 623618 405746 623854
rect 405982 623618 406066 623854
rect 406302 623618 433746 623854
rect 433982 623618 434066 623854
rect 434302 623618 461746 623854
rect 461982 623618 462066 623854
rect 462302 623618 489746 623854
rect 489982 623618 490066 623854
rect 490302 623618 517746 623854
rect 517982 623618 518066 623854
rect 518302 623618 545746 623854
rect 545982 623618 546066 623854
rect 546302 623618 573746 623854
rect 573982 623618 574066 623854
rect 574302 623618 585342 623854
rect 585578 623618 585662 623854
rect 585898 623618 592650 623854
rect -8726 623586 592650 623618
rect -8726 620454 592650 620486
rect -8726 620218 -2934 620454
rect -2698 620218 -2614 620454
rect -2378 620218 38026 620454
rect 38262 620218 38346 620454
rect 38582 620218 66026 620454
rect 66262 620218 66346 620454
rect 66582 620218 94026 620454
rect 94262 620218 94346 620454
rect 94582 620218 122026 620454
rect 122262 620218 122346 620454
rect 122582 620218 150026 620454
rect 150262 620218 150346 620454
rect 150582 620218 178026 620454
rect 178262 620218 178346 620454
rect 178582 620218 206026 620454
rect 206262 620218 206346 620454
rect 206582 620218 234026 620454
rect 234262 620218 234346 620454
rect 234582 620218 262026 620454
rect 262262 620218 262346 620454
rect 262582 620218 290026 620454
rect 290262 620218 290346 620454
rect 290582 620218 318026 620454
rect 318262 620218 318346 620454
rect 318582 620218 346026 620454
rect 346262 620218 346346 620454
rect 346582 620218 374026 620454
rect 374262 620218 374346 620454
rect 374582 620218 402026 620454
rect 402262 620218 402346 620454
rect 402582 620218 430026 620454
rect 430262 620218 430346 620454
rect 430582 620218 458026 620454
rect 458262 620218 458346 620454
rect 458582 620218 486026 620454
rect 486262 620218 486346 620454
rect 486582 620218 514026 620454
rect 514262 620218 514346 620454
rect 514582 620218 542026 620454
rect 542262 620218 542346 620454
rect 542582 620218 570026 620454
rect 570262 620218 570346 620454
rect 570582 620218 586302 620454
rect 586538 620218 586622 620454
rect 586858 620218 592650 620454
rect -8726 620134 592650 620218
rect -8726 619898 -2934 620134
rect -2698 619898 -2614 620134
rect -2378 619898 38026 620134
rect 38262 619898 38346 620134
rect 38582 619898 66026 620134
rect 66262 619898 66346 620134
rect 66582 619898 94026 620134
rect 94262 619898 94346 620134
rect 94582 619898 122026 620134
rect 122262 619898 122346 620134
rect 122582 619898 150026 620134
rect 150262 619898 150346 620134
rect 150582 619898 178026 620134
rect 178262 619898 178346 620134
rect 178582 619898 206026 620134
rect 206262 619898 206346 620134
rect 206582 619898 234026 620134
rect 234262 619898 234346 620134
rect 234582 619898 262026 620134
rect 262262 619898 262346 620134
rect 262582 619898 290026 620134
rect 290262 619898 290346 620134
rect 290582 619898 318026 620134
rect 318262 619898 318346 620134
rect 318582 619898 346026 620134
rect 346262 619898 346346 620134
rect 346582 619898 374026 620134
rect 374262 619898 374346 620134
rect 374582 619898 402026 620134
rect 402262 619898 402346 620134
rect 402582 619898 430026 620134
rect 430262 619898 430346 620134
rect 430582 619898 458026 620134
rect 458262 619898 458346 620134
rect 458582 619898 486026 620134
rect 486262 619898 486346 620134
rect 486582 619898 514026 620134
rect 514262 619898 514346 620134
rect 514582 619898 542026 620134
rect 542262 619898 542346 620134
rect 542582 619898 570026 620134
rect 570262 619898 570346 620134
rect 570582 619898 586302 620134
rect 586538 619898 586622 620134
rect 586858 619898 592650 620134
rect -8726 619866 592650 619898
rect -8726 587174 592650 587206
rect -8726 586938 -1974 587174
rect -1738 586938 -1654 587174
rect -1418 586938 41746 587174
rect 41982 586938 42066 587174
rect 42302 586938 69746 587174
rect 69982 586938 70066 587174
rect 70302 586938 97746 587174
rect 97982 586938 98066 587174
rect 98302 586938 125746 587174
rect 125982 586938 126066 587174
rect 126302 586938 153746 587174
rect 153982 586938 154066 587174
rect 154302 586938 181746 587174
rect 181982 586938 182066 587174
rect 182302 586938 209746 587174
rect 209982 586938 210066 587174
rect 210302 586938 237746 587174
rect 237982 586938 238066 587174
rect 238302 586938 265746 587174
rect 265982 586938 266066 587174
rect 266302 586938 293746 587174
rect 293982 586938 294066 587174
rect 294302 586938 321746 587174
rect 321982 586938 322066 587174
rect 322302 586938 349746 587174
rect 349982 586938 350066 587174
rect 350302 586938 377746 587174
rect 377982 586938 378066 587174
rect 378302 586938 405746 587174
rect 405982 586938 406066 587174
rect 406302 586938 433746 587174
rect 433982 586938 434066 587174
rect 434302 586938 461746 587174
rect 461982 586938 462066 587174
rect 462302 586938 489746 587174
rect 489982 586938 490066 587174
rect 490302 586938 517746 587174
rect 517982 586938 518066 587174
rect 518302 586938 545746 587174
rect 545982 586938 546066 587174
rect 546302 586938 573746 587174
rect 573982 586938 574066 587174
rect 574302 586938 585342 587174
rect 585578 586938 585662 587174
rect 585898 586938 592650 587174
rect -8726 586854 592650 586938
rect -8726 586618 -1974 586854
rect -1738 586618 -1654 586854
rect -1418 586618 41746 586854
rect 41982 586618 42066 586854
rect 42302 586618 69746 586854
rect 69982 586618 70066 586854
rect 70302 586618 97746 586854
rect 97982 586618 98066 586854
rect 98302 586618 125746 586854
rect 125982 586618 126066 586854
rect 126302 586618 153746 586854
rect 153982 586618 154066 586854
rect 154302 586618 181746 586854
rect 181982 586618 182066 586854
rect 182302 586618 209746 586854
rect 209982 586618 210066 586854
rect 210302 586618 237746 586854
rect 237982 586618 238066 586854
rect 238302 586618 265746 586854
rect 265982 586618 266066 586854
rect 266302 586618 293746 586854
rect 293982 586618 294066 586854
rect 294302 586618 321746 586854
rect 321982 586618 322066 586854
rect 322302 586618 349746 586854
rect 349982 586618 350066 586854
rect 350302 586618 377746 586854
rect 377982 586618 378066 586854
rect 378302 586618 405746 586854
rect 405982 586618 406066 586854
rect 406302 586618 433746 586854
rect 433982 586618 434066 586854
rect 434302 586618 461746 586854
rect 461982 586618 462066 586854
rect 462302 586618 489746 586854
rect 489982 586618 490066 586854
rect 490302 586618 517746 586854
rect 517982 586618 518066 586854
rect 518302 586618 545746 586854
rect 545982 586618 546066 586854
rect 546302 586618 573746 586854
rect 573982 586618 574066 586854
rect 574302 586618 585342 586854
rect 585578 586618 585662 586854
rect 585898 586618 592650 586854
rect -8726 586586 592650 586618
rect -8726 583454 592650 583486
rect -8726 583218 -2934 583454
rect -2698 583218 -2614 583454
rect -2378 583218 38026 583454
rect 38262 583218 38346 583454
rect 38582 583218 66026 583454
rect 66262 583218 66346 583454
rect 66582 583218 94026 583454
rect 94262 583218 94346 583454
rect 94582 583218 122026 583454
rect 122262 583218 122346 583454
rect 122582 583218 150026 583454
rect 150262 583218 150346 583454
rect 150582 583218 178026 583454
rect 178262 583218 178346 583454
rect 178582 583218 206026 583454
rect 206262 583218 206346 583454
rect 206582 583218 234026 583454
rect 234262 583218 234346 583454
rect 234582 583218 262026 583454
rect 262262 583218 262346 583454
rect 262582 583218 290026 583454
rect 290262 583218 290346 583454
rect 290582 583218 318026 583454
rect 318262 583218 318346 583454
rect 318582 583218 346026 583454
rect 346262 583218 346346 583454
rect 346582 583218 374026 583454
rect 374262 583218 374346 583454
rect 374582 583218 402026 583454
rect 402262 583218 402346 583454
rect 402582 583218 430026 583454
rect 430262 583218 430346 583454
rect 430582 583218 458026 583454
rect 458262 583218 458346 583454
rect 458582 583218 486026 583454
rect 486262 583218 486346 583454
rect 486582 583218 514026 583454
rect 514262 583218 514346 583454
rect 514582 583218 542026 583454
rect 542262 583218 542346 583454
rect 542582 583218 570026 583454
rect 570262 583218 570346 583454
rect 570582 583218 586302 583454
rect 586538 583218 586622 583454
rect 586858 583218 592650 583454
rect -8726 583134 592650 583218
rect -8726 582898 -2934 583134
rect -2698 582898 -2614 583134
rect -2378 582898 38026 583134
rect 38262 582898 38346 583134
rect 38582 582898 66026 583134
rect 66262 582898 66346 583134
rect 66582 582898 94026 583134
rect 94262 582898 94346 583134
rect 94582 582898 122026 583134
rect 122262 582898 122346 583134
rect 122582 582898 150026 583134
rect 150262 582898 150346 583134
rect 150582 582898 178026 583134
rect 178262 582898 178346 583134
rect 178582 582898 206026 583134
rect 206262 582898 206346 583134
rect 206582 582898 234026 583134
rect 234262 582898 234346 583134
rect 234582 582898 262026 583134
rect 262262 582898 262346 583134
rect 262582 582898 290026 583134
rect 290262 582898 290346 583134
rect 290582 582898 318026 583134
rect 318262 582898 318346 583134
rect 318582 582898 346026 583134
rect 346262 582898 346346 583134
rect 346582 582898 374026 583134
rect 374262 582898 374346 583134
rect 374582 582898 402026 583134
rect 402262 582898 402346 583134
rect 402582 582898 430026 583134
rect 430262 582898 430346 583134
rect 430582 582898 458026 583134
rect 458262 582898 458346 583134
rect 458582 582898 486026 583134
rect 486262 582898 486346 583134
rect 486582 582898 514026 583134
rect 514262 582898 514346 583134
rect 514582 582898 542026 583134
rect 542262 582898 542346 583134
rect 542582 582898 570026 583134
rect 570262 582898 570346 583134
rect 570582 582898 586302 583134
rect 586538 582898 586622 583134
rect 586858 582898 592650 583134
rect -8726 582866 592650 582898
rect -8726 550174 592650 550206
rect -8726 549938 -1974 550174
rect -1738 549938 -1654 550174
rect -1418 549938 41746 550174
rect 41982 549938 42066 550174
rect 42302 549938 69746 550174
rect 69982 549938 70066 550174
rect 70302 549938 97746 550174
rect 97982 549938 98066 550174
rect 98302 549938 125746 550174
rect 125982 549938 126066 550174
rect 126302 549938 153746 550174
rect 153982 549938 154066 550174
rect 154302 549938 181746 550174
rect 181982 549938 182066 550174
rect 182302 549938 209746 550174
rect 209982 549938 210066 550174
rect 210302 549938 237746 550174
rect 237982 549938 238066 550174
rect 238302 549938 265746 550174
rect 265982 549938 266066 550174
rect 266302 549938 293746 550174
rect 293982 549938 294066 550174
rect 294302 549938 321746 550174
rect 321982 549938 322066 550174
rect 322302 549938 349746 550174
rect 349982 549938 350066 550174
rect 350302 549938 377746 550174
rect 377982 549938 378066 550174
rect 378302 549938 405746 550174
rect 405982 549938 406066 550174
rect 406302 549938 433746 550174
rect 433982 549938 434066 550174
rect 434302 549938 461746 550174
rect 461982 549938 462066 550174
rect 462302 549938 489746 550174
rect 489982 549938 490066 550174
rect 490302 549938 517746 550174
rect 517982 549938 518066 550174
rect 518302 549938 545746 550174
rect 545982 549938 546066 550174
rect 546302 549938 573746 550174
rect 573982 549938 574066 550174
rect 574302 549938 585342 550174
rect 585578 549938 585662 550174
rect 585898 549938 592650 550174
rect -8726 549854 592650 549938
rect -8726 549618 -1974 549854
rect -1738 549618 -1654 549854
rect -1418 549618 41746 549854
rect 41982 549618 42066 549854
rect 42302 549618 69746 549854
rect 69982 549618 70066 549854
rect 70302 549618 97746 549854
rect 97982 549618 98066 549854
rect 98302 549618 125746 549854
rect 125982 549618 126066 549854
rect 126302 549618 153746 549854
rect 153982 549618 154066 549854
rect 154302 549618 181746 549854
rect 181982 549618 182066 549854
rect 182302 549618 209746 549854
rect 209982 549618 210066 549854
rect 210302 549618 237746 549854
rect 237982 549618 238066 549854
rect 238302 549618 265746 549854
rect 265982 549618 266066 549854
rect 266302 549618 293746 549854
rect 293982 549618 294066 549854
rect 294302 549618 321746 549854
rect 321982 549618 322066 549854
rect 322302 549618 349746 549854
rect 349982 549618 350066 549854
rect 350302 549618 377746 549854
rect 377982 549618 378066 549854
rect 378302 549618 405746 549854
rect 405982 549618 406066 549854
rect 406302 549618 433746 549854
rect 433982 549618 434066 549854
rect 434302 549618 461746 549854
rect 461982 549618 462066 549854
rect 462302 549618 489746 549854
rect 489982 549618 490066 549854
rect 490302 549618 517746 549854
rect 517982 549618 518066 549854
rect 518302 549618 545746 549854
rect 545982 549618 546066 549854
rect 546302 549618 573746 549854
rect 573982 549618 574066 549854
rect 574302 549618 585342 549854
rect 585578 549618 585662 549854
rect 585898 549618 592650 549854
rect -8726 549586 592650 549618
rect -8726 546454 592650 546486
rect -8726 546218 -2934 546454
rect -2698 546218 -2614 546454
rect -2378 546218 38026 546454
rect 38262 546218 38346 546454
rect 38582 546218 66026 546454
rect 66262 546218 66346 546454
rect 66582 546218 94026 546454
rect 94262 546218 94346 546454
rect 94582 546218 122026 546454
rect 122262 546218 122346 546454
rect 122582 546218 150026 546454
rect 150262 546218 150346 546454
rect 150582 546218 178026 546454
rect 178262 546218 178346 546454
rect 178582 546218 206026 546454
rect 206262 546218 206346 546454
rect 206582 546218 234026 546454
rect 234262 546218 234346 546454
rect 234582 546218 262026 546454
rect 262262 546218 262346 546454
rect 262582 546218 290026 546454
rect 290262 546218 290346 546454
rect 290582 546218 318026 546454
rect 318262 546218 318346 546454
rect 318582 546218 346026 546454
rect 346262 546218 346346 546454
rect 346582 546218 374026 546454
rect 374262 546218 374346 546454
rect 374582 546218 402026 546454
rect 402262 546218 402346 546454
rect 402582 546218 430026 546454
rect 430262 546218 430346 546454
rect 430582 546218 458026 546454
rect 458262 546218 458346 546454
rect 458582 546218 486026 546454
rect 486262 546218 486346 546454
rect 486582 546218 514026 546454
rect 514262 546218 514346 546454
rect 514582 546218 542026 546454
rect 542262 546218 542346 546454
rect 542582 546218 570026 546454
rect 570262 546218 570346 546454
rect 570582 546218 586302 546454
rect 586538 546218 586622 546454
rect 586858 546218 592650 546454
rect -8726 546134 592650 546218
rect -8726 545898 -2934 546134
rect -2698 545898 -2614 546134
rect -2378 545898 38026 546134
rect 38262 545898 38346 546134
rect 38582 545898 66026 546134
rect 66262 545898 66346 546134
rect 66582 545898 94026 546134
rect 94262 545898 94346 546134
rect 94582 545898 122026 546134
rect 122262 545898 122346 546134
rect 122582 545898 150026 546134
rect 150262 545898 150346 546134
rect 150582 545898 178026 546134
rect 178262 545898 178346 546134
rect 178582 545898 206026 546134
rect 206262 545898 206346 546134
rect 206582 545898 234026 546134
rect 234262 545898 234346 546134
rect 234582 545898 262026 546134
rect 262262 545898 262346 546134
rect 262582 545898 290026 546134
rect 290262 545898 290346 546134
rect 290582 545898 318026 546134
rect 318262 545898 318346 546134
rect 318582 545898 346026 546134
rect 346262 545898 346346 546134
rect 346582 545898 374026 546134
rect 374262 545898 374346 546134
rect 374582 545898 402026 546134
rect 402262 545898 402346 546134
rect 402582 545898 430026 546134
rect 430262 545898 430346 546134
rect 430582 545898 458026 546134
rect 458262 545898 458346 546134
rect 458582 545898 486026 546134
rect 486262 545898 486346 546134
rect 486582 545898 514026 546134
rect 514262 545898 514346 546134
rect 514582 545898 542026 546134
rect 542262 545898 542346 546134
rect 542582 545898 570026 546134
rect 570262 545898 570346 546134
rect 570582 545898 586302 546134
rect 586538 545898 586622 546134
rect 586858 545898 592650 546134
rect -8726 545866 592650 545898
rect -8726 513174 592650 513206
rect -8726 512938 -1974 513174
rect -1738 512938 -1654 513174
rect -1418 512938 41746 513174
rect 41982 512938 42066 513174
rect 42302 512938 69746 513174
rect 69982 512938 70066 513174
rect 70302 512938 97746 513174
rect 97982 512938 98066 513174
rect 98302 512938 125746 513174
rect 125982 512938 126066 513174
rect 126302 512938 153746 513174
rect 153982 512938 154066 513174
rect 154302 512938 181746 513174
rect 181982 512938 182066 513174
rect 182302 512938 209746 513174
rect 209982 512938 210066 513174
rect 210302 512938 237746 513174
rect 237982 512938 238066 513174
rect 238302 512938 265746 513174
rect 265982 512938 266066 513174
rect 266302 512938 293746 513174
rect 293982 512938 294066 513174
rect 294302 512938 321746 513174
rect 321982 512938 322066 513174
rect 322302 512938 349746 513174
rect 349982 512938 350066 513174
rect 350302 512938 377746 513174
rect 377982 512938 378066 513174
rect 378302 512938 405746 513174
rect 405982 512938 406066 513174
rect 406302 512938 433746 513174
rect 433982 512938 434066 513174
rect 434302 512938 461746 513174
rect 461982 512938 462066 513174
rect 462302 512938 489746 513174
rect 489982 512938 490066 513174
rect 490302 512938 517746 513174
rect 517982 512938 518066 513174
rect 518302 512938 545746 513174
rect 545982 512938 546066 513174
rect 546302 512938 573746 513174
rect 573982 512938 574066 513174
rect 574302 512938 585342 513174
rect 585578 512938 585662 513174
rect 585898 512938 592650 513174
rect -8726 512854 592650 512938
rect -8726 512618 -1974 512854
rect -1738 512618 -1654 512854
rect -1418 512618 41746 512854
rect 41982 512618 42066 512854
rect 42302 512618 69746 512854
rect 69982 512618 70066 512854
rect 70302 512618 97746 512854
rect 97982 512618 98066 512854
rect 98302 512618 125746 512854
rect 125982 512618 126066 512854
rect 126302 512618 153746 512854
rect 153982 512618 154066 512854
rect 154302 512618 181746 512854
rect 181982 512618 182066 512854
rect 182302 512618 209746 512854
rect 209982 512618 210066 512854
rect 210302 512618 237746 512854
rect 237982 512618 238066 512854
rect 238302 512618 265746 512854
rect 265982 512618 266066 512854
rect 266302 512618 293746 512854
rect 293982 512618 294066 512854
rect 294302 512618 321746 512854
rect 321982 512618 322066 512854
rect 322302 512618 349746 512854
rect 349982 512618 350066 512854
rect 350302 512618 377746 512854
rect 377982 512618 378066 512854
rect 378302 512618 405746 512854
rect 405982 512618 406066 512854
rect 406302 512618 433746 512854
rect 433982 512618 434066 512854
rect 434302 512618 461746 512854
rect 461982 512618 462066 512854
rect 462302 512618 489746 512854
rect 489982 512618 490066 512854
rect 490302 512618 517746 512854
rect 517982 512618 518066 512854
rect 518302 512618 545746 512854
rect 545982 512618 546066 512854
rect 546302 512618 573746 512854
rect 573982 512618 574066 512854
rect 574302 512618 585342 512854
rect 585578 512618 585662 512854
rect 585898 512618 592650 512854
rect -8726 512586 592650 512618
rect -8726 509454 592650 509486
rect -8726 509218 -2934 509454
rect -2698 509218 -2614 509454
rect -2378 509218 38026 509454
rect 38262 509218 38346 509454
rect 38582 509218 66026 509454
rect 66262 509218 66346 509454
rect 66582 509218 94026 509454
rect 94262 509218 94346 509454
rect 94582 509218 122026 509454
rect 122262 509218 122346 509454
rect 122582 509218 150026 509454
rect 150262 509218 150346 509454
rect 150582 509218 178026 509454
rect 178262 509218 178346 509454
rect 178582 509218 206026 509454
rect 206262 509218 206346 509454
rect 206582 509218 234026 509454
rect 234262 509218 234346 509454
rect 234582 509218 262026 509454
rect 262262 509218 262346 509454
rect 262582 509218 290026 509454
rect 290262 509218 290346 509454
rect 290582 509218 318026 509454
rect 318262 509218 318346 509454
rect 318582 509218 346026 509454
rect 346262 509218 346346 509454
rect 346582 509218 374026 509454
rect 374262 509218 374346 509454
rect 374582 509218 402026 509454
rect 402262 509218 402346 509454
rect 402582 509218 430026 509454
rect 430262 509218 430346 509454
rect 430582 509218 458026 509454
rect 458262 509218 458346 509454
rect 458582 509218 486026 509454
rect 486262 509218 486346 509454
rect 486582 509218 514026 509454
rect 514262 509218 514346 509454
rect 514582 509218 542026 509454
rect 542262 509218 542346 509454
rect 542582 509218 570026 509454
rect 570262 509218 570346 509454
rect 570582 509218 586302 509454
rect 586538 509218 586622 509454
rect 586858 509218 592650 509454
rect -8726 509134 592650 509218
rect -8726 508898 -2934 509134
rect -2698 508898 -2614 509134
rect -2378 508898 38026 509134
rect 38262 508898 38346 509134
rect 38582 508898 66026 509134
rect 66262 508898 66346 509134
rect 66582 508898 94026 509134
rect 94262 508898 94346 509134
rect 94582 508898 122026 509134
rect 122262 508898 122346 509134
rect 122582 508898 150026 509134
rect 150262 508898 150346 509134
rect 150582 508898 178026 509134
rect 178262 508898 178346 509134
rect 178582 508898 206026 509134
rect 206262 508898 206346 509134
rect 206582 508898 234026 509134
rect 234262 508898 234346 509134
rect 234582 508898 262026 509134
rect 262262 508898 262346 509134
rect 262582 508898 290026 509134
rect 290262 508898 290346 509134
rect 290582 508898 318026 509134
rect 318262 508898 318346 509134
rect 318582 508898 346026 509134
rect 346262 508898 346346 509134
rect 346582 508898 374026 509134
rect 374262 508898 374346 509134
rect 374582 508898 402026 509134
rect 402262 508898 402346 509134
rect 402582 508898 430026 509134
rect 430262 508898 430346 509134
rect 430582 508898 458026 509134
rect 458262 508898 458346 509134
rect 458582 508898 486026 509134
rect 486262 508898 486346 509134
rect 486582 508898 514026 509134
rect 514262 508898 514346 509134
rect 514582 508898 542026 509134
rect 542262 508898 542346 509134
rect 542582 508898 570026 509134
rect 570262 508898 570346 509134
rect 570582 508898 586302 509134
rect 586538 508898 586622 509134
rect 586858 508898 592650 509134
rect -8726 508866 592650 508898
rect -8726 476174 592650 476206
rect -8726 475938 -1974 476174
rect -1738 475938 -1654 476174
rect -1418 475938 41746 476174
rect 41982 475938 42066 476174
rect 42302 475938 69746 476174
rect 69982 475938 70066 476174
rect 70302 475938 97746 476174
rect 97982 475938 98066 476174
rect 98302 475938 125746 476174
rect 125982 475938 126066 476174
rect 126302 475938 153746 476174
rect 153982 475938 154066 476174
rect 154302 475938 181746 476174
rect 181982 475938 182066 476174
rect 182302 475938 209746 476174
rect 209982 475938 210066 476174
rect 210302 475938 237746 476174
rect 237982 475938 238066 476174
rect 238302 475938 265746 476174
rect 265982 475938 266066 476174
rect 266302 475938 293746 476174
rect 293982 475938 294066 476174
rect 294302 475938 321746 476174
rect 321982 475938 322066 476174
rect 322302 475938 349746 476174
rect 349982 475938 350066 476174
rect 350302 475938 377746 476174
rect 377982 475938 378066 476174
rect 378302 475938 405746 476174
rect 405982 475938 406066 476174
rect 406302 475938 433746 476174
rect 433982 475938 434066 476174
rect 434302 475938 461746 476174
rect 461982 475938 462066 476174
rect 462302 475938 489746 476174
rect 489982 475938 490066 476174
rect 490302 475938 517746 476174
rect 517982 475938 518066 476174
rect 518302 475938 545746 476174
rect 545982 475938 546066 476174
rect 546302 475938 573746 476174
rect 573982 475938 574066 476174
rect 574302 475938 585342 476174
rect 585578 475938 585662 476174
rect 585898 475938 592650 476174
rect -8726 475854 592650 475938
rect -8726 475618 -1974 475854
rect -1738 475618 -1654 475854
rect -1418 475618 41746 475854
rect 41982 475618 42066 475854
rect 42302 475618 69746 475854
rect 69982 475618 70066 475854
rect 70302 475618 97746 475854
rect 97982 475618 98066 475854
rect 98302 475618 125746 475854
rect 125982 475618 126066 475854
rect 126302 475618 153746 475854
rect 153982 475618 154066 475854
rect 154302 475618 181746 475854
rect 181982 475618 182066 475854
rect 182302 475618 209746 475854
rect 209982 475618 210066 475854
rect 210302 475618 237746 475854
rect 237982 475618 238066 475854
rect 238302 475618 265746 475854
rect 265982 475618 266066 475854
rect 266302 475618 293746 475854
rect 293982 475618 294066 475854
rect 294302 475618 321746 475854
rect 321982 475618 322066 475854
rect 322302 475618 349746 475854
rect 349982 475618 350066 475854
rect 350302 475618 377746 475854
rect 377982 475618 378066 475854
rect 378302 475618 405746 475854
rect 405982 475618 406066 475854
rect 406302 475618 433746 475854
rect 433982 475618 434066 475854
rect 434302 475618 461746 475854
rect 461982 475618 462066 475854
rect 462302 475618 489746 475854
rect 489982 475618 490066 475854
rect 490302 475618 517746 475854
rect 517982 475618 518066 475854
rect 518302 475618 545746 475854
rect 545982 475618 546066 475854
rect 546302 475618 573746 475854
rect 573982 475618 574066 475854
rect 574302 475618 585342 475854
rect 585578 475618 585662 475854
rect 585898 475618 592650 475854
rect -8726 475586 592650 475618
rect -8726 472454 592650 472486
rect -8726 472218 -2934 472454
rect -2698 472218 -2614 472454
rect -2378 472218 38026 472454
rect 38262 472218 38346 472454
rect 38582 472218 66026 472454
rect 66262 472218 66346 472454
rect 66582 472218 94026 472454
rect 94262 472218 94346 472454
rect 94582 472218 122026 472454
rect 122262 472218 122346 472454
rect 122582 472218 150026 472454
rect 150262 472218 150346 472454
rect 150582 472218 178026 472454
rect 178262 472218 178346 472454
rect 178582 472218 206026 472454
rect 206262 472218 206346 472454
rect 206582 472218 234026 472454
rect 234262 472218 234346 472454
rect 234582 472218 262026 472454
rect 262262 472218 262346 472454
rect 262582 472218 290026 472454
rect 290262 472218 290346 472454
rect 290582 472218 318026 472454
rect 318262 472218 318346 472454
rect 318582 472218 346026 472454
rect 346262 472218 346346 472454
rect 346582 472218 374026 472454
rect 374262 472218 374346 472454
rect 374582 472218 402026 472454
rect 402262 472218 402346 472454
rect 402582 472218 430026 472454
rect 430262 472218 430346 472454
rect 430582 472218 458026 472454
rect 458262 472218 458346 472454
rect 458582 472218 486026 472454
rect 486262 472218 486346 472454
rect 486582 472218 514026 472454
rect 514262 472218 514346 472454
rect 514582 472218 542026 472454
rect 542262 472218 542346 472454
rect 542582 472218 570026 472454
rect 570262 472218 570346 472454
rect 570582 472218 586302 472454
rect 586538 472218 586622 472454
rect 586858 472218 592650 472454
rect -8726 472134 592650 472218
rect -8726 471898 -2934 472134
rect -2698 471898 -2614 472134
rect -2378 471898 38026 472134
rect 38262 471898 38346 472134
rect 38582 471898 66026 472134
rect 66262 471898 66346 472134
rect 66582 471898 94026 472134
rect 94262 471898 94346 472134
rect 94582 471898 122026 472134
rect 122262 471898 122346 472134
rect 122582 471898 150026 472134
rect 150262 471898 150346 472134
rect 150582 471898 178026 472134
rect 178262 471898 178346 472134
rect 178582 471898 206026 472134
rect 206262 471898 206346 472134
rect 206582 471898 234026 472134
rect 234262 471898 234346 472134
rect 234582 471898 262026 472134
rect 262262 471898 262346 472134
rect 262582 471898 290026 472134
rect 290262 471898 290346 472134
rect 290582 471898 318026 472134
rect 318262 471898 318346 472134
rect 318582 471898 346026 472134
rect 346262 471898 346346 472134
rect 346582 471898 374026 472134
rect 374262 471898 374346 472134
rect 374582 471898 402026 472134
rect 402262 471898 402346 472134
rect 402582 471898 430026 472134
rect 430262 471898 430346 472134
rect 430582 471898 458026 472134
rect 458262 471898 458346 472134
rect 458582 471898 486026 472134
rect 486262 471898 486346 472134
rect 486582 471898 514026 472134
rect 514262 471898 514346 472134
rect 514582 471898 542026 472134
rect 542262 471898 542346 472134
rect 542582 471898 570026 472134
rect 570262 471898 570346 472134
rect 570582 471898 586302 472134
rect 586538 471898 586622 472134
rect 586858 471898 592650 472134
rect -8726 471866 592650 471898
rect -8726 439174 592650 439206
rect -8726 438938 -1974 439174
rect -1738 438938 -1654 439174
rect -1418 438938 41746 439174
rect 41982 438938 42066 439174
rect 42302 438938 69746 439174
rect 69982 438938 70066 439174
rect 70302 438938 97746 439174
rect 97982 438938 98066 439174
rect 98302 438938 125746 439174
rect 125982 438938 126066 439174
rect 126302 438938 153746 439174
rect 153982 438938 154066 439174
rect 154302 438938 181746 439174
rect 181982 438938 182066 439174
rect 182302 438938 209746 439174
rect 209982 438938 210066 439174
rect 210302 438938 237746 439174
rect 237982 438938 238066 439174
rect 238302 438938 265746 439174
rect 265982 438938 266066 439174
rect 266302 438938 293746 439174
rect 293982 438938 294066 439174
rect 294302 438938 321746 439174
rect 321982 438938 322066 439174
rect 322302 438938 349746 439174
rect 349982 438938 350066 439174
rect 350302 438938 377746 439174
rect 377982 438938 378066 439174
rect 378302 438938 405746 439174
rect 405982 438938 406066 439174
rect 406302 438938 433746 439174
rect 433982 438938 434066 439174
rect 434302 438938 461746 439174
rect 461982 438938 462066 439174
rect 462302 438938 489746 439174
rect 489982 438938 490066 439174
rect 490302 438938 517746 439174
rect 517982 438938 518066 439174
rect 518302 438938 545746 439174
rect 545982 438938 546066 439174
rect 546302 438938 573746 439174
rect 573982 438938 574066 439174
rect 574302 438938 585342 439174
rect 585578 438938 585662 439174
rect 585898 438938 592650 439174
rect -8726 438854 592650 438938
rect -8726 438618 -1974 438854
rect -1738 438618 -1654 438854
rect -1418 438618 41746 438854
rect 41982 438618 42066 438854
rect 42302 438618 69746 438854
rect 69982 438618 70066 438854
rect 70302 438618 97746 438854
rect 97982 438618 98066 438854
rect 98302 438618 125746 438854
rect 125982 438618 126066 438854
rect 126302 438618 153746 438854
rect 153982 438618 154066 438854
rect 154302 438618 181746 438854
rect 181982 438618 182066 438854
rect 182302 438618 209746 438854
rect 209982 438618 210066 438854
rect 210302 438618 237746 438854
rect 237982 438618 238066 438854
rect 238302 438618 265746 438854
rect 265982 438618 266066 438854
rect 266302 438618 293746 438854
rect 293982 438618 294066 438854
rect 294302 438618 321746 438854
rect 321982 438618 322066 438854
rect 322302 438618 349746 438854
rect 349982 438618 350066 438854
rect 350302 438618 377746 438854
rect 377982 438618 378066 438854
rect 378302 438618 405746 438854
rect 405982 438618 406066 438854
rect 406302 438618 433746 438854
rect 433982 438618 434066 438854
rect 434302 438618 461746 438854
rect 461982 438618 462066 438854
rect 462302 438618 489746 438854
rect 489982 438618 490066 438854
rect 490302 438618 517746 438854
rect 517982 438618 518066 438854
rect 518302 438618 545746 438854
rect 545982 438618 546066 438854
rect 546302 438618 573746 438854
rect 573982 438618 574066 438854
rect 574302 438618 585342 438854
rect 585578 438618 585662 438854
rect 585898 438618 592650 438854
rect -8726 438586 592650 438618
rect -8726 435454 592650 435486
rect -8726 435218 -2934 435454
rect -2698 435218 -2614 435454
rect -2378 435218 38026 435454
rect 38262 435218 38346 435454
rect 38582 435218 66026 435454
rect 66262 435218 66346 435454
rect 66582 435218 94026 435454
rect 94262 435218 94346 435454
rect 94582 435218 122026 435454
rect 122262 435218 122346 435454
rect 122582 435218 150026 435454
rect 150262 435218 150346 435454
rect 150582 435218 178026 435454
rect 178262 435218 178346 435454
rect 178582 435218 206026 435454
rect 206262 435218 206346 435454
rect 206582 435218 234026 435454
rect 234262 435218 234346 435454
rect 234582 435218 262026 435454
rect 262262 435218 262346 435454
rect 262582 435218 290026 435454
rect 290262 435218 290346 435454
rect 290582 435218 318026 435454
rect 318262 435218 318346 435454
rect 318582 435218 346026 435454
rect 346262 435218 346346 435454
rect 346582 435218 374026 435454
rect 374262 435218 374346 435454
rect 374582 435218 402026 435454
rect 402262 435218 402346 435454
rect 402582 435218 430026 435454
rect 430262 435218 430346 435454
rect 430582 435218 458026 435454
rect 458262 435218 458346 435454
rect 458582 435218 486026 435454
rect 486262 435218 486346 435454
rect 486582 435218 514026 435454
rect 514262 435218 514346 435454
rect 514582 435218 542026 435454
rect 542262 435218 542346 435454
rect 542582 435218 570026 435454
rect 570262 435218 570346 435454
rect 570582 435218 586302 435454
rect 586538 435218 586622 435454
rect 586858 435218 592650 435454
rect -8726 435134 592650 435218
rect -8726 434898 -2934 435134
rect -2698 434898 -2614 435134
rect -2378 434898 38026 435134
rect 38262 434898 38346 435134
rect 38582 434898 66026 435134
rect 66262 434898 66346 435134
rect 66582 434898 94026 435134
rect 94262 434898 94346 435134
rect 94582 434898 122026 435134
rect 122262 434898 122346 435134
rect 122582 434898 150026 435134
rect 150262 434898 150346 435134
rect 150582 434898 178026 435134
rect 178262 434898 178346 435134
rect 178582 434898 206026 435134
rect 206262 434898 206346 435134
rect 206582 434898 234026 435134
rect 234262 434898 234346 435134
rect 234582 434898 262026 435134
rect 262262 434898 262346 435134
rect 262582 434898 290026 435134
rect 290262 434898 290346 435134
rect 290582 434898 318026 435134
rect 318262 434898 318346 435134
rect 318582 434898 346026 435134
rect 346262 434898 346346 435134
rect 346582 434898 374026 435134
rect 374262 434898 374346 435134
rect 374582 434898 402026 435134
rect 402262 434898 402346 435134
rect 402582 434898 430026 435134
rect 430262 434898 430346 435134
rect 430582 434898 458026 435134
rect 458262 434898 458346 435134
rect 458582 434898 486026 435134
rect 486262 434898 486346 435134
rect 486582 434898 514026 435134
rect 514262 434898 514346 435134
rect 514582 434898 542026 435134
rect 542262 434898 542346 435134
rect 542582 434898 570026 435134
rect 570262 434898 570346 435134
rect 570582 434898 586302 435134
rect 586538 434898 586622 435134
rect 586858 434898 592650 435134
rect -8726 434866 592650 434898
rect -8726 402174 592650 402206
rect -8726 401938 -1974 402174
rect -1738 401938 -1654 402174
rect -1418 401938 41746 402174
rect 41982 401938 42066 402174
rect 42302 401938 69746 402174
rect 69982 401938 70066 402174
rect 70302 401938 97746 402174
rect 97982 401938 98066 402174
rect 98302 401938 125746 402174
rect 125982 401938 126066 402174
rect 126302 401938 153746 402174
rect 153982 401938 154066 402174
rect 154302 401938 181746 402174
rect 181982 401938 182066 402174
rect 182302 401938 209746 402174
rect 209982 401938 210066 402174
rect 210302 401938 237746 402174
rect 237982 401938 238066 402174
rect 238302 401938 265746 402174
rect 265982 401938 266066 402174
rect 266302 401938 293746 402174
rect 293982 401938 294066 402174
rect 294302 401938 321746 402174
rect 321982 401938 322066 402174
rect 322302 401938 349746 402174
rect 349982 401938 350066 402174
rect 350302 401938 377746 402174
rect 377982 401938 378066 402174
rect 378302 401938 405746 402174
rect 405982 401938 406066 402174
rect 406302 401938 433746 402174
rect 433982 401938 434066 402174
rect 434302 401938 461746 402174
rect 461982 401938 462066 402174
rect 462302 401938 489746 402174
rect 489982 401938 490066 402174
rect 490302 401938 517746 402174
rect 517982 401938 518066 402174
rect 518302 401938 545746 402174
rect 545982 401938 546066 402174
rect 546302 401938 573746 402174
rect 573982 401938 574066 402174
rect 574302 401938 585342 402174
rect 585578 401938 585662 402174
rect 585898 401938 592650 402174
rect -8726 401854 592650 401938
rect -8726 401618 -1974 401854
rect -1738 401618 -1654 401854
rect -1418 401618 41746 401854
rect 41982 401618 42066 401854
rect 42302 401618 69746 401854
rect 69982 401618 70066 401854
rect 70302 401618 97746 401854
rect 97982 401618 98066 401854
rect 98302 401618 125746 401854
rect 125982 401618 126066 401854
rect 126302 401618 153746 401854
rect 153982 401618 154066 401854
rect 154302 401618 181746 401854
rect 181982 401618 182066 401854
rect 182302 401618 209746 401854
rect 209982 401618 210066 401854
rect 210302 401618 237746 401854
rect 237982 401618 238066 401854
rect 238302 401618 265746 401854
rect 265982 401618 266066 401854
rect 266302 401618 293746 401854
rect 293982 401618 294066 401854
rect 294302 401618 321746 401854
rect 321982 401618 322066 401854
rect 322302 401618 349746 401854
rect 349982 401618 350066 401854
rect 350302 401618 377746 401854
rect 377982 401618 378066 401854
rect 378302 401618 405746 401854
rect 405982 401618 406066 401854
rect 406302 401618 433746 401854
rect 433982 401618 434066 401854
rect 434302 401618 461746 401854
rect 461982 401618 462066 401854
rect 462302 401618 489746 401854
rect 489982 401618 490066 401854
rect 490302 401618 517746 401854
rect 517982 401618 518066 401854
rect 518302 401618 545746 401854
rect 545982 401618 546066 401854
rect 546302 401618 573746 401854
rect 573982 401618 574066 401854
rect 574302 401618 585342 401854
rect 585578 401618 585662 401854
rect 585898 401618 592650 401854
rect -8726 401586 592650 401618
rect -8726 398454 592650 398486
rect -8726 398218 -2934 398454
rect -2698 398218 -2614 398454
rect -2378 398218 38026 398454
rect 38262 398218 38346 398454
rect 38582 398218 66026 398454
rect 66262 398218 66346 398454
rect 66582 398218 94026 398454
rect 94262 398218 94346 398454
rect 94582 398218 122026 398454
rect 122262 398218 122346 398454
rect 122582 398218 150026 398454
rect 150262 398218 150346 398454
rect 150582 398218 178026 398454
rect 178262 398218 178346 398454
rect 178582 398218 206026 398454
rect 206262 398218 206346 398454
rect 206582 398218 234026 398454
rect 234262 398218 234346 398454
rect 234582 398218 262026 398454
rect 262262 398218 262346 398454
rect 262582 398218 290026 398454
rect 290262 398218 290346 398454
rect 290582 398218 318026 398454
rect 318262 398218 318346 398454
rect 318582 398218 346026 398454
rect 346262 398218 346346 398454
rect 346582 398218 374026 398454
rect 374262 398218 374346 398454
rect 374582 398218 402026 398454
rect 402262 398218 402346 398454
rect 402582 398218 430026 398454
rect 430262 398218 430346 398454
rect 430582 398218 458026 398454
rect 458262 398218 458346 398454
rect 458582 398218 486026 398454
rect 486262 398218 486346 398454
rect 486582 398218 514026 398454
rect 514262 398218 514346 398454
rect 514582 398218 542026 398454
rect 542262 398218 542346 398454
rect 542582 398218 570026 398454
rect 570262 398218 570346 398454
rect 570582 398218 586302 398454
rect 586538 398218 586622 398454
rect 586858 398218 592650 398454
rect -8726 398134 592650 398218
rect -8726 397898 -2934 398134
rect -2698 397898 -2614 398134
rect -2378 397898 38026 398134
rect 38262 397898 38346 398134
rect 38582 397898 66026 398134
rect 66262 397898 66346 398134
rect 66582 397898 94026 398134
rect 94262 397898 94346 398134
rect 94582 397898 122026 398134
rect 122262 397898 122346 398134
rect 122582 397898 150026 398134
rect 150262 397898 150346 398134
rect 150582 397898 178026 398134
rect 178262 397898 178346 398134
rect 178582 397898 206026 398134
rect 206262 397898 206346 398134
rect 206582 397898 234026 398134
rect 234262 397898 234346 398134
rect 234582 397898 262026 398134
rect 262262 397898 262346 398134
rect 262582 397898 290026 398134
rect 290262 397898 290346 398134
rect 290582 397898 318026 398134
rect 318262 397898 318346 398134
rect 318582 397898 346026 398134
rect 346262 397898 346346 398134
rect 346582 397898 374026 398134
rect 374262 397898 374346 398134
rect 374582 397898 402026 398134
rect 402262 397898 402346 398134
rect 402582 397898 430026 398134
rect 430262 397898 430346 398134
rect 430582 397898 458026 398134
rect 458262 397898 458346 398134
rect 458582 397898 486026 398134
rect 486262 397898 486346 398134
rect 486582 397898 514026 398134
rect 514262 397898 514346 398134
rect 514582 397898 542026 398134
rect 542262 397898 542346 398134
rect 542582 397898 570026 398134
rect 570262 397898 570346 398134
rect 570582 397898 586302 398134
rect 586538 397898 586622 398134
rect 586858 397898 592650 398134
rect -8726 397866 592650 397898
rect -8726 365174 592650 365206
rect -8726 364938 -1974 365174
rect -1738 364938 -1654 365174
rect -1418 364938 41746 365174
rect 41982 364938 42066 365174
rect 42302 364938 69746 365174
rect 69982 364938 70066 365174
rect 70302 364938 97746 365174
rect 97982 364938 98066 365174
rect 98302 364938 125746 365174
rect 125982 364938 126066 365174
rect 126302 364938 153746 365174
rect 153982 364938 154066 365174
rect 154302 364938 181746 365174
rect 181982 364938 182066 365174
rect 182302 364938 209746 365174
rect 209982 364938 210066 365174
rect 210302 364938 237746 365174
rect 237982 364938 238066 365174
rect 238302 364938 265746 365174
rect 265982 364938 266066 365174
rect 266302 364938 293746 365174
rect 293982 364938 294066 365174
rect 294302 364938 321746 365174
rect 321982 364938 322066 365174
rect 322302 364938 349746 365174
rect 349982 364938 350066 365174
rect 350302 364938 377746 365174
rect 377982 364938 378066 365174
rect 378302 364938 405746 365174
rect 405982 364938 406066 365174
rect 406302 364938 433746 365174
rect 433982 364938 434066 365174
rect 434302 364938 461746 365174
rect 461982 364938 462066 365174
rect 462302 364938 489746 365174
rect 489982 364938 490066 365174
rect 490302 364938 517746 365174
rect 517982 364938 518066 365174
rect 518302 364938 545746 365174
rect 545982 364938 546066 365174
rect 546302 364938 573746 365174
rect 573982 364938 574066 365174
rect 574302 364938 585342 365174
rect 585578 364938 585662 365174
rect 585898 364938 592650 365174
rect -8726 364854 592650 364938
rect -8726 364618 -1974 364854
rect -1738 364618 -1654 364854
rect -1418 364618 41746 364854
rect 41982 364618 42066 364854
rect 42302 364618 69746 364854
rect 69982 364618 70066 364854
rect 70302 364618 97746 364854
rect 97982 364618 98066 364854
rect 98302 364618 125746 364854
rect 125982 364618 126066 364854
rect 126302 364618 153746 364854
rect 153982 364618 154066 364854
rect 154302 364618 181746 364854
rect 181982 364618 182066 364854
rect 182302 364618 209746 364854
rect 209982 364618 210066 364854
rect 210302 364618 237746 364854
rect 237982 364618 238066 364854
rect 238302 364618 265746 364854
rect 265982 364618 266066 364854
rect 266302 364618 293746 364854
rect 293982 364618 294066 364854
rect 294302 364618 321746 364854
rect 321982 364618 322066 364854
rect 322302 364618 349746 364854
rect 349982 364618 350066 364854
rect 350302 364618 377746 364854
rect 377982 364618 378066 364854
rect 378302 364618 405746 364854
rect 405982 364618 406066 364854
rect 406302 364618 433746 364854
rect 433982 364618 434066 364854
rect 434302 364618 461746 364854
rect 461982 364618 462066 364854
rect 462302 364618 489746 364854
rect 489982 364618 490066 364854
rect 490302 364618 517746 364854
rect 517982 364618 518066 364854
rect 518302 364618 545746 364854
rect 545982 364618 546066 364854
rect 546302 364618 573746 364854
rect 573982 364618 574066 364854
rect 574302 364618 585342 364854
rect 585578 364618 585662 364854
rect 585898 364618 592650 364854
rect -8726 364586 592650 364618
rect -8726 361454 592650 361486
rect -8726 361218 -2934 361454
rect -2698 361218 -2614 361454
rect -2378 361218 38026 361454
rect 38262 361218 38346 361454
rect 38582 361218 66026 361454
rect 66262 361218 66346 361454
rect 66582 361218 94026 361454
rect 94262 361218 94346 361454
rect 94582 361218 122026 361454
rect 122262 361218 122346 361454
rect 122582 361218 150026 361454
rect 150262 361218 150346 361454
rect 150582 361218 178026 361454
rect 178262 361218 178346 361454
rect 178582 361218 206026 361454
rect 206262 361218 206346 361454
rect 206582 361218 234026 361454
rect 234262 361218 234346 361454
rect 234582 361218 262026 361454
rect 262262 361218 262346 361454
rect 262582 361218 290026 361454
rect 290262 361218 290346 361454
rect 290582 361218 318026 361454
rect 318262 361218 318346 361454
rect 318582 361218 346026 361454
rect 346262 361218 346346 361454
rect 346582 361218 374026 361454
rect 374262 361218 374346 361454
rect 374582 361218 402026 361454
rect 402262 361218 402346 361454
rect 402582 361218 430026 361454
rect 430262 361218 430346 361454
rect 430582 361218 458026 361454
rect 458262 361218 458346 361454
rect 458582 361218 486026 361454
rect 486262 361218 486346 361454
rect 486582 361218 514026 361454
rect 514262 361218 514346 361454
rect 514582 361218 542026 361454
rect 542262 361218 542346 361454
rect 542582 361218 570026 361454
rect 570262 361218 570346 361454
rect 570582 361218 586302 361454
rect 586538 361218 586622 361454
rect 586858 361218 592650 361454
rect -8726 361134 592650 361218
rect -8726 360898 -2934 361134
rect -2698 360898 -2614 361134
rect -2378 360898 38026 361134
rect 38262 360898 38346 361134
rect 38582 360898 66026 361134
rect 66262 360898 66346 361134
rect 66582 360898 94026 361134
rect 94262 360898 94346 361134
rect 94582 360898 122026 361134
rect 122262 360898 122346 361134
rect 122582 360898 150026 361134
rect 150262 360898 150346 361134
rect 150582 360898 178026 361134
rect 178262 360898 178346 361134
rect 178582 360898 206026 361134
rect 206262 360898 206346 361134
rect 206582 360898 234026 361134
rect 234262 360898 234346 361134
rect 234582 360898 262026 361134
rect 262262 360898 262346 361134
rect 262582 360898 290026 361134
rect 290262 360898 290346 361134
rect 290582 360898 318026 361134
rect 318262 360898 318346 361134
rect 318582 360898 346026 361134
rect 346262 360898 346346 361134
rect 346582 360898 374026 361134
rect 374262 360898 374346 361134
rect 374582 360898 402026 361134
rect 402262 360898 402346 361134
rect 402582 360898 430026 361134
rect 430262 360898 430346 361134
rect 430582 360898 458026 361134
rect 458262 360898 458346 361134
rect 458582 360898 486026 361134
rect 486262 360898 486346 361134
rect 486582 360898 514026 361134
rect 514262 360898 514346 361134
rect 514582 360898 542026 361134
rect 542262 360898 542346 361134
rect 542582 360898 570026 361134
rect 570262 360898 570346 361134
rect 570582 360898 586302 361134
rect 586538 360898 586622 361134
rect 586858 360898 592650 361134
rect -8726 360866 592650 360898
rect -8726 328174 592650 328206
rect -8726 327938 -1974 328174
rect -1738 327938 -1654 328174
rect -1418 327938 41746 328174
rect 41982 327938 42066 328174
rect 42302 327938 69746 328174
rect 69982 327938 70066 328174
rect 70302 327938 97746 328174
rect 97982 327938 98066 328174
rect 98302 327938 125746 328174
rect 125982 327938 126066 328174
rect 126302 327938 153746 328174
rect 153982 327938 154066 328174
rect 154302 327938 181746 328174
rect 181982 327938 182066 328174
rect 182302 327938 209746 328174
rect 209982 327938 210066 328174
rect 210302 327938 237746 328174
rect 237982 327938 238066 328174
rect 238302 327938 265746 328174
rect 265982 327938 266066 328174
rect 266302 327938 293746 328174
rect 293982 327938 294066 328174
rect 294302 327938 321746 328174
rect 321982 327938 322066 328174
rect 322302 327938 349746 328174
rect 349982 327938 350066 328174
rect 350302 327938 377746 328174
rect 377982 327938 378066 328174
rect 378302 327938 405746 328174
rect 405982 327938 406066 328174
rect 406302 327938 433746 328174
rect 433982 327938 434066 328174
rect 434302 327938 461746 328174
rect 461982 327938 462066 328174
rect 462302 327938 489746 328174
rect 489982 327938 490066 328174
rect 490302 327938 517746 328174
rect 517982 327938 518066 328174
rect 518302 327938 545746 328174
rect 545982 327938 546066 328174
rect 546302 327938 573746 328174
rect 573982 327938 574066 328174
rect 574302 327938 585342 328174
rect 585578 327938 585662 328174
rect 585898 327938 592650 328174
rect -8726 327854 592650 327938
rect -8726 327618 -1974 327854
rect -1738 327618 -1654 327854
rect -1418 327618 41746 327854
rect 41982 327618 42066 327854
rect 42302 327618 69746 327854
rect 69982 327618 70066 327854
rect 70302 327618 97746 327854
rect 97982 327618 98066 327854
rect 98302 327618 125746 327854
rect 125982 327618 126066 327854
rect 126302 327618 153746 327854
rect 153982 327618 154066 327854
rect 154302 327618 181746 327854
rect 181982 327618 182066 327854
rect 182302 327618 209746 327854
rect 209982 327618 210066 327854
rect 210302 327618 237746 327854
rect 237982 327618 238066 327854
rect 238302 327618 265746 327854
rect 265982 327618 266066 327854
rect 266302 327618 293746 327854
rect 293982 327618 294066 327854
rect 294302 327618 321746 327854
rect 321982 327618 322066 327854
rect 322302 327618 349746 327854
rect 349982 327618 350066 327854
rect 350302 327618 377746 327854
rect 377982 327618 378066 327854
rect 378302 327618 405746 327854
rect 405982 327618 406066 327854
rect 406302 327618 433746 327854
rect 433982 327618 434066 327854
rect 434302 327618 461746 327854
rect 461982 327618 462066 327854
rect 462302 327618 489746 327854
rect 489982 327618 490066 327854
rect 490302 327618 517746 327854
rect 517982 327618 518066 327854
rect 518302 327618 545746 327854
rect 545982 327618 546066 327854
rect 546302 327618 573746 327854
rect 573982 327618 574066 327854
rect 574302 327618 585342 327854
rect 585578 327618 585662 327854
rect 585898 327618 592650 327854
rect -8726 327586 592650 327618
rect -8726 324454 592650 324486
rect -8726 324218 -2934 324454
rect -2698 324218 -2614 324454
rect -2378 324218 38026 324454
rect 38262 324218 38346 324454
rect 38582 324218 66026 324454
rect 66262 324218 66346 324454
rect 66582 324218 94026 324454
rect 94262 324218 94346 324454
rect 94582 324218 122026 324454
rect 122262 324218 122346 324454
rect 122582 324218 150026 324454
rect 150262 324218 150346 324454
rect 150582 324218 178026 324454
rect 178262 324218 178346 324454
rect 178582 324218 206026 324454
rect 206262 324218 206346 324454
rect 206582 324218 234026 324454
rect 234262 324218 234346 324454
rect 234582 324218 262026 324454
rect 262262 324218 262346 324454
rect 262582 324218 290026 324454
rect 290262 324218 290346 324454
rect 290582 324218 318026 324454
rect 318262 324218 318346 324454
rect 318582 324218 346026 324454
rect 346262 324218 346346 324454
rect 346582 324218 374026 324454
rect 374262 324218 374346 324454
rect 374582 324218 402026 324454
rect 402262 324218 402346 324454
rect 402582 324218 430026 324454
rect 430262 324218 430346 324454
rect 430582 324218 458026 324454
rect 458262 324218 458346 324454
rect 458582 324218 486026 324454
rect 486262 324218 486346 324454
rect 486582 324218 514026 324454
rect 514262 324218 514346 324454
rect 514582 324218 542026 324454
rect 542262 324218 542346 324454
rect 542582 324218 570026 324454
rect 570262 324218 570346 324454
rect 570582 324218 586302 324454
rect 586538 324218 586622 324454
rect 586858 324218 592650 324454
rect -8726 324134 592650 324218
rect -8726 323898 -2934 324134
rect -2698 323898 -2614 324134
rect -2378 323898 38026 324134
rect 38262 323898 38346 324134
rect 38582 323898 66026 324134
rect 66262 323898 66346 324134
rect 66582 323898 94026 324134
rect 94262 323898 94346 324134
rect 94582 323898 122026 324134
rect 122262 323898 122346 324134
rect 122582 323898 150026 324134
rect 150262 323898 150346 324134
rect 150582 323898 178026 324134
rect 178262 323898 178346 324134
rect 178582 323898 206026 324134
rect 206262 323898 206346 324134
rect 206582 323898 234026 324134
rect 234262 323898 234346 324134
rect 234582 323898 262026 324134
rect 262262 323898 262346 324134
rect 262582 323898 290026 324134
rect 290262 323898 290346 324134
rect 290582 323898 318026 324134
rect 318262 323898 318346 324134
rect 318582 323898 346026 324134
rect 346262 323898 346346 324134
rect 346582 323898 374026 324134
rect 374262 323898 374346 324134
rect 374582 323898 402026 324134
rect 402262 323898 402346 324134
rect 402582 323898 430026 324134
rect 430262 323898 430346 324134
rect 430582 323898 458026 324134
rect 458262 323898 458346 324134
rect 458582 323898 486026 324134
rect 486262 323898 486346 324134
rect 486582 323898 514026 324134
rect 514262 323898 514346 324134
rect 514582 323898 542026 324134
rect 542262 323898 542346 324134
rect 542582 323898 570026 324134
rect 570262 323898 570346 324134
rect 570582 323898 586302 324134
rect 586538 323898 586622 324134
rect 586858 323898 592650 324134
rect -8726 323866 592650 323898
rect -8726 291174 592650 291206
rect -8726 290938 -1974 291174
rect -1738 290938 -1654 291174
rect -1418 290938 41746 291174
rect 41982 290938 42066 291174
rect 42302 290938 69746 291174
rect 69982 290938 70066 291174
rect 70302 290938 97746 291174
rect 97982 290938 98066 291174
rect 98302 290938 125746 291174
rect 125982 290938 126066 291174
rect 126302 290938 153746 291174
rect 153982 290938 154066 291174
rect 154302 290938 181746 291174
rect 181982 290938 182066 291174
rect 182302 290938 209746 291174
rect 209982 290938 210066 291174
rect 210302 290938 237746 291174
rect 237982 290938 238066 291174
rect 238302 290938 265746 291174
rect 265982 290938 266066 291174
rect 266302 290938 293746 291174
rect 293982 290938 294066 291174
rect 294302 290938 321746 291174
rect 321982 290938 322066 291174
rect 322302 290938 349746 291174
rect 349982 290938 350066 291174
rect 350302 290938 377746 291174
rect 377982 290938 378066 291174
rect 378302 290938 405746 291174
rect 405982 290938 406066 291174
rect 406302 290938 433746 291174
rect 433982 290938 434066 291174
rect 434302 290938 461746 291174
rect 461982 290938 462066 291174
rect 462302 290938 489746 291174
rect 489982 290938 490066 291174
rect 490302 290938 517746 291174
rect 517982 290938 518066 291174
rect 518302 290938 545746 291174
rect 545982 290938 546066 291174
rect 546302 290938 573746 291174
rect 573982 290938 574066 291174
rect 574302 290938 585342 291174
rect 585578 290938 585662 291174
rect 585898 290938 592650 291174
rect -8726 290854 592650 290938
rect -8726 290618 -1974 290854
rect -1738 290618 -1654 290854
rect -1418 290618 41746 290854
rect 41982 290618 42066 290854
rect 42302 290618 69746 290854
rect 69982 290618 70066 290854
rect 70302 290618 97746 290854
rect 97982 290618 98066 290854
rect 98302 290618 125746 290854
rect 125982 290618 126066 290854
rect 126302 290618 153746 290854
rect 153982 290618 154066 290854
rect 154302 290618 181746 290854
rect 181982 290618 182066 290854
rect 182302 290618 209746 290854
rect 209982 290618 210066 290854
rect 210302 290618 237746 290854
rect 237982 290618 238066 290854
rect 238302 290618 265746 290854
rect 265982 290618 266066 290854
rect 266302 290618 293746 290854
rect 293982 290618 294066 290854
rect 294302 290618 321746 290854
rect 321982 290618 322066 290854
rect 322302 290618 349746 290854
rect 349982 290618 350066 290854
rect 350302 290618 377746 290854
rect 377982 290618 378066 290854
rect 378302 290618 405746 290854
rect 405982 290618 406066 290854
rect 406302 290618 433746 290854
rect 433982 290618 434066 290854
rect 434302 290618 461746 290854
rect 461982 290618 462066 290854
rect 462302 290618 489746 290854
rect 489982 290618 490066 290854
rect 490302 290618 517746 290854
rect 517982 290618 518066 290854
rect 518302 290618 545746 290854
rect 545982 290618 546066 290854
rect 546302 290618 573746 290854
rect 573982 290618 574066 290854
rect 574302 290618 585342 290854
rect 585578 290618 585662 290854
rect 585898 290618 592650 290854
rect -8726 290586 592650 290618
rect -8726 287454 592650 287486
rect -8726 287218 -2934 287454
rect -2698 287218 -2614 287454
rect -2378 287218 38026 287454
rect 38262 287218 38346 287454
rect 38582 287218 66026 287454
rect 66262 287218 66346 287454
rect 66582 287218 94026 287454
rect 94262 287218 94346 287454
rect 94582 287218 122026 287454
rect 122262 287218 122346 287454
rect 122582 287218 150026 287454
rect 150262 287218 150346 287454
rect 150582 287218 178026 287454
rect 178262 287218 178346 287454
rect 178582 287218 206026 287454
rect 206262 287218 206346 287454
rect 206582 287218 234026 287454
rect 234262 287218 234346 287454
rect 234582 287218 262026 287454
rect 262262 287218 262346 287454
rect 262582 287218 290026 287454
rect 290262 287218 290346 287454
rect 290582 287218 318026 287454
rect 318262 287218 318346 287454
rect 318582 287218 346026 287454
rect 346262 287218 346346 287454
rect 346582 287218 374026 287454
rect 374262 287218 374346 287454
rect 374582 287218 402026 287454
rect 402262 287218 402346 287454
rect 402582 287218 430026 287454
rect 430262 287218 430346 287454
rect 430582 287218 458026 287454
rect 458262 287218 458346 287454
rect 458582 287218 486026 287454
rect 486262 287218 486346 287454
rect 486582 287218 514026 287454
rect 514262 287218 514346 287454
rect 514582 287218 542026 287454
rect 542262 287218 542346 287454
rect 542582 287218 570026 287454
rect 570262 287218 570346 287454
rect 570582 287218 586302 287454
rect 586538 287218 586622 287454
rect 586858 287218 592650 287454
rect -8726 287134 592650 287218
rect -8726 286898 -2934 287134
rect -2698 286898 -2614 287134
rect -2378 286898 38026 287134
rect 38262 286898 38346 287134
rect 38582 286898 66026 287134
rect 66262 286898 66346 287134
rect 66582 286898 94026 287134
rect 94262 286898 94346 287134
rect 94582 286898 122026 287134
rect 122262 286898 122346 287134
rect 122582 286898 150026 287134
rect 150262 286898 150346 287134
rect 150582 286898 178026 287134
rect 178262 286898 178346 287134
rect 178582 286898 206026 287134
rect 206262 286898 206346 287134
rect 206582 286898 234026 287134
rect 234262 286898 234346 287134
rect 234582 286898 262026 287134
rect 262262 286898 262346 287134
rect 262582 286898 290026 287134
rect 290262 286898 290346 287134
rect 290582 286898 318026 287134
rect 318262 286898 318346 287134
rect 318582 286898 346026 287134
rect 346262 286898 346346 287134
rect 346582 286898 374026 287134
rect 374262 286898 374346 287134
rect 374582 286898 402026 287134
rect 402262 286898 402346 287134
rect 402582 286898 430026 287134
rect 430262 286898 430346 287134
rect 430582 286898 458026 287134
rect 458262 286898 458346 287134
rect 458582 286898 486026 287134
rect 486262 286898 486346 287134
rect 486582 286898 514026 287134
rect 514262 286898 514346 287134
rect 514582 286898 542026 287134
rect 542262 286898 542346 287134
rect 542582 286898 570026 287134
rect 570262 286898 570346 287134
rect 570582 286898 586302 287134
rect 586538 286898 586622 287134
rect 586858 286898 592650 287134
rect -8726 286866 592650 286898
rect -8726 254174 592650 254206
rect -8726 253938 -1974 254174
rect -1738 253938 -1654 254174
rect -1418 253938 41746 254174
rect 41982 253938 42066 254174
rect 42302 253938 69746 254174
rect 69982 253938 70066 254174
rect 70302 253938 97746 254174
rect 97982 253938 98066 254174
rect 98302 253938 125746 254174
rect 125982 253938 126066 254174
rect 126302 253938 153746 254174
rect 153982 253938 154066 254174
rect 154302 253938 181746 254174
rect 181982 253938 182066 254174
rect 182302 253938 209746 254174
rect 209982 253938 210066 254174
rect 210302 253938 237746 254174
rect 237982 253938 238066 254174
rect 238302 253938 265746 254174
rect 265982 253938 266066 254174
rect 266302 253938 293746 254174
rect 293982 253938 294066 254174
rect 294302 253938 321746 254174
rect 321982 253938 322066 254174
rect 322302 253938 349746 254174
rect 349982 253938 350066 254174
rect 350302 253938 377746 254174
rect 377982 253938 378066 254174
rect 378302 253938 405746 254174
rect 405982 253938 406066 254174
rect 406302 253938 433746 254174
rect 433982 253938 434066 254174
rect 434302 253938 461746 254174
rect 461982 253938 462066 254174
rect 462302 253938 489746 254174
rect 489982 253938 490066 254174
rect 490302 253938 517746 254174
rect 517982 253938 518066 254174
rect 518302 253938 545746 254174
rect 545982 253938 546066 254174
rect 546302 253938 573746 254174
rect 573982 253938 574066 254174
rect 574302 253938 585342 254174
rect 585578 253938 585662 254174
rect 585898 253938 592650 254174
rect -8726 253854 592650 253938
rect -8726 253618 -1974 253854
rect -1738 253618 -1654 253854
rect -1418 253618 41746 253854
rect 41982 253618 42066 253854
rect 42302 253618 69746 253854
rect 69982 253618 70066 253854
rect 70302 253618 97746 253854
rect 97982 253618 98066 253854
rect 98302 253618 125746 253854
rect 125982 253618 126066 253854
rect 126302 253618 153746 253854
rect 153982 253618 154066 253854
rect 154302 253618 181746 253854
rect 181982 253618 182066 253854
rect 182302 253618 209746 253854
rect 209982 253618 210066 253854
rect 210302 253618 237746 253854
rect 237982 253618 238066 253854
rect 238302 253618 265746 253854
rect 265982 253618 266066 253854
rect 266302 253618 293746 253854
rect 293982 253618 294066 253854
rect 294302 253618 321746 253854
rect 321982 253618 322066 253854
rect 322302 253618 349746 253854
rect 349982 253618 350066 253854
rect 350302 253618 377746 253854
rect 377982 253618 378066 253854
rect 378302 253618 405746 253854
rect 405982 253618 406066 253854
rect 406302 253618 433746 253854
rect 433982 253618 434066 253854
rect 434302 253618 461746 253854
rect 461982 253618 462066 253854
rect 462302 253618 489746 253854
rect 489982 253618 490066 253854
rect 490302 253618 517746 253854
rect 517982 253618 518066 253854
rect 518302 253618 545746 253854
rect 545982 253618 546066 253854
rect 546302 253618 573746 253854
rect 573982 253618 574066 253854
rect 574302 253618 585342 253854
rect 585578 253618 585662 253854
rect 585898 253618 592650 253854
rect -8726 253586 592650 253618
rect -8726 250454 592650 250486
rect -8726 250218 -2934 250454
rect -2698 250218 -2614 250454
rect -2378 250218 38026 250454
rect 38262 250218 38346 250454
rect 38582 250218 66026 250454
rect 66262 250218 66346 250454
rect 66582 250218 94026 250454
rect 94262 250218 94346 250454
rect 94582 250218 122026 250454
rect 122262 250218 122346 250454
rect 122582 250218 150026 250454
rect 150262 250218 150346 250454
rect 150582 250218 178026 250454
rect 178262 250218 178346 250454
rect 178582 250218 206026 250454
rect 206262 250218 206346 250454
rect 206582 250218 234026 250454
rect 234262 250218 234346 250454
rect 234582 250218 262026 250454
rect 262262 250218 262346 250454
rect 262582 250218 290026 250454
rect 290262 250218 290346 250454
rect 290582 250218 318026 250454
rect 318262 250218 318346 250454
rect 318582 250218 346026 250454
rect 346262 250218 346346 250454
rect 346582 250218 374026 250454
rect 374262 250218 374346 250454
rect 374582 250218 402026 250454
rect 402262 250218 402346 250454
rect 402582 250218 430026 250454
rect 430262 250218 430346 250454
rect 430582 250218 458026 250454
rect 458262 250218 458346 250454
rect 458582 250218 486026 250454
rect 486262 250218 486346 250454
rect 486582 250218 514026 250454
rect 514262 250218 514346 250454
rect 514582 250218 542026 250454
rect 542262 250218 542346 250454
rect 542582 250218 570026 250454
rect 570262 250218 570346 250454
rect 570582 250218 586302 250454
rect 586538 250218 586622 250454
rect 586858 250218 592650 250454
rect -8726 250134 592650 250218
rect -8726 249898 -2934 250134
rect -2698 249898 -2614 250134
rect -2378 249898 38026 250134
rect 38262 249898 38346 250134
rect 38582 249898 66026 250134
rect 66262 249898 66346 250134
rect 66582 249898 94026 250134
rect 94262 249898 94346 250134
rect 94582 249898 122026 250134
rect 122262 249898 122346 250134
rect 122582 249898 150026 250134
rect 150262 249898 150346 250134
rect 150582 249898 178026 250134
rect 178262 249898 178346 250134
rect 178582 249898 206026 250134
rect 206262 249898 206346 250134
rect 206582 249898 234026 250134
rect 234262 249898 234346 250134
rect 234582 249898 262026 250134
rect 262262 249898 262346 250134
rect 262582 249898 290026 250134
rect 290262 249898 290346 250134
rect 290582 249898 318026 250134
rect 318262 249898 318346 250134
rect 318582 249898 346026 250134
rect 346262 249898 346346 250134
rect 346582 249898 374026 250134
rect 374262 249898 374346 250134
rect 374582 249898 402026 250134
rect 402262 249898 402346 250134
rect 402582 249898 430026 250134
rect 430262 249898 430346 250134
rect 430582 249898 458026 250134
rect 458262 249898 458346 250134
rect 458582 249898 486026 250134
rect 486262 249898 486346 250134
rect 486582 249898 514026 250134
rect 514262 249898 514346 250134
rect 514582 249898 542026 250134
rect 542262 249898 542346 250134
rect 542582 249898 570026 250134
rect 570262 249898 570346 250134
rect 570582 249898 586302 250134
rect 586538 249898 586622 250134
rect 586858 249898 592650 250134
rect -8726 249866 592650 249898
rect -8726 217174 592650 217206
rect -8726 216938 -1974 217174
rect -1738 216938 -1654 217174
rect -1418 216938 41746 217174
rect 41982 216938 42066 217174
rect 42302 216938 69746 217174
rect 69982 216938 70066 217174
rect 70302 216938 97746 217174
rect 97982 216938 98066 217174
rect 98302 216938 125746 217174
rect 125982 216938 126066 217174
rect 126302 216938 153746 217174
rect 153982 216938 154066 217174
rect 154302 216938 181746 217174
rect 181982 216938 182066 217174
rect 182302 216938 209746 217174
rect 209982 216938 210066 217174
rect 210302 216938 237746 217174
rect 237982 216938 238066 217174
rect 238302 216938 265746 217174
rect 265982 216938 266066 217174
rect 266302 216938 293746 217174
rect 293982 216938 294066 217174
rect 294302 216938 321746 217174
rect 321982 216938 322066 217174
rect 322302 216938 349746 217174
rect 349982 216938 350066 217174
rect 350302 216938 377746 217174
rect 377982 216938 378066 217174
rect 378302 216938 405746 217174
rect 405982 216938 406066 217174
rect 406302 216938 433746 217174
rect 433982 216938 434066 217174
rect 434302 216938 461746 217174
rect 461982 216938 462066 217174
rect 462302 216938 489746 217174
rect 489982 216938 490066 217174
rect 490302 216938 517746 217174
rect 517982 216938 518066 217174
rect 518302 216938 545746 217174
rect 545982 216938 546066 217174
rect 546302 216938 573746 217174
rect 573982 216938 574066 217174
rect 574302 216938 585342 217174
rect 585578 216938 585662 217174
rect 585898 216938 592650 217174
rect -8726 216854 592650 216938
rect -8726 216618 -1974 216854
rect -1738 216618 -1654 216854
rect -1418 216618 41746 216854
rect 41982 216618 42066 216854
rect 42302 216618 69746 216854
rect 69982 216618 70066 216854
rect 70302 216618 97746 216854
rect 97982 216618 98066 216854
rect 98302 216618 125746 216854
rect 125982 216618 126066 216854
rect 126302 216618 153746 216854
rect 153982 216618 154066 216854
rect 154302 216618 181746 216854
rect 181982 216618 182066 216854
rect 182302 216618 209746 216854
rect 209982 216618 210066 216854
rect 210302 216618 237746 216854
rect 237982 216618 238066 216854
rect 238302 216618 265746 216854
rect 265982 216618 266066 216854
rect 266302 216618 293746 216854
rect 293982 216618 294066 216854
rect 294302 216618 321746 216854
rect 321982 216618 322066 216854
rect 322302 216618 349746 216854
rect 349982 216618 350066 216854
rect 350302 216618 377746 216854
rect 377982 216618 378066 216854
rect 378302 216618 405746 216854
rect 405982 216618 406066 216854
rect 406302 216618 433746 216854
rect 433982 216618 434066 216854
rect 434302 216618 461746 216854
rect 461982 216618 462066 216854
rect 462302 216618 489746 216854
rect 489982 216618 490066 216854
rect 490302 216618 517746 216854
rect 517982 216618 518066 216854
rect 518302 216618 545746 216854
rect 545982 216618 546066 216854
rect 546302 216618 573746 216854
rect 573982 216618 574066 216854
rect 574302 216618 585342 216854
rect 585578 216618 585662 216854
rect 585898 216618 592650 216854
rect -8726 216586 592650 216618
rect -8726 213454 592650 213486
rect -8726 213218 -2934 213454
rect -2698 213218 -2614 213454
rect -2378 213218 38026 213454
rect 38262 213218 38346 213454
rect 38582 213218 66026 213454
rect 66262 213218 66346 213454
rect 66582 213218 94026 213454
rect 94262 213218 94346 213454
rect 94582 213218 122026 213454
rect 122262 213218 122346 213454
rect 122582 213218 150026 213454
rect 150262 213218 150346 213454
rect 150582 213218 178026 213454
rect 178262 213218 178346 213454
rect 178582 213218 206026 213454
rect 206262 213218 206346 213454
rect 206582 213218 234026 213454
rect 234262 213218 234346 213454
rect 234582 213218 262026 213454
rect 262262 213218 262346 213454
rect 262582 213218 290026 213454
rect 290262 213218 290346 213454
rect 290582 213218 318026 213454
rect 318262 213218 318346 213454
rect 318582 213218 346026 213454
rect 346262 213218 346346 213454
rect 346582 213218 374026 213454
rect 374262 213218 374346 213454
rect 374582 213218 402026 213454
rect 402262 213218 402346 213454
rect 402582 213218 430026 213454
rect 430262 213218 430346 213454
rect 430582 213218 458026 213454
rect 458262 213218 458346 213454
rect 458582 213218 486026 213454
rect 486262 213218 486346 213454
rect 486582 213218 514026 213454
rect 514262 213218 514346 213454
rect 514582 213218 542026 213454
rect 542262 213218 542346 213454
rect 542582 213218 570026 213454
rect 570262 213218 570346 213454
rect 570582 213218 586302 213454
rect 586538 213218 586622 213454
rect 586858 213218 592650 213454
rect -8726 213134 592650 213218
rect -8726 212898 -2934 213134
rect -2698 212898 -2614 213134
rect -2378 212898 38026 213134
rect 38262 212898 38346 213134
rect 38582 212898 66026 213134
rect 66262 212898 66346 213134
rect 66582 212898 94026 213134
rect 94262 212898 94346 213134
rect 94582 212898 122026 213134
rect 122262 212898 122346 213134
rect 122582 212898 150026 213134
rect 150262 212898 150346 213134
rect 150582 212898 178026 213134
rect 178262 212898 178346 213134
rect 178582 212898 206026 213134
rect 206262 212898 206346 213134
rect 206582 212898 234026 213134
rect 234262 212898 234346 213134
rect 234582 212898 262026 213134
rect 262262 212898 262346 213134
rect 262582 212898 290026 213134
rect 290262 212898 290346 213134
rect 290582 212898 318026 213134
rect 318262 212898 318346 213134
rect 318582 212898 346026 213134
rect 346262 212898 346346 213134
rect 346582 212898 374026 213134
rect 374262 212898 374346 213134
rect 374582 212898 402026 213134
rect 402262 212898 402346 213134
rect 402582 212898 430026 213134
rect 430262 212898 430346 213134
rect 430582 212898 458026 213134
rect 458262 212898 458346 213134
rect 458582 212898 486026 213134
rect 486262 212898 486346 213134
rect 486582 212898 514026 213134
rect 514262 212898 514346 213134
rect 514582 212898 542026 213134
rect 542262 212898 542346 213134
rect 542582 212898 570026 213134
rect 570262 212898 570346 213134
rect 570582 212898 586302 213134
rect 586538 212898 586622 213134
rect 586858 212898 592650 213134
rect -8726 212866 592650 212898
rect -8726 180174 592650 180206
rect -8726 179938 -1974 180174
rect -1738 179938 -1654 180174
rect -1418 179938 41746 180174
rect 41982 179938 42066 180174
rect 42302 179938 69746 180174
rect 69982 179938 70066 180174
rect 70302 179938 97746 180174
rect 97982 179938 98066 180174
rect 98302 179938 125746 180174
rect 125982 179938 126066 180174
rect 126302 179938 153746 180174
rect 153982 179938 154066 180174
rect 154302 179938 181746 180174
rect 181982 179938 182066 180174
rect 182302 179938 209746 180174
rect 209982 179938 210066 180174
rect 210302 179938 237746 180174
rect 237982 179938 238066 180174
rect 238302 179938 265746 180174
rect 265982 179938 266066 180174
rect 266302 179938 293746 180174
rect 293982 179938 294066 180174
rect 294302 179938 321746 180174
rect 321982 179938 322066 180174
rect 322302 179938 349746 180174
rect 349982 179938 350066 180174
rect 350302 179938 377746 180174
rect 377982 179938 378066 180174
rect 378302 179938 405746 180174
rect 405982 179938 406066 180174
rect 406302 179938 433746 180174
rect 433982 179938 434066 180174
rect 434302 179938 461746 180174
rect 461982 179938 462066 180174
rect 462302 179938 489746 180174
rect 489982 179938 490066 180174
rect 490302 179938 517746 180174
rect 517982 179938 518066 180174
rect 518302 179938 545746 180174
rect 545982 179938 546066 180174
rect 546302 179938 573746 180174
rect 573982 179938 574066 180174
rect 574302 179938 585342 180174
rect 585578 179938 585662 180174
rect 585898 179938 592650 180174
rect -8726 179854 592650 179938
rect -8726 179618 -1974 179854
rect -1738 179618 -1654 179854
rect -1418 179618 41746 179854
rect 41982 179618 42066 179854
rect 42302 179618 69746 179854
rect 69982 179618 70066 179854
rect 70302 179618 97746 179854
rect 97982 179618 98066 179854
rect 98302 179618 125746 179854
rect 125982 179618 126066 179854
rect 126302 179618 153746 179854
rect 153982 179618 154066 179854
rect 154302 179618 181746 179854
rect 181982 179618 182066 179854
rect 182302 179618 209746 179854
rect 209982 179618 210066 179854
rect 210302 179618 237746 179854
rect 237982 179618 238066 179854
rect 238302 179618 265746 179854
rect 265982 179618 266066 179854
rect 266302 179618 293746 179854
rect 293982 179618 294066 179854
rect 294302 179618 321746 179854
rect 321982 179618 322066 179854
rect 322302 179618 349746 179854
rect 349982 179618 350066 179854
rect 350302 179618 377746 179854
rect 377982 179618 378066 179854
rect 378302 179618 405746 179854
rect 405982 179618 406066 179854
rect 406302 179618 433746 179854
rect 433982 179618 434066 179854
rect 434302 179618 461746 179854
rect 461982 179618 462066 179854
rect 462302 179618 489746 179854
rect 489982 179618 490066 179854
rect 490302 179618 517746 179854
rect 517982 179618 518066 179854
rect 518302 179618 545746 179854
rect 545982 179618 546066 179854
rect 546302 179618 573746 179854
rect 573982 179618 574066 179854
rect 574302 179618 585342 179854
rect 585578 179618 585662 179854
rect 585898 179618 592650 179854
rect -8726 179586 592650 179618
rect -8726 176454 592650 176486
rect -8726 176218 -2934 176454
rect -2698 176218 -2614 176454
rect -2378 176218 38026 176454
rect 38262 176218 38346 176454
rect 38582 176218 66026 176454
rect 66262 176218 66346 176454
rect 66582 176218 94026 176454
rect 94262 176218 94346 176454
rect 94582 176218 122026 176454
rect 122262 176218 122346 176454
rect 122582 176218 150026 176454
rect 150262 176218 150346 176454
rect 150582 176218 178026 176454
rect 178262 176218 178346 176454
rect 178582 176218 206026 176454
rect 206262 176218 206346 176454
rect 206582 176218 234026 176454
rect 234262 176218 234346 176454
rect 234582 176218 262026 176454
rect 262262 176218 262346 176454
rect 262582 176218 290026 176454
rect 290262 176218 290346 176454
rect 290582 176218 318026 176454
rect 318262 176218 318346 176454
rect 318582 176218 346026 176454
rect 346262 176218 346346 176454
rect 346582 176218 374026 176454
rect 374262 176218 374346 176454
rect 374582 176218 402026 176454
rect 402262 176218 402346 176454
rect 402582 176218 430026 176454
rect 430262 176218 430346 176454
rect 430582 176218 458026 176454
rect 458262 176218 458346 176454
rect 458582 176218 486026 176454
rect 486262 176218 486346 176454
rect 486582 176218 514026 176454
rect 514262 176218 514346 176454
rect 514582 176218 542026 176454
rect 542262 176218 542346 176454
rect 542582 176218 570026 176454
rect 570262 176218 570346 176454
rect 570582 176218 586302 176454
rect 586538 176218 586622 176454
rect 586858 176218 592650 176454
rect -8726 176134 592650 176218
rect -8726 175898 -2934 176134
rect -2698 175898 -2614 176134
rect -2378 175898 38026 176134
rect 38262 175898 38346 176134
rect 38582 175898 66026 176134
rect 66262 175898 66346 176134
rect 66582 175898 94026 176134
rect 94262 175898 94346 176134
rect 94582 175898 122026 176134
rect 122262 175898 122346 176134
rect 122582 175898 150026 176134
rect 150262 175898 150346 176134
rect 150582 175898 178026 176134
rect 178262 175898 178346 176134
rect 178582 175898 206026 176134
rect 206262 175898 206346 176134
rect 206582 175898 234026 176134
rect 234262 175898 234346 176134
rect 234582 175898 262026 176134
rect 262262 175898 262346 176134
rect 262582 175898 290026 176134
rect 290262 175898 290346 176134
rect 290582 175898 318026 176134
rect 318262 175898 318346 176134
rect 318582 175898 346026 176134
rect 346262 175898 346346 176134
rect 346582 175898 374026 176134
rect 374262 175898 374346 176134
rect 374582 175898 402026 176134
rect 402262 175898 402346 176134
rect 402582 175898 430026 176134
rect 430262 175898 430346 176134
rect 430582 175898 458026 176134
rect 458262 175898 458346 176134
rect 458582 175898 486026 176134
rect 486262 175898 486346 176134
rect 486582 175898 514026 176134
rect 514262 175898 514346 176134
rect 514582 175898 542026 176134
rect 542262 175898 542346 176134
rect 542582 175898 570026 176134
rect 570262 175898 570346 176134
rect 570582 175898 586302 176134
rect 586538 175898 586622 176134
rect 586858 175898 592650 176134
rect -8726 175866 592650 175898
rect -8726 143174 592650 143206
rect -8726 142938 -1974 143174
rect -1738 142938 -1654 143174
rect -1418 142938 41746 143174
rect 41982 142938 42066 143174
rect 42302 142938 69746 143174
rect 69982 142938 70066 143174
rect 70302 142938 97746 143174
rect 97982 142938 98066 143174
rect 98302 142938 125746 143174
rect 125982 142938 126066 143174
rect 126302 142938 153746 143174
rect 153982 142938 154066 143174
rect 154302 142938 181746 143174
rect 181982 142938 182066 143174
rect 182302 142938 209746 143174
rect 209982 142938 210066 143174
rect 210302 142938 237746 143174
rect 237982 142938 238066 143174
rect 238302 142938 265746 143174
rect 265982 142938 266066 143174
rect 266302 142938 293746 143174
rect 293982 142938 294066 143174
rect 294302 142938 321746 143174
rect 321982 142938 322066 143174
rect 322302 142938 349746 143174
rect 349982 142938 350066 143174
rect 350302 142938 377746 143174
rect 377982 142938 378066 143174
rect 378302 142938 405746 143174
rect 405982 142938 406066 143174
rect 406302 142938 433746 143174
rect 433982 142938 434066 143174
rect 434302 142938 461746 143174
rect 461982 142938 462066 143174
rect 462302 142938 489746 143174
rect 489982 142938 490066 143174
rect 490302 142938 517746 143174
rect 517982 142938 518066 143174
rect 518302 142938 545746 143174
rect 545982 142938 546066 143174
rect 546302 142938 573746 143174
rect 573982 142938 574066 143174
rect 574302 142938 585342 143174
rect 585578 142938 585662 143174
rect 585898 142938 592650 143174
rect -8726 142854 592650 142938
rect -8726 142618 -1974 142854
rect -1738 142618 -1654 142854
rect -1418 142618 41746 142854
rect 41982 142618 42066 142854
rect 42302 142618 69746 142854
rect 69982 142618 70066 142854
rect 70302 142618 97746 142854
rect 97982 142618 98066 142854
rect 98302 142618 125746 142854
rect 125982 142618 126066 142854
rect 126302 142618 153746 142854
rect 153982 142618 154066 142854
rect 154302 142618 181746 142854
rect 181982 142618 182066 142854
rect 182302 142618 209746 142854
rect 209982 142618 210066 142854
rect 210302 142618 237746 142854
rect 237982 142618 238066 142854
rect 238302 142618 265746 142854
rect 265982 142618 266066 142854
rect 266302 142618 293746 142854
rect 293982 142618 294066 142854
rect 294302 142618 321746 142854
rect 321982 142618 322066 142854
rect 322302 142618 349746 142854
rect 349982 142618 350066 142854
rect 350302 142618 377746 142854
rect 377982 142618 378066 142854
rect 378302 142618 405746 142854
rect 405982 142618 406066 142854
rect 406302 142618 433746 142854
rect 433982 142618 434066 142854
rect 434302 142618 461746 142854
rect 461982 142618 462066 142854
rect 462302 142618 489746 142854
rect 489982 142618 490066 142854
rect 490302 142618 517746 142854
rect 517982 142618 518066 142854
rect 518302 142618 545746 142854
rect 545982 142618 546066 142854
rect 546302 142618 573746 142854
rect 573982 142618 574066 142854
rect 574302 142618 585342 142854
rect 585578 142618 585662 142854
rect 585898 142618 592650 142854
rect -8726 142586 592650 142618
rect -8726 139454 592650 139486
rect -8726 139218 -2934 139454
rect -2698 139218 -2614 139454
rect -2378 139218 38026 139454
rect 38262 139218 38346 139454
rect 38582 139218 66026 139454
rect 66262 139218 66346 139454
rect 66582 139218 94026 139454
rect 94262 139218 94346 139454
rect 94582 139218 122026 139454
rect 122262 139218 122346 139454
rect 122582 139218 150026 139454
rect 150262 139218 150346 139454
rect 150582 139218 178026 139454
rect 178262 139218 178346 139454
rect 178582 139218 206026 139454
rect 206262 139218 206346 139454
rect 206582 139218 234026 139454
rect 234262 139218 234346 139454
rect 234582 139218 262026 139454
rect 262262 139218 262346 139454
rect 262582 139218 290026 139454
rect 290262 139218 290346 139454
rect 290582 139218 318026 139454
rect 318262 139218 318346 139454
rect 318582 139218 346026 139454
rect 346262 139218 346346 139454
rect 346582 139218 374026 139454
rect 374262 139218 374346 139454
rect 374582 139218 402026 139454
rect 402262 139218 402346 139454
rect 402582 139218 430026 139454
rect 430262 139218 430346 139454
rect 430582 139218 458026 139454
rect 458262 139218 458346 139454
rect 458582 139218 486026 139454
rect 486262 139218 486346 139454
rect 486582 139218 514026 139454
rect 514262 139218 514346 139454
rect 514582 139218 542026 139454
rect 542262 139218 542346 139454
rect 542582 139218 570026 139454
rect 570262 139218 570346 139454
rect 570582 139218 586302 139454
rect 586538 139218 586622 139454
rect 586858 139218 592650 139454
rect -8726 139134 592650 139218
rect -8726 138898 -2934 139134
rect -2698 138898 -2614 139134
rect -2378 138898 38026 139134
rect 38262 138898 38346 139134
rect 38582 138898 66026 139134
rect 66262 138898 66346 139134
rect 66582 138898 94026 139134
rect 94262 138898 94346 139134
rect 94582 138898 122026 139134
rect 122262 138898 122346 139134
rect 122582 138898 150026 139134
rect 150262 138898 150346 139134
rect 150582 138898 178026 139134
rect 178262 138898 178346 139134
rect 178582 138898 206026 139134
rect 206262 138898 206346 139134
rect 206582 138898 234026 139134
rect 234262 138898 234346 139134
rect 234582 138898 262026 139134
rect 262262 138898 262346 139134
rect 262582 138898 290026 139134
rect 290262 138898 290346 139134
rect 290582 138898 318026 139134
rect 318262 138898 318346 139134
rect 318582 138898 346026 139134
rect 346262 138898 346346 139134
rect 346582 138898 374026 139134
rect 374262 138898 374346 139134
rect 374582 138898 402026 139134
rect 402262 138898 402346 139134
rect 402582 138898 430026 139134
rect 430262 138898 430346 139134
rect 430582 138898 458026 139134
rect 458262 138898 458346 139134
rect 458582 138898 486026 139134
rect 486262 138898 486346 139134
rect 486582 138898 514026 139134
rect 514262 138898 514346 139134
rect 514582 138898 542026 139134
rect 542262 138898 542346 139134
rect 542582 138898 570026 139134
rect 570262 138898 570346 139134
rect 570582 138898 586302 139134
rect 586538 138898 586622 139134
rect 586858 138898 592650 139134
rect -8726 138866 592650 138898
rect -8726 106174 592650 106206
rect -8726 105938 -1974 106174
rect -1738 105938 -1654 106174
rect -1418 105938 41746 106174
rect 41982 105938 42066 106174
rect 42302 105938 69746 106174
rect 69982 105938 70066 106174
rect 70302 105938 97746 106174
rect 97982 105938 98066 106174
rect 98302 105938 125746 106174
rect 125982 105938 126066 106174
rect 126302 105938 153746 106174
rect 153982 105938 154066 106174
rect 154302 105938 181746 106174
rect 181982 105938 182066 106174
rect 182302 105938 209746 106174
rect 209982 105938 210066 106174
rect 210302 105938 237746 106174
rect 237982 105938 238066 106174
rect 238302 105938 265746 106174
rect 265982 105938 266066 106174
rect 266302 105938 293746 106174
rect 293982 105938 294066 106174
rect 294302 105938 321746 106174
rect 321982 105938 322066 106174
rect 322302 105938 349746 106174
rect 349982 105938 350066 106174
rect 350302 105938 377746 106174
rect 377982 105938 378066 106174
rect 378302 105938 405746 106174
rect 405982 105938 406066 106174
rect 406302 105938 433746 106174
rect 433982 105938 434066 106174
rect 434302 105938 461746 106174
rect 461982 105938 462066 106174
rect 462302 105938 489746 106174
rect 489982 105938 490066 106174
rect 490302 105938 517746 106174
rect 517982 105938 518066 106174
rect 518302 105938 545746 106174
rect 545982 105938 546066 106174
rect 546302 105938 573746 106174
rect 573982 105938 574066 106174
rect 574302 105938 585342 106174
rect 585578 105938 585662 106174
rect 585898 105938 592650 106174
rect -8726 105854 592650 105938
rect -8726 105618 -1974 105854
rect -1738 105618 -1654 105854
rect -1418 105618 41746 105854
rect 41982 105618 42066 105854
rect 42302 105618 69746 105854
rect 69982 105618 70066 105854
rect 70302 105618 97746 105854
rect 97982 105618 98066 105854
rect 98302 105618 125746 105854
rect 125982 105618 126066 105854
rect 126302 105618 153746 105854
rect 153982 105618 154066 105854
rect 154302 105618 181746 105854
rect 181982 105618 182066 105854
rect 182302 105618 209746 105854
rect 209982 105618 210066 105854
rect 210302 105618 237746 105854
rect 237982 105618 238066 105854
rect 238302 105618 265746 105854
rect 265982 105618 266066 105854
rect 266302 105618 293746 105854
rect 293982 105618 294066 105854
rect 294302 105618 321746 105854
rect 321982 105618 322066 105854
rect 322302 105618 349746 105854
rect 349982 105618 350066 105854
rect 350302 105618 377746 105854
rect 377982 105618 378066 105854
rect 378302 105618 405746 105854
rect 405982 105618 406066 105854
rect 406302 105618 433746 105854
rect 433982 105618 434066 105854
rect 434302 105618 461746 105854
rect 461982 105618 462066 105854
rect 462302 105618 489746 105854
rect 489982 105618 490066 105854
rect 490302 105618 517746 105854
rect 517982 105618 518066 105854
rect 518302 105618 545746 105854
rect 545982 105618 546066 105854
rect 546302 105618 573746 105854
rect 573982 105618 574066 105854
rect 574302 105618 585342 105854
rect 585578 105618 585662 105854
rect 585898 105618 592650 105854
rect -8726 105586 592650 105618
rect -8726 102454 592650 102486
rect -8726 102218 -2934 102454
rect -2698 102218 -2614 102454
rect -2378 102218 38026 102454
rect 38262 102218 38346 102454
rect 38582 102218 66026 102454
rect 66262 102218 66346 102454
rect 66582 102218 94026 102454
rect 94262 102218 94346 102454
rect 94582 102218 122026 102454
rect 122262 102218 122346 102454
rect 122582 102218 150026 102454
rect 150262 102218 150346 102454
rect 150582 102218 178026 102454
rect 178262 102218 178346 102454
rect 178582 102218 206026 102454
rect 206262 102218 206346 102454
rect 206582 102218 234026 102454
rect 234262 102218 234346 102454
rect 234582 102218 262026 102454
rect 262262 102218 262346 102454
rect 262582 102218 290026 102454
rect 290262 102218 290346 102454
rect 290582 102218 318026 102454
rect 318262 102218 318346 102454
rect 318582 102218 346026 102454
rect 346262 102218 346346 102454
rect 346582 102218 374026 102454
rect 374262 102218 374346 102454
rect 374582 102218 402026 102454
rect 402262 102218 402346 102454
rect 402582 102218 430026 102454
rect 430262 102218 430346 102454
rect 430582 102218 458026 102454
rect 458262 102218 458346 102454
rect 458582 102218 486026 102454
rect 486262 102218 486346 102454
rect 486582 102218 514026 102454
rect 514262 102218 514346 102454
rect 514582 102218 542026 102454
rect 542262 102218 542346 102454
rect 542582 102218 570026 102454
rect 570262 102218 570346 102454
rect 570582 102218 586302 102454
rect 586538 102218 586622 102454
rect 586858 102218 592650 102454
rect -8726 102134 592650 102218
rect -8726 101898 -2934 102134
rect -2698 101898 -2614 102134
rect -2378 101898 38026 102134
rect 38262 101898 38346 102134
rect 38582 101898 66026 102134
rect 66262 101898 66346 102134
rect 66582 101898 94026 102134
rect 94262 101898 94346 102134
rect 94582 101898 122026 102134
rect 122262 101898 122346 102134
rect 122582 101898 150026 102134
rect 150262 101898 150346 102134
rect 150582 101898 178026 102134
rect 178262 101898 178346 102134
rect 178582 101898 206026 102134
rect 206262 101898 206346 102134
rect 206582 101898 234026 102134
rect 234262 101898 234346 102134
rect 234582 101898 262026 102134
rect 262262 101898 262346 102134
rect 262582 101898 290026 102134
rect 290262 101898 290346 102134
rect 290582 101898 318026 102134
rect 318262 101898 318346 102134
rect 318582 101898 346026 102134
rect 346262 101898 346346 102134
rect 346582 101898 374026 102134
rect 374262 101898 374346 102134
rect 374582 101898 402026 102134
rect 402262 101898 402346 102134
rect 402582 101898 430026 102134
rect 430262 101898 430346 102134
rect 430582 101898 458026 102134
rect 458262 101898 458346 102134
rect 458582 101898 486026 102134
rect 486262 101898 486346 102134
rect 486582 101898 514026 102134
rect 514262 101898 514346 102134
rect 514582 101898 542026 102134
rect 542262 101898 542346 102134
rect 542582 101898 570026 102134
rect 570262 101898 570346 102134
rect 570582 101898 586302 102134
rect 586538 101898 586622 102134
rect 586858 101898 592650 102134
rect -8726 101866 592650 101898
rect -8726 69174 592650 69206
rect -8726 68938 -1974 69174
rect -1738 68938 -1654 69174
rect -1418 68938 41746 69174
rect 41982 68938 42066 69174
rect 42302 68938 69746 69174
rect 69982 68938 70066 69174
rect 70302 68938 97746 69174
rect 97982 68938 98066 69174
rect 98302 68938 125746 69174
rect 125982 68938 126066 69174
rect 126302 68938 153746 69174
rect 153982 68938 154066 69174
rect 154302 68938 181746 69174
rect 181982 68938 182066 69174
rect 182302 68938 209746 69174
rect 209982 68938 210066 69174
rect 210302 68938 237746 69174
rect 237982 68938 238066 69174
rect 238302 68938 265746 69174
rect 265982 68938 266066 69174
rect 266302 68938 293746 69174
rect 293982 68938 294066 69174
rect 294302 68938 321746 69174
rect 321982 68938 322066 69174
rect 322302 68938 349746 69174
rect 349982 68938 350066 69174
rect 350302 68938 377746 69174
rect 377982 68938 378066 69174
rect 378302 68938 405746 69174
rect 405982 68938 406066 69174
rect 406302 68938 433746 69174
rect 433982 68938 434066 69174
rect 434302 68938 461746 69174
rect 461982 68938 462066 69174
rect 462302 68938 489746 69174
rect 489982 68938 490066 69174
rect 490302 68938 517746 69174
rect 517982 68938 518066 69174
rect 518302 68938 545746 69174
rect 545982 68938 546066 69174
rect 546302 68938 573746 69174
rect 573982 68938 574066 69174
rect 574302 68938 585342 69174
rect 585578 68938 585662 69174
rect 585898 68938 592650 69174
rect -8726 68854 592650 68938
rect -8726 68618 -1974 68854
rect -1738 68618 -1654 68854
rect -1418 68618 41746 68854
rect 41982 68618 42066 68854
rect 42302 68618 69746 68854
rect 69982 68618 70066 68854
rect 70302 68618 97746 68854
rect 97982 68618 98066 68854
rect 98302 68618 125746 68854
rect 125982 68618 126066 68854
rect 126302 68618 153746 68854
rect 153982 68618 154066 68854
rect 154302 68618 181746 68854
rect 181982 68618 182066 68854
rect 182302 68618 209746 68854
rect 209982 68618 210066 68854
rect 210302 68618 237746 68854
rect 237982 68618 238066 68854
rect 238302 68618 265746 68854
rect 265982 68618 266066 68854
rect 266302 68618 293746 68854
rect 293982 68618 294066 68854
rect 294302 68618 321746 68854
rect 321982 68618 322066 68854
rect 322302 68618 349746 68854
rect 349982 68618 350066 68854
rect 350302 68618 377746 68854
rect 377982 68618 378066 68854
rect 378302 68618 405746 68854
rect 405982 68618 406066 68854
rect 406302 68618 433746 68854
rect 433982 68618 434066 68854
rect 434302 68618 461746 68854
rect 461982 68618 462066 68854
rect 462302 68618 489746 68854
rect 489982 68618 490066 68854
rect 490302 68618 517746 68854
rect 517982 68618 518066 68854
rect 518302 68618 545746 68854
rect 545982 68618 546066 68854
rect 546302 68618 573746 68854
rect 573982 68618 574066 68854
rect 574302 68618 585342 68854
rect 585578 68618 585662 68854
rect 585898 68618 592650 68854
rect -8726 68586 592650 68618
rect -8726 65454 592650 65486
rect -8726 65218 -2934 65454
rect -2698 65218 -2614 65454
rect -2378 65218 38026 65454
rect 38262 65218 38346 65454
rect 38582 65218 66026 65454
rect 66262 65218 66346 65454
rect 66582 65218 94026 65454
rect 94262 65218 94346 65454
rect 94582 65218 122026 65454
rect 122262 65218 122346 65454
rect 122582 65218 150026 65454
rect 150262 65218 150346 65454
rect 150582 65218 178026 65454
rect 178262 65218 178346 65454
rect 178582 65218 206026 65454
rect 206262 65218 206346 65454
rect 206582 65218 234026 65454
rect 234262 65218 234346 65454
rect 234582 65218 262026 65454
rect 262262 65218 262346 65454
rect 262582 65218 290026 65454
rect 290262 65218 290346 65454
rect 290582 65218 318026 65454
rect 318262 65218 318346 65454
rect 318582 65218 346026 65454
rect 346262 65218 346346 65454
rect 346582 65218 374026 65454
rect 374262 65218 374346 65454
rect 374582 65218 402026 65454
rect 402262 65218 402346 65454
rect 402582 65218 430026 65454
rect 430262 65218 430346 65454
rect 430582 65218 458026 65454
rect 458262 65218 458346 65454
rect 458582 65218 486026 65454
rect 486262 65218 486346 65454
rect 486582 65218 514026 65454
rect 514262 65218 514346 65454
rect 514582 65218 542026 65454
rect 542262 65218 542346 65454
rect 542582 65218 570026 65454
rect 570262 65218 570346 65454
rect 570582 65218 586302 65454
rect 586538 65218 586622 65454
rect 586858 65218 592650 65454
rect -8726 65134 592650 65218
rect -8726 64898 -2934 65134
rect -2698 64898 -2614 65134
rect -2378 64898 38026 65134
rect 38262 64898 38346 65134
rect 38582 64898 66026 65134
rect 66262 64898 66346 65134
rect 66582 64898 94026 65134
rect 94262 64898 94346 65134
rect 94582 64898 122026 65134
rect 122262 64898 122346 65134
rect 122582 64898 150026 65134
rect 150262 64898 150346 65134
rect 150582 64898 178026 65134
rect 178262 64898 178346 65134
rect 178582 64898 206026 65134
rect 206262 64898 206346 65134
rect 206582 64898 234026 65134
rect 234262 64898 234346 65134
rect 234582 64898 262026 65134
rect 262262 64898 262346 65134
rect 262582 64898 290026 65134
rect 290262 64898 290346 65134
rect 290582 64898 318026 65134
rect 318262 64898 318346 65134
rect 318582 64898 346026 65134
rect 346262 64898 346346 65134
rect 346582 64898 374026 65134
rect 374262 64898 374346 65134
rect 374582 64898 402026 65134
rect 402262 64898 402346 65134
rect 402582 64898 430026 65134
rect 430262 64898 430346 65134
rect 430582 64898 458026 65134
rect 458262 64898 458346 65134
rect 458582 64898 486026 65134
rect 486262 64898 486346 65134
rect 486582 64898 514026 65134
rect 514262 64898 514346 65134
rect 514582 64898 542026 65134
rect 542262 64898 542346 65134
rect 542582 64898 570026 65134
rect 570262 64898 570346 65134
rect 570582 64898 586302 65134
rect 586538 64898 586622 65134
rect 586858 64898 592650 65134
rect -8726 64866 592650 64898
rect -8726 32174 592650 32206
rect -8726 31938 -1974 32174
rect -1738 31938 -1654 32174
rect -1418 31938 26460 32174
rect 26696 31938 37408 32174
rect 37644 31938 41746 32174
rect 41982 31938 42066 32174
rect 42302 31938 48356 32174
rect 48592 31938 59304 32174
rect 59540 31938 69746 32174
rect 69982 31938 70066 32174
rect 70302 31938 91860 32174
rect 92096 31938 92808 32174
rect 93044 31938 93756 32174
rect 93992 31938 94704 32174
rect 94940 31938 97746 32174
rect 97982 31938 98066 32174
rect 98302 31938 102059 32174
rect 102295 31938 109005 32174
rect 109241 31938 115951 32174
rect 116187 31938 122897 32174
rect 123133 31938 132060 32174
rect 132296 31938 133008 32174
rect 133244 31938 133956 32174
rect 134192 31938 134904 32174
rect 135140 31938 142259 32174
rect 142495 31938 149205 32174
rect 149441 31938 153746 32174
rect 153982 31938 154066 32174
rect 154302 31938 156151 32174
rect 156387 31938 163097 32174
rect 163333 31938 172260 32174
rect 172496 31938 173208 32174
rect 173444 31938 174156 32174
rect 174392 31938 175104 32174
rect 175340 31938 181746 32174
rect 181982 31938 182066 32174
rect 182302 31938 182459 32174
rect 182695 31938 189405 32174
rect 189641 31938 196351 32174
rect 196587 31938 203297 32174
rect 203533 31938 209746 32174
rect 209982 31938 210066 32174
rect 210302 31938 212460 32174
rect 212696 31938 213408 32174
rect 213644 31938 214356 32174
rect 214592 31938 215304 32174
rect 215540 31938 222659 32174
rect 222895 31938 229605 32174
rect 229841 31938 236551 32174
rect 236787 31938 243497 32174
rect 243733 31938 252660 32174
rect 252896 31938 253608 32174
rect 253844 31938 254556 32174
rect 254792 31938 255504 32174
rect 255740 31938 262859 32174
rect 263095 31938 269805 32174
rect 270041 31938 276751 32174
rect 276987 31938 283697 32174
rect 283933 31938 293746 32174
rect 293982 31938 294066 32174
rect 294302 31938 321746 32174
rect 321982 31938 322066 32174
rect 322302 31938 349746 32174
rect 349982 31938 350066 32174
rect 350302 31938 377746 32174
rect 377982 31938 378066 32174
rect 378302 31938 405746 32174
rect 405982 31938 406066 32174
rect 406302 31938 433746 32174
rect 433982 31938 434066 32174
rect 434302 31938 461746 32174
rect 461982 31938 462066 32174
rect 462302 31938 489746 32174
rect 489982 31938 490066 32174
rect 490302 31938 517746 32174
rect 517982 31938 518066 32174
rect 518302 31938 545746 32174
rect 545982 31938 546066 32174
rect 546302 31938 573746 32174
rect 573982 31938 574066 32174
rect 574302 31938 585342 32174
rect 585578 31938 585662 32174
rect 585898 31938 592650 32174
rect -8726 31854 592650 31938
rect -8726 31618 -1974 31854
rect -1738 31618 -1654 31854
rect -1418 31618 26460 31854
rect 26696 31618 37408 31854
rect 37644 31618 41746 31854
rect 41982 31618 42066 31854
rect 42302 31618 48356 31854
rect 48592 31618 59304 31854
rect 59540 31618 69746 31854
rect 69982 31618 70066 31854
rect 70302 31618 91860 31854
rect 92096 31618 92808 31854
rect 93044 31618 93756 31854
rect 93992 31618 94704 31854
rect 94940 31618 97746 31854
rect 97982 31618 98066 31854
rect 98302 31618 102059 31854
rect 102295 31618 109005 31854
rect 109241 31618 115951 31854
rect 116187 31618 122897 31854
rect 123133 31618 132060 31854
rect 132296 31618 133008 31854
rect 133244 31618 133956 31854
rect 134192 31618 134904 31854
rect 135140 31618 142259 31854
rect 142495 31618 149205 31854
rect 149441 31618 153746 31854
rect 153982 31618 154066 31854
rect 154302 31618 156151 31854
rect 156387 31618 163097 31854
rect 163333 31618 172260 31854
rect 172496 31618 173208 31854
rect 173444 31618 174156 31854
rect 174392 31618 175104 31854
rect 175340 31618 181746 31854
rect 181982 31618 182066 31854
rect 182302 31618 182459 31854
rect 182695 31618 189405 31854
rect 189641 31618 196351 31854
rect 196587 31618 203297 31854
rect 203533 31618 209746 31854
rect 209982 31618 210066 31854
rect 210302 31618 212460 31854
rect 212696 31618 213408 31854
rect 213644 31618 214356 31854
rect 214592 31618 215304 31854
rect 215540 31618 222659 31854
rect 222895 31618 229605 31854
rect 229841 31618 236551 31854
rect 236787 31618 243497 31854
rect 243733 31618 252660 31854
rect 252896 31618 253608 31854
rect 253844 31618 254556 31854
rect 254792 31618 255504 31854
rect 255740 31618 262859 31854
rect 263095 31618 269805 31854
rect 270041 31618 276751 31854
rect 276987 31618 283697 31854
rect 283933 31618 293746 31854
rect 293982 31618 294066 31854
rect 294302 31618 321746 31854
rect 321982 31618 322066 31854
rect 322302 31618 349746 31854
rect 349982 31618 350066 31854
rect 350302 31618 377746 31854
rect 377982 31618 378066 31854
rect 378302 31618 405746 31854
rect 405982 31618 406066 31854
rect 406302 31618 433746 31854
rect 433982 31618 434066 31854
rect 434302 31618 461746 31854
rect 461982 31618 462066 31854
rect 462302 31618 489746 31854
rect 489982 31618 490066 31854
rect 490302 31618 517746 31854
rect 517982 31618 518066 31854
rect 518302 31618 545746 31854
rect 545982 31618 546066 31854
rect 546302 31618 573746 31854
rect 573982 31618 574066 31854
rect 574302 31618 585342 31854
rect 585578 31618 585662 31854
rect 585898 31618 592650 31854
rect -8726 31586 592650 31618
rect -8726 28454 592650 28486
rect -8726 28218 -2934 28454
rect -2698 28218 -2614 28454
rect -2378 28218 31934 28454
rect 32170 28218 38026 28454
rect 38262 28218 38346 28454
rect 38582 28218 42882 28454
rect 43118 28218 53830 28454
rect 54066 28218 64778 28454
rect 65014 28218 66026 28454
rect 66262 28218 66346 28454
rect 66582 28218 92334 28454
rect 92570 28218 93282 28454
rect 93518 28218 94230 28454
rect 94466 28218 105532 28454
rect 105768 28218 112478 28454
rect 112714 28218 119424 28454
rect 119660 28218 122026 28454
rect 122262 28218 122346 28454
rect 122582 28218 126370 28454
rect 126606 28218 132534 28454
rect 132770 28218 133482 28454
rect 133718 28218 134430 28454
rect 134666 28218 145732 28454
rect 145968 28218 150026 28454
rect 150262 28218 150346 28454
rect 150582 28218 152678 28454
rect 152914 28218 159624 28454
rect 159860 28218 166570 28454
rect 166806 28218 172734 28454
rect 172970 28218 173682 28454
rect 173918 28218 174630 28454
rect 174866 28218 178026 28454
rect 178262 28218 178346 28454
rect 178582 28218 185932 28454
rect 186168 28218 192878 28454
rect 193114 28218 199824 28454
rect 200060 28218 206026 28454
rect 206262 28218 206346 28454
rect 206582 28218 206770 28454
rect 207006 28218 212934 28454
rect 213170 28218 213882 28454
rect 214118 28218 214830 28454
rect 215066 28218 226132 28454
rect 226368 28218 233078 28454
rect 233314 28218 240024 28454
rect 240260 28218 246970 28454
rect 247206 28218 253134 28454
rect 253370 28218 254082 28454
rect 254318 28218 255030 28454
rect 255266 28218 266332 28454
rect 266568 28218 273278 28454
rect 273514 28218 280224 28454
rect 280460 28218 287170 28454
rect 287406 28218 290026 28454
rect 290262 28218 290346 28454
rect 290582 28218 318026 28454
rect 318262 28218 318346 28454
rect 318582 28218 346026 28454
rect 346262 28218 346346 28454
rect 346582 28218 374026 28454
rect 374262 28218 374346 28454
rect 374582 28218 402026 28454
rect 402262 28218 402346 28454
rect 402582 28218 430026 28454
rect 430262 28218 430346 28454
rect 430582 28218 458026 28454
rect 458262 28218 458346 28454
rect 458582 28218 486026 28454
rect 486262 28218 486346 28454
rect 486582 28218 514026 28454
rect 514262 28218 514346 28454
rect 514582 28218 542026 28454
rect 542262 28218 542346 28454
rect 542582 28218 570026 28454
rect 570262 28218 570346 28454
rect 570582 28218 586302 28454
rect 586538 28218 586622 28454
rect 586858 28218 592650 28454
rect -8726 28134 592650 28218
rect -8726 27898 -2934 28134
rect -2698 27898 -2614 28134
rect -2378 27898 31934 28134
rect 32170 27898 38026 28134
rect 38262 27898 38346 28134
rect 38582 27898 42882 28134
rect 43118 27898 53830 28134
rect 54066 27898 64778 28134
rect 65014 27898 66026 28134
rect 66262 27898 66346 28134
rect 66582 27898 92334 28134
rect 92570 27898 93282 28134
rect 93518 27898 94230 28134
rect 94466 27898 105532 28134
rect 105768 27898 112478 28134
rect 112714 27898 119424 28134
rect 119660 27898 122026 28134
rect 122262 27898 122346 28134
rect 122582 27898 126370 28134
rect 126606 27898 132534 28134
rect 132770 27898 133482 28134
rect 133718 27898 134430 28134
rect 134666 27898 145732 28134
rect 145968 27898 150026 28134
rect 150262 27898 150346 28134
rect 150582 27898 152678 28134
rect 152914 27898 159624 28134
rect 159860 27898 166570 28134
rect 166806 27898 172734 28134
rect 172970 27898 173682 28134
rect 173918 27898 174630 28134
rect 174866 27898 178026 28134
rect 178262 27898 178346 28134
rect 178582 27898 185932 28134
rect 186168 27898 192878 28134
rect 193114 27898 199824 28134
rect 200060 27898 206026 28134
rect 206262 27898 206346 28134
rect 206582 27898 206770 28134
rect 207006 27898 212934 28134
rect 213170 27898 213882 28134
rect 214118 27898 214830 28134
rect 215066 27898 226132 28134
rect 226368 27898 233078 28134
rect 233314 27898 240024 28134
rect 240260 27898 246970 28134
rect 247206 27898 253134 28134
rect 253370 27898 254082 28134
rect 254318 27898 255030 28134
rect 255266 27898 266332 28134
rect 266568 27898 273278 28134
rect 273514 27898 280224 28134
rect 280460 27898 287170 28134
rect 287406 27898 290026 28134
rect 290262 27898 290346 28134
rect 290582 27898 318026 28134
rect 318262 27898 318346 28134
rect 318582 27898 346026 28134
rect 346262 27898 346346 28134
rect 346582 27898 374026 28134
rect 374262 27898 374346 28134
rect 374582 27898 402026 28134
rect 402262 27898 402346 28134
rect 402582 27898 430026 28134
rect 430262 27898 430346 28134
rect 430582 27898 458026 28134
rect 458262 27898 458346 28134
rect 458582 27898 486026 28134
rect 486262 27898 486346 28134
rect 486582 27898 514026 28134
rect 514262 27898 514346 28134
rect 514582 27898 542026 28134
rect 542262 27898 542346 28134
rect 542582 27898 570026 28134
rect 570262 27898 570346 28134
rect 570582 27898 586302 28134
rect 586538 27898 586622 28134
rect 586858 27898 592650 28134
rect -8726 27866 592650 27898
rect -2006 -346 585930 -314
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 41746 -346
rect 41982 -582 42066 -346
rect 42302 -582 69746 -346
rect 69982 -582 70066 -346
rect 70302 -582 97746 -346
rect 97982 -582 98066 -346
rect 98302 -582 153746 -346
rect 153982 -582 154066 -346
rect 154302 -582 181746 -346
rect 181982 -582 182066 -346
rect 182302 -582 209746 -346
rect 209982 -582 210066 -346
rect 210302 -582 293746 -346
rect 293982 -582 294066 -346
rect 294302 -582 321746 -346
rect 321982 -582 322066 -346
rect 322302 -582 349746 -346
rect 349982 -582 350066 -346
rect 350302 -582 377746 -346
rect 377982 -582 378066 -346
rect 378302 -582 405746 -346
rect 405982 -582 406066 -346
rect 406302 -582 433746 -346
rect 433982 -582 434066 -346
rect 434302 -582 461746 -346
rect 461982 -582 462066 -346
rect 462302 -582 489746 -346
rect 489982 -582 490066 -346
rect 490302 -582 517746 -346
rect 517982 -582 518066 -346
rect 518302 -582 545746 -346
rect 545982 -582 546066 -346
rect 546302 -582 573746 -346
rect 573982 -582 574066 -346
rect 574302 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect -2006 -666 585930 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 41746 -666
rect 41982 -902 42066 -666
rect 42302 -902 69746 -666
rect 69982 -902 70066 -666
rect 70302 -902 97746 -666
rect 97982 -902 98066 -666
rect 98302 -902 153746 -666
rect 153982 -902 154066 -666
rect 154302 -902 181746 -666
rect 181982 -902 182066 -666
rect 182302 -902 209746 -666
rect 209982 -902 210066 -666
rect 210302 -902 293746 -666
rect 293982 -902 294066 -666
rect 294302 -902 321746 -666
rect 321982 -902 322066 -666
rect 322302 -902 349746 -666
rect 349982 -902 350066 -666
rect 350302 -902 377746 -666
rect 377982 -902 378066 -666
rect 378302 -902 405746 -666
rect 405982 -902 406066 -666
rect 406302 -902 433746 -666
rect 433982 -902 434066 -666
rect 434302 -902 461746 -666
rect 461982 -902 462066 -666
rect 462302 -902 489746 -666
rect 489982 -902 490066 -666
rect 490302 -902 517746 -666
rect 517982 -902 518066 -666
rect 518302 -902 545746 -666
rect 545982 -902 546066 -666
rect 546302 -902 573746 -666
rect 573982 -902 574066 -666
rect 574302 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect -2006 -934 585930 -902
rect -2966 -1306 586890 -1274
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 38026 -1306
rect 38262 -1542 38346 -1306
rect 38582 -1542 66026 -1306
rect 66262 -1542 66346 -1306
rect 66582 -1542 122026 -1306
rect 122262 -1542 122346 -1306
rect 122582 -1542 150026 -1306
rect 150262 -1542 150346 -1306
rect 150582 -1542 178026 -1306
rect 178262 -1542 178346 -1306
rect 178582 -1542 206026 -1306
rect 206262 -1542 206346 -1306
rect 206582 -1542 290026 -1306
rect 290262 -1542 290346 -1306
rect 290582 -1542 318026 -1306
rect 318262 -1542 318346 -1306
rect 318582 -1542 346026 -1306
rect 346262 -1542 346346 -1306
rect 346582 -1542 374026 -1306
rect 374262 -1542 374346 -1306
rect 374582 -1542 402026 -1306
rect 402262 -1542 402346 -1306
rect 402582 -1542 430026 -1306
rect 430262 -1542 430346 -1306
rect 430582 -1542 458026 -1306
rect 458262 -1542 458346 -1306
rect 458582 -1542 486026 -1306
rect 486262 -1542 486346 -1306
rect 486582 -1542 514026 -1306
rect 514262 -1542 514346 -1306
rect 514582 -1542 542026 -1306
rect 542262 -1542 542346 -1306
rect 542582 -1542 570026 -1306
rect 570262 -1542 570346 -1306
rect 570582 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect -2966 -1626 586890 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 38026 -1626
rect 38262 -1862 38346 -1626
rect 38582 -1862 66026 -1626
rect 66262 -1862 66346 -1626
rect 66582 -1862 122026 -1626
rect 122262 -1862 122346 -1626
rect 122582 -1862 150026 -1626
rect 150262 -1862 150346 -1626
rect 150582 -1862 178026 -1626
rect 178262 -1862 178346 -1626
rect 178582 -1862 206026 -1626
rect 206262 -1862 206346 -1626
rect 206582 -1862 290026 -1626
rect 290262 -1862 290346 -1626
rect 290582 -1862 318026 -1626
rect 318262 -1862 318346 -1626
rect 318582 -1862 346026 -1626
rect 346262 -1862 346346 -1626
rect 346582 -1862 374026 -1626
rect 374262 -1862 374346 -1626
rect 374582 -1862 402026 -1626
rect 402262 -1862 402346 -1626
rect 402582 -1862 430026 -1626
rect 430262 -1862 430346 -1626
rect 430582 -1862 458026 -1626
rect 458262 -1862 458346 -1626
rect 458582 -1862 486026 -1626
rect 486262 -1862 486346 -1626
rect 486582 -1862 514026 -1626
rect 514262 -1862 514346 -1626
rect 514582 -1862 542026 -1626
rect 542262 -1862 542346 -1626
rect 542582 -1862 570026 -1626
rect 570262 -1862 570346 -1626
rect 570582 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect -2966 -1894 586890 -1862
rect -3926 -2266 587850 -2234
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect -3926 -2586 587850 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect -3926 -2854 587850 -2822
rect -4886 -3226 588810 -3194
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect -4886 -3546 588810 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect -4886 -3814 588810 -3782
rect -5846 -4186 589770 -4154
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect -5846 -4506 589770 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect -5846 -4774 589770 -4742
rect -6806 -5146 590730 -5114
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect -6806 -5466 590730 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect -6806 -5734 590730 -5702
rect -7766 -6106 591690 -6074
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect -7766 -6426 591690 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect -7766 -6694 591690 -6662
rect -8726 -7066 592650 -7034
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect -8726 -7386 592650 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect -8726 -7654 592650 -7622
use meiniki_pi  meiniki_pi_003
timestamp 0
transform 1 0 218200 0 1 19000
box 0 31 29979 33425
use scan_controller  scan_controller
timestamp 0
transform 1 0 20000 0 1 20000
box -10 0 46000 20000
use scanchain  scanchain_000
timestamp 0
transform 1 0 90400 0 1 19000
box 0 688 6000 23248
use scanchain  scanchain_001
timestamp 0
transform 1 0 130600 0 1 19000
box 0 688 6000 23248
use scanchain  scanchain_002
timestamp 0
transform 1 0 170800 0 1 19000
box 0 688 6000 23248
use scanchain  scanchain_003
timestamp 0
transform 1 0 211000 0 1 19000
box 0 688 6000 23248
use scanchain  scanchain_004
timestamp 0
transform 1 0 251200 0 1 19000
box 0 688 6000 23248
use user_module_357464855584307201  user_module_357464855584307201_000
timestamp 0
transform 1 0 97600 0 1 19000
box 0 1040 29048 32688
use user_module_357752736742764545  user_module_357752736742764545_002
timestamp 0
transform 1 0 178000 0 1 19000
box 0 1040 29048 32688
use weverest_top  weverest_top_001
timestamp 0
transform 1 0 137800 0 1 19000
box 0 614 29048 32688
use wormy_top  wormy_top_004
timestamp 0
transform 1 0 258400 0 1 19000
box 0 818 29048 32688
<< labels >>
flabel metal3 s 583520 285276 584960 285516 0 FreeSans 960 0 0 0 analog_io[0]
port 0 nsew signal bidirectional
flabel metal2 s 446098 703520 446210 704960 0 FreeSans 448 90 0 0 analog_io[10]
port 1 nsew signal bidirectional
flabel metal2 s 381146 703520 381258 704960 0 FreeSans 448 90 0 0 analog_io[11]
port 2 nsew signal bidirectional
flabel metal2 s 316286 703520 316398 704960 0 FreeSans 448 90 0 0 analog_io[12]
port 3 nsew signal bidirectional
flabel metal2 s 251426 703520 251538 704960 0 FreeSans 448 90 0 0 analog_io[13]
port 4 nsew signal bidirectional
flabel metal2 s 186474 703520 186586 704960 0 FreeSans 448 90 0 0 analog_io[14]
port 5 nsew signal bidirectional
flabel metal2 s 121614 703520 121726 704960 0 FreeSans 448 90 0 0 analog_io[15]
port 6 nsew signal bidirectional
flabel metal2 s 56754 703520 56866 704960 0 FreeSans 448 90 0 0 analog_io[16]
port 7 nsew signal bidirectional
flabel metal3 s -960 697220 480 697460 0 FreeSans 960 0 0 0 analog_io[17]
port 8 nsew signal bidirectional
flabel metal3 s -960 644996 480 645236 0 FreeSans 960 0 0 0 analog_io[18]
port 9 nsew signal bidirectional
flabel metal3 s -960 592908 480 593148 0 FreeSans 960 0 0 0 analog_io[19]
port 10 nsew signal bidirectional
flabel metal3 s 583520 338452 584960 338692 0 FreeSans 960 0 0 0 analog_io[1]
port 11 nsew signal bidirectional
flabel metal3 s -960 540684 480 540924 0 FreeSans 960 0 0 0 analog_io[20]
port 12 nsew signal bidirectional
flabel metal3 s -960 488596 480 488836 0 FreeSans 960 0 0 0 analog_io[21]
port 13 nsew signal bidirectional
flabel metal3 s -960 436508 480 436748 0 FreeSans 960 0 0 0 analog_io[22]
port 14 nsew signal bidirectional
flabel metal3 s -960 384284 480 384524 0 FreeSans 960 0 0 0 analog_io[23]
port 15 nsew signal bidirectional
flabel metal3 s -960 332196 480 332436 0 FreeSans 960 0 0 0 analog_io[24]
port 16 nsew signal bidirectional
flabel metal3 s -960 279972 480 280212 0 FreeSans 960 0 0 0 analog_io[25]
port 17 nsew signal bidirectional
flabel metal3 s -960 227884 480 228124 0 FreeSans 960 0 0 0 analog_io[26]
port 18 nsew signal bidirectional
flabel metal3 s -960 175796 480 176036 0 FreeSans 960 0 0 0 analog_io[27]
port 19 nsew signal bidirectional
flabel metal3 s -960 123572 480 123812 0 FreeSans 960 0 0 0 analog_io[28]
port 20 nsew signal bidirectional
flabel metal3 s 583520 391628 584960 391868 0 FreeSans 960 0 0 0 analog_io[2]
port 21 nsew signal bidirectional
flabel metal3 s 583520 444668 584960 444908 0 FreeSans 960 0 0 0 analog_io[3]
port 22 nsew signal bidirectional
flabel metal3 s 583520 497844 584960 498084 0 FreeSans 960 0 0 0 analog_io[4]
port 23 nsew signal bidirectional
flabel metal3 s 583520 551020 584960 551260 0 FreeSans 960 0 0 0 analog_io[5]
port 24 nsew signal bidirectional
flabel metal3 s 583520 604060 584960 604300 0 FreeSans 960 0 0 0 analog_io[6]
port 25 nsew signal bidirectional
flabel metal3 s 583520 657236 584960 657476 0 FreeSans 960 0 0 0 analog_io[7]
port 26 nsew signal bidirectional
flabel metal2 s 575818 703520 575930 704960 0 FreeSans 448 90 0 0 analog_io[8]
port 27 nsew signal bidirectional
flabel metal2 s 510958 703520 511070 704960 0 FreeSans 448 90 0 0 analog_io[9]
port 28 nsew signal bidirectional
flabel metal3 s 583520 6476 584960 6716 0 FreeSans 960 0 0 0 io_in[0]
port 29 nsew signal input
flabel metal3 s 583520 457996 584960 458236 0 FreeSans 960 0 0 0 io_in[10]
port 30 nsew signal input
flabel metal3 s 583520 511172 584960 511412 0 FreeSans 960 0 0 0 io_in[11]
port 31 nsew signal input
flabel metal3 s 583520 564212 584960 564452 0 FreeSans 960 0 0 0 io_in[12]
port 32 nsew signal input
flabel metal3 s 583520 617388 584960 617628 0 FreeSans 960 0 0 0 io_in[13]
port 33 nsew signal input
flabel metal3 s 583520 670564 584960 670804 0 FreeSans 960 0 0 0 io_in[14]
port 34 nsew signal input
flabel metal2 s 559626 703520 559738 704960 0 FreeSans 448 90 0 0 io_in[15]
port 35 nsew signal input
flabel metal2 s 494766 703520 494878 704960 0 FreeSans 448 90 0 0 io_in[16]
port 36 nsew signal input
flabel metal2 s 429814 703520 429926 704960 0 FreeSans 448 90 0 0 io_in[17]
port 37 nsew signal input
flabel metal2 s 364954 703520 365066 704960 0 FreeSans 448 90 0 0 io_in[18]
port 38 nsew signal input
flabel metal2 s 300094 703520 300206 704960 0 FreeSans 448 90 0 0 io_in[19]
port 39 nsew signal input
flabel metal3 s 583520 46188 584960 46428 0 FreeSans 960 0 0 0 io_in[1]
port 40 nsew signal input
flabel metal2 s 235142 703520 235254 704960 0 FreeSans 448 90 0 0 io_in[20]
port 41 nsew signal input
flabel metal2 s 170282 703520 170394 704960 0 FreeSans 448 90 0 0 io_in[21]
port 42 nsew signal input
flabel metal2 s 105422 703520 105534 704960 0 FreeSans 448 90 0 0 io_in[22]
port 43 nsew signal input
flabel metal2 s 40470 703520 40582 704960 0 FreeSans 448 90 0 0 io_in[23]
port 44 nsew signal input
flabel metal3 s -960 684164 480 684404 0 FreeSans 960 0 0 0 io_in[24]
port 45 nsew signal input
flabel metal3 s -960 631940 480 632180 0 FreeSans 960 0 0 0 io_in[25]
port 46 nsew signal input
flabel metal3 s -960 579852 480 580092 0 FreeSans 960 0 0 0 io_in[26]
port 47 nsew signal input
flabel metal3 s -960 527764 480 528004 0 FreeSans 960 0 0 0 io_in[27]
port 48 nsew signal input
flabel metal3 s -960 475540 480 475780 0 FreeSans 960 0 0 0 io_in[28]
port 49 nsew signal input
flabel metal3 s -960 423452 480 423692 0 FreeSans 960 0 0 0 io_in[29]
port 50 nsew signal input
flabel metal3 s 583520 86036 584960 86276 0 FreeSans 960 0 0 0 io_in[2]
port 51 nsew signal input
flabel metal3 s -960 371228 480 371468 0 FreeSans 960 0 0 0 io_in[30]
port 52 nsew signal input
flabel metal3 s -960 319140 480 319380 0 FreeSans 960 0 0 0 io_in[31]
port 53 nsew signal input
flabel metal3 s -960 267052 480 267292 0 FreeSans 960 0 0 0 io_in[32]
port 54 nsew signal input
flabel metal3 s -960 214828 480 215068 0 FreeSans 960 0 0 0 io_in[33]
port 55 nsew signal input
flabel metal3 s -960 162740 480 162980 0 FreeSans 960 0 0 0 io_in[34]
port 56 nsew signal input
flabel metal3 s -960 110516 480 110756 0 FreeSans 960 0 0 0 io_in[35]
port 57 nsew signal input
flabel metal3 s -960 71484 480 71724 0 FreeSans 960 0 0 0 io_in[36]
port 58 nsew signal input
flabel metal3 s -960 32316 480 32556 0 FreeSans 960 0 0 0 io_in[37]
port 59 nsew signal input
flabel metal3 s 583520 125884 584960 126124 0 FreeSans 960 0 0 0 io_in[3]
port 60 nsew signal input
flabel metal3 s 583520 165732 584960 165972 0 FreeSans 960 0 0 0 io_in[4]
port 61 nsew signal input
flabel metal3 s 583520 205580 584960 205820 0 FreeSans 960 0 0 0 io_in[5]
port 62 nsew signal input
flabel metal3 s 583520 245428 584960 245668 0 FreeSans 960 0 0 0 io_in[6]
port 63 nsew signal input
flabel metal3 s 583520 298604 584960 298844 0 FreeSans 960 0 0 0 io_in[7]
port 64 nsew signal input
flabel metal3 s 583520 351780 584960 352020 0 FreeSans 960 0 0 0 io_in[8]
port 65 nsew signal input
flabel metal3 s 583520 404820 584960 405060 0 FreeSans 960 0 0 0 io_in[9]
port 66 nsew signal input
flabel metal3 s 583520 32996 584960 33236 0 FreeSans 960 0 0 0 io_oeb[0]
port 67 nsew signal tristate
flabel metal3 s 583520 484516 584960 484756 0 FreeSans 960 0 0 0 io_oeb[10]
port 68 nsew signal tristate
flabel metal3 s 583520 537692 584960 537932 0 FreeSans 960 0 0 0 io_oeb[11]
port 69 nsew signal tristate
flabel metal3 s 583520 590868 584960 591108 0 FreeSans 960 0 0 0 io_oeb[12]
port 70 nsew signal tristate
flabel metal3 s 583520 643908 584960 644148 0 FreeSans 960 0 0 0 io_oeb[13]
port 71 nsew signal tristate
flabel metal3 s 583520 697084 584960 697324 0 FreeSans 960 0 0 0 io_oeb[14]
port 72 nsew signal tristate
flabel metal2 s 527150 703520 527262 704960 0 FreeSans 448 90 0 0 io_oeb[15]
port 73 nsew signal tristate
flabel metal2 s 462290 703520 462402 704960 0 FreeSans 448 90 0 0 io_oeb[16]
port 74 nsew signal tristate
flabel metal2 s 397430 703520 397542 704960 0 FreeSans 448 90 0 0 io_oeb[17]
port 75 nsew signal tristate
flabel metal2 s 332478 703520 332590 704960 0 FreeSans 448 90 0 0 io_oeb[18]
port 76 nsew signal tristate
flabel metal2 s 267618 703520 267730 704960 0 FreeSans 448 90 0 0 io_oeb[19]
port 77 nsew signal tristate
flabel metal3 s 583520 72844 584960 73084 0 FreeSans 960 0 0 0 io_oeb[1]
port 78 nsew signal tristate
flabel metal2 s 202758 703520 202870 704960 0 FreeSans 448 90 0 0 io_oeb[20]
port 79 nsew signal tristate
flabel metal2 s 137806 703520 137918 704960 0 FreeSans 448 90 0 0 io_oeb[21]
port 80 nsew signal tristate
flabel metal2 s 72946 703520 73058 704960 0 FreeSans 448 90 0 0 io_oeb[22]
port 81 nsew signal tristate
flabel metal2 s 8086 703520 8198 704960 0 FreeSans 448 90 0 0 io_oeb[23]
port 82 nsew signal tristate
flabel metal3 s -960 658052 480 658292 0 FreeSans 960 0 0 0 io_oeb[24]
port 83 nsew signal tristate
flabel metal3 s -960 605964 480 606204 0 FreeSans 960 0 0 0 io_oeb[25]
port 84 nsew signal tristate
flabel metal3 s -960 553740 480 553980 0 FreeSans 960 0 0 0 io_oeb[26]
port 85 nsew signal tristate
flabel metal3 s -960 501652 480 501892 0 FreeSans 960 0 0 0 io_oeb[27]
port 86 nsew signal tristate
flabel metal3 s -960 449428 480 449668 0 FreeSans 960 0 0 0 io_oeb[28]
port 87 nsew signal tristate
flabel metal3 s -960 397340 480 397580 0 FreeSans 960 0 0 0 io_oeb[29]
port 88 nsew signal tristate
flabel metal3 s 583520 112692 584960 112932 0 FreeSans 960 0 0 0 io_oeb[2]
port 89 nsew signal tristate
flabel metal3 s -960 345252 480 345492 0 FreeSans 960 0 0 0 io_oeb[30]
port 90 nsew signal tristate
flabel metal3 s -960 293028 480 293268 0 FreeSans 960 0 0 0 io_oeb[31]
port 91 nsew signal tristate
flabel metal3 s -960 240940 480 241180 0 FreeSans 960 0 0 0 io_oeb[32]
port 92 nsew signal tristate
flabel metal3 s -960 188716 480 188956 0 FreeSans 960 0 0 0 io_oeb[33]
port 93 nsew signal tristate
flabel metal3 s -960 136628 480 136868 0 FreeSans 960 0 0 0 io_oeb[34]
port 94 nsew signal tristate
flabel metal3 s -960 84540 480 84780 0 FreeSans 960 0 0 0 io_oeb[35]
port 95 nsew signal tristate
flabel metal3 s -960 45372 480 45612 0 FreeSans 960 0 0 0 io_oeb[36]
port 96 nsew signal tristate
flabel metal3 s -960 6340 480 6580 0 FreeSans 960 0 0 0 io_oeb[37]
port 97 nsew signal tristate
flabel metal3 s 583520 152540 584960 152780 0 FreeSans 960 0 0 0 io_oeb[3]
port 98 nsew signal tristate
flabel metal3 s 583520 192388 584960 192628 0 FreeSans 960 0 0 0 io_oeb[4]
port 99 nsew signal tristate
flabel metal3 s 583520 232236 584960 232476 0 FreeSans 960 0 0 0 io_oeb[5]
port 100 nsew signal tristate
flabel metal3 s 583520 272084 584960 272324 0 FreeSans 960 0 0 0 io_oeb[6]
port 101 nsew signal tristate
flabel metal3 s 583520 325124 584960 325364 0 FreeSans 960 0 0 0 io_oeb[7]
port 102 nsew signal tristate
flabel metal3 s 583520 378300 584960 378540 0 FreeSans 960 0 0 0 io_oeb[8]
port 103 nsew signal tristate
flabel metal3 s 583520 431476 584960 431716 0 FreeSans 960 0 0 0 io_oeb[9]
port 104 nsew signal tristate
flabel metal3 s 583520 19668 584960 19908 0 FreeSans 960 0 0 0 io_out[0]
port 105 nsew signal tristate
flabel metal3 s 583520 471324 584960 471564 0 FreeSans 960 0 0 0 io_out[10]
port 106 nsew signal tristate
flabel metal3 s 583520 524364 584960 524604 0 FreeSans 960 0 0 0 io_out[11]
port 107 nsew signal tristate
flabel metal3 s 583520 577540 584960 577780 0 FreeSans 960 0 0 0 io_out[12]
port 108 nsew signal tristate
flabel metal3 s 583520 630716 584960 630956 0 FreeSans 960 0 0 0 io_out[13]
port 109 nsew signal tristate
flabel metal3 s 583520 683756 584960 683996 0 FreeSans 960 0 0 0 io_out[14]
port 110 nsew signal tristate
flabel metal2 s 543434 703520 543546 704960 0 FreeSans 448 90 0 0 io_out[15]
port 111 nsew signal tristate
flabel metal2 s 478482 703520 478594 704960 0 FreeSans 448 90 0 0 io_out[16]
port 112 nsew signal tristate
flabel metal2 s 413622 703520 413734 704960 0 FreeSans 448 90 0 0 io_out[17]
port 113 nsew signal tristate
flabel metal2 s 348762 703520 348874 704960 0 FreeSans 448 90 0 0 io_out[18]
port 114 nsew signal tristate
flabel metal2 s 283810 703520 283922 704960 0 FreeSans 448 90 0 0 io_out[19]
port 115 nsew signal tristate
flabel metal3 s 583520 59516 584960 59756 0 FreeSans 960 0 0 0 io_out[1]
port 116 nsew signal tristate
flabel metal2 s 218950 703520 219062 704960 0 FreeSans 448 90 0 0 io_out[20]
port 117 nsew signal tristate
flabel metal2 s 154090 703520 154202 704960 0 FreeSans 448 90 0 0 io_out[21]
port 118 nsew signal tristate
flabel metal2 s 89138 703520 89250 704960 0 FreeSans 448 90 0 0 io_out[22]
port 119 nsew signal tristate
flabel metal2 s 24278 703520 24390 704960 0 FreeSans 448 90 0 0 io_out[23]
port 120 nsew signal tristate
flabel metal3 s -960 671108 480 671348 0 FreeSans 960 0 0 0 io_out[24]
port 121 nsew signal tristate
flabel metal3 s -960 619020 480 619260 0 FreeSans 960 0 0 0 io_out[25]
port 122 nsew signal tristate
flabel metal3 s -960 566796 480 567036 0 FreeSans 960 0 0 0 io_out[26]
port 123 nsew signal tristate
flabel metal3 s -960 514708 480 514948 0 FreeSans 960 0 0 0 io_out[27]
port 124 nsew signal tristate
flabel metal3 s -960 462484 480 462724 0 FreeSans 960 0 0 0 io_out[28]
port 125 nsew signal tristate
flabel metal3 s -960 410396 480 410636 0 FreeSans 960 0 0 0 io_out[29]
port 126 nsew signal tristate
flabel metal3 s 583520 99364 584960 99604 0 FreeSans 960 0 0 0 io_out[2]
port 127 nsew signal tristate
flabel metal3 s -960 358308 480 358548 0 FreeSans 960 0 0 0 io_out[30]
port 128 nsew signal tristate
flabel metal3 s -960 306084 480 306324 0 FreeSans 960 0 0 0 io_out[31]
port 129 nsew signal tristate
flabel metal3 s -960 253996 480 254236 0 FreeSans 960 0 0 0 io_out[32]
port 130 nsew signal tristate
flabel metal3 s -960 201772 480 202012 0 FreeSans 960 0 0 0 io_out[33]
port 131 nsew signal tristate
flabel metal3 s -960 149684 480 149924 0 FreeSans 960 0 0 0 io_out[34]
port 132 nsew signal tristate
flabel metal3 s -960 97460 480 97700 0 FreeSans 960 0 0 0 io_out[35]
port 133 nsew signal tristate
flabel metal3 s -960 58428 480 58668 0 FreeSans 960 0 0 0 io_out[36]
port 134 nsew signal tristate
flabel metal3 s -960 19260 480 19500 0 FreeSans 960 0 0 0 io_out[37]
port 135 nsew signal tristate
flabel metal3 s 583520 139212 584960 139452 0 FreeSans 960 0 0 0 io_out[3]
port 136 nsew signal tristate
flabel metal3 s 583520 179060 584960 179300 0 FreeSans 960 0 0 0 io_out[4]
port 137 nsew signal tristate
flabel metal3 s 583520 218908 584960 219148 0 FreeSans 960 0 0 0 io_out[5]
port 138 nsew signal tristate
flabel metal3 s 583520 258756 584960 258996 0 FreeSans 960 0 0 0 io_out[6]
port 139 nsew signal tristate
flabel metal3 s 583520 311932 584960 312172 0 FreeSans 960 0 0 0 io_out[7]
port 140 nsew signal tristate
flabel metal3 s 583520 364972 584960 365212 0 FreeSans 960 0 0 0 io_out[8]
port 141 nsew signal tristate
flabel metal3 s 583520 418148 584960 418388 0 FreeSans 960 0 0 0 io_out[9]
port 142 nsew signal tristate
flabel metal2 s 125846 -960 125958 480 0 FreeSans 448 90 0 0 la_data_in[0]
port 143 nsew signal input
flabel metal2 s 480506 -960 480618 480 0 FreeSans 448 90 0 0 la_data_in[100]
port 144 nsew signal input
flabel metal2 s 484002 -960 484114 480 0 FreeSans 448 90 0 0 la_data_in[101]
port 145 nsew signal input
flabel metal2 s 487590 -960 487702 480 0 FreeSans 448 90 0 0 la_data_in[102]
port 146 nsew signal input
flabel metal2 s 491086 -960 491198 480 0 FreeSans 448 90 0 0 la_data_in[103]
port 147 nsew signal input
flabel metal2 s 494674 -960 494786 480 0 FreeSans 448 90 0 0 la_data_in[104]
port 148 nsew signal input
flabel metal2 s 498170 -960 498282 480 0 FreeSans 448 90 0 0 la_data_in[105]
port 149 nsew signal input
flabel metal2 s 501758 -960 501870 480 0 FreeSans 448 90 0 0 la_data_in[106]
port 150 nsew signal input
flabel metal2 s 505346 -960 505458 480 0 FreeSans 448 90 0 0 la_data_in[107]
port 151 nsew signal input
flabel metal2 s 508842 -960 508954 480 0 FreeSans 448 90 0 0 la_data_in[108]
port 152 nsew signal input
flabel metal2 s 512430 -960 512542 480 0 FreeSans 448 90 0 0 la_data_in[109]
port 153 nsew signal input
flabel metal2 s 161266 -960 161378 480 0 FreeSans 448 90 0 0 la_data_in[10]
port 154 nsew signal input
flabel metal2 s 515926 -960 516038 480 0 FreeSans 448 90 0 0 la_data_in[110]
port 155 nsew signal input
flabel metal2 s 519514 -960 519626 480 0 FreeSans 448 90 0 0 la_data_in[111]
port 156 nsew signal input
flabel metal2 s 523010 -960 523122 480 0 FreeSans 448 90 0 0 la_data_in[112]
port 157 nsew signal input
flabel metal2 s 526598 -960 526710 480 0 FreeSans 448 90 0 0 la_data_in[113]
port 158 nsew signal input
flabel metal2 s 530094 -960 530206 480 0 FreeSans 448 90 0 0 la_data_in[114]
port 159 nsew signal input
flabel metal2 s 533682 -960 533794 480 0 FreeSans 448 90 0 0 la_data_in[115]
port 160 nsew signal input
flabel metal2 s 537178 -960 537290 480 0 FreeSans 448 90 0 0 la_data_in[116]
port 161 nsew signal input
flabel metal2 s 540766 -960 540878 480 0 FreeSans 448 90 0 0 la_data_in[117]
port 162 nsew signal input
flabel metal2 s 544354 -960 544466 480 0 FreeSans 448 90 0 0 la_data_in[118]
port 163 nsew signal input
flabel metal2 s 547850 -960 547962 480 0 FreeSans 448 90 0 0 la_data_in[119]
port 164 nsew signal input
flabel metal2 s 164854 -960 164966 480 0 FreeSans 448 90 0 0 la_data_in[11]
port 165 nsew signal input
flabel metal2 s 551438 -960 551550 480 0 FreeSans 448 90 0 0 la_data_in[120]
port 166 nsew signal input
flabel metal2 s 554934 -960 555046 480 0 FreeSans 448 90 0 0 la_data_in[121]
port 167 nsew signal input
flabel metal2 s 558522 -960 558634 480 0 FreeSans 448 90 0 0 la_data_in[122]
port 168 nsew signal input
flabel metal2 s 562018 -960 562130 480 0 FreeSans 448 90 0 0 la_data_in[123]
port 169 nsew signal input
flabel metal2 s 565606 -960 565718 480 0 FreeSans 448 90 0 0 la_data_in[124]
port 170 nsew signal input
flabel metal2 s 569102 -960 569214 480 0 FreeSans 448 90 0 0 la_data_in[125]
port 171 nsew signal input
flabel metal2 s 572690 -960 572802 480 0 FreeSans 448 90 0 0 la_data_in[126]
port 172 nsew signal input
flabel metal2 s 576278 -960 576390 480 0 FreeSans 448 90 0 0 la_data_in[127]
port 173 nsew signal input
flabel metal2 s 168350 -960 168462 480 0 FreeSans 448 90 0 0 la_data_in[12]
port 174 nsew signal input
flabel metal2 s 171938 -960 172050 480 0 FreeSans 448 90 0 0 la_data_in[13]
port 175 nsew signal input
flabel metal2 s 175434 -960 175546 480 0 FreeSans 448 90 0 0 la_data_in[14]
port 176 nsew signal input
flabel metal2 s 179022 -960 179134 480 0 FreeSans 448 90 0 0 la_data_in[15]
port 177 nsew signal input
flabel metal2 s 182518 -960 182630 480 0 FreeSans 448 90 0 0 la_data_in[16]
port 178 nsew signal input
flabel metal2 s 186106 -960 186218 480 0 FreeSans 448 90 0 0 la_data_in[17]
port 179 nsew signal input
flabel metal2 s 189694 -960 189806 480 0 FreeSans 448 90 0 0 la_data_in[18]
port 180 nsew signal input
flabel metal2 s 193190 -960 193302 480 0 FreeSans 448 90 0 0 la_data_in[19]
port 181 nsew signal input
flabel metal2 s 129342 -960 129454 480 0 FreeSans 448 90 0 0 la_data_in[1]
port 182 nsew signal input
flabel metal2 s 196778 -960 196890 480 0 FreeSans 448 90 0 0 la_data_in[20]
port 183 nsew signal input
flabel metal2 s 200274 -960 200386 480 0 FreeSans 448 90 0 0 la_data_in[21]
port 184 nsew signal input
flabel metal2 s 203862 -960 203974 480 0 FreeSans 448 90 0 0 la_data_in[22]
port 185 nsew signal input
flabel metal2 s 207358 -960 207470 480 0 FreeSans 448 90 0 0 la_data_in[23]
port 186 nsew signal input
flabel metal2 s 210946 -960 211058 480 0 FreeSans 448 90 0 0 la_data_in[24]
port 187 nsew signal input
flabel metal2 s 214442 -960 214554 480 0 FreeSans 448 90 0 0 la_data_in[25]
port 188 nsew signal input
flabel metal2 s 218030 -960 218142 480 0 FreeSans 448 90 0 0 la_data_in[26]
port 189 nsew signal input
flabel metal2 s 221526 -960 221638 480 0 FreeSans 448 90 0 0 la_data_in[27]
port 190 nsew signal input
flabel metal2 s 225114 -960 225226 480 0 FreeSans 448 90 0 0 la_data_in[28]
port 191 nsew signal input
flabel metal2 s 228702 -960 228814 480 0 FreeSans 448 90 0 0 la_data_in[29]
port 192 nsew signal input
flabel metal2 s 132930 -960 133042 480 0 FreeSans 448 90 0 0 la_data_in[2]
port 193 nsew signal input
flabel metal2 s 232198 -960 232310 480 0 FreeSans 448 90 0 0 la_data_in[30]
port 194 nsew signal input
flabel metal2 s 235786 -960 235898 480 0 FreeSans 448 90 0 0 la_data_in[31]
port 195 nsew signal input
flabel metal2 s 239282 -960 239394 480 0 FreeSans 448 90 0 0 la_data_in[32]
port 196 nsew signal input
flabel metal2 s 242870 -960 242982 480 0 FreeSans 448 90 0 0 la_data_in[33]
port 197 nsew signal input
flabel metal2 s 246366 -960 246478 480 0 FreeSans 448 90 0 0 la_data_in[34]
port 198 nsew signal input
flabel metal2 s 249954 -960 250066 480 0 FreeSans 448 90 0 0 la_data_in[35]
port 199 nsew signal input
flabel metal2 s 253450 -960 253562 480 0 FreeSans 448 90 0 0 la_data_in[36]
port 200 nsew signal input
flabel metal2 s 257038 -960 257150 480 0 FreeSans 448 90 0 0 la_data_in[37]
port 201 nsew signal input
flabel metal2 s 260626 -960 260738 480 0 FreeSans 448 90 0 0 la_data_in[38]
port 202 nsew signal input
flabel metal2 s 264122 -960 264234 480 0 FreeSans 448 90 0 0 la_data_in[39]
port 203 nsew signal input
flabel metal2 s 136426 -960 136538 480 0 FreeSans 448 90 0 0 la_data_in[3]
port 204 nsew signal input
flabel metal2 s 267710 -960 267822 480 0 FreeSans 448 90 0 0 la_data_in[40]
port 205 nsew signal input
flabel metal2 s 271206 -960 271318 480 0 FreeSans 448 90 0 0 la_data_in[41]
port 206 nsew signal input
flabel metal2 s 274794 -960 274906 480 0 FreeSans 448 90 0 0 la_data_in[42]
port 207 nsew signal input
flabel metal2 s 278290 -960 278402 480 0 FreeSans 448 90 0 0 la_data_in[43]
port 208 nsew signal input
flabel metal2 s 281878 -960 281990 480 0 FreeSans 448 90 0 0 la_data_in[44]
port 209 nsew signal input
flabel metal2 s 285374 -960 285486 480 0 FreeSans 448 90 0 0 la_data_in[45]
port 210 nsew signal input
flabel metal2 s 288962 -960 289074 480 0 FreeSans 448 90 0 0 la_data_in[46]
port 211 nsew signal input
flabel metal2 s 292550 -960 292662 480 0 FreeSans 448 90 0 0 la_data_in[47]
port 212 nsew signal input
flabel metal2 s 296046 -960 296158 480 0 FreeSans 448 90 0 0 la_data_in[48]
port 213 nsew signal input
flabel metal2 s 299634 -960 299746 480 0 FreeSans 448 90 0 0 la_data_in[49]
port 214 nsew signal input
flabel metal2 s 140014 -960 140126 480 0 FreeSans 448 90 0 0 la_data_in[4]
port 215 nsew signal input
flabel metal2 s 303130 -960 303242 480 0 FreeSans 448 90 0 0 la_data_in[50]
port 216 nsew signal input
flabel metal2 s 306718 -960 306830 480 0 FreeSans 448 90 0 0 la_data_in[51]
port 217 nsew signal input
flabel metal2 s 310214 -960 310326 480 0 FreeSans 448 90 0 0 la_data_in[52]
port 218 nsew signal input
flabel metal2 s 313802 -960 313914 480 0 FreeSans 448 90 0 0 la_data_in[53]
port 219 nsew signal input
flabel metal2 s 317298 -960 317410 480 0 FreeSans 448 90 0 0 la_data_in[54]
port 220 nsew signal input
flabel metal2 s 320886 -960 320998 480 0 FreeSans 448 90 0 0 la_data_in[55]
port 221 nsew signal input
flabel metal2 s 324382 -960 324494 480 0 FreeSans 448 90 0 0 la_data_in[56]
port 222 nsew signal input
flabel metal2 s 327970 -960 328082 480 0 FreeSans 448 90 0 0 la_data_in[57]
port 223 nsew signal input
flabel metal2 s 331558 -960 331670 480 0 FreeSans 448 90 0 0 la_data_in[58]
port 224 nsew signal input
flabel metal2 s 335054 -960 335166 480 0 FreeSans 448 90 0 0 la_data_in[59]
port 225 nsew signal input
flabel metal2 s 143510 -960 143622 480 0 FreeSans 448 90 0 0 la_data_in[5]
port 226 nsew signal input
flabel metal2 s 338642 -960 338754 480 0 FreeSans 448 90 0 0 la_data_in[60]
port 227 nsew signal input
flabel metal2 s 342138 -960 342250 480 0 FreeSans 448 90 0 0 la_data_in[61]
port 228 nsew signal input
flabel metal2 s 345726 -960 345838 480 0 FreeSans 448 90 0 0 la_data_in[62]
port 229 nsew signal input
flabel metal2 s 349222 -960 349334 480 0 FreeSans 448 90 0 0 la_data_in[63]
port 230 nsew signal input
flabel metal2 s 352810 -960 352922 480 0 FreeSans 448 90 0 0 la_data_in[64]
port 231 nsew signal input
flabel metal2 s 356306 -960 356418 480 0 FreeSans 448 90 0 0 la_data_in[65]
port 232 nsew signal input
flabel metal2 s 359894 -960 360006 480 0 FreeSans 448 90 0 0 la_data_in[66]
port 233 nsew signal input
flabel metal2 s 363482 -960 363594 480 0 FreeSans 448 90 0 0 la_data_in[67]
port 234 nsew signal input
flabel metal2 s 366978 -960 367090 480 0 FreeSans 448 90 0 0 la_data_in[68]
port 235 nsew signal input
flabel metal2 s 370566 -960 370678 480 0 FreeSans 448 90 0 0 la_data_in[69]
port 236 nsew signal input
flabel metal2 s 147098 -960 147210 480 0 FreeSans 448 90 0 0 la_data_in[6]
port 237 nsew signal input
flabel metal2 s 374062 -960 374174 480 0 FreeSans 448 90 0 0 la_data_in[70]
port 238 nsew signal input
flabel metal2 s 377650 -960 377762 480 0 FreeSans 448 90 0 0 la_data_in[71]
port 239 nsew signal input
flabel metal2 s 381146 -960 381258 480 0 FreeSans 448 90 0 0 la_data_in[72]
port 240 nsew signal input
flabel metal2 s 384734 -960 384846 480 0 FreeSans 448 90 0 0 la_data_in[73]
port 241 nsew signal input
flabel metal2 s 388230 -960 388342 480 0 FreeSans 448 90 0 0 la_data_in[74]
port 242 nsew signal input
flabel metal2 s 391818 -960 391930 480 0 FreeSans 448 90 0 0 la_data_in[75]
port 243 nsew signal input
flabel metal2 s 395314 -960 395426 480 0 FreeSans 448 90 0 0 la_data_in[76]
port 244 nsew signal input
flabel metal2 s 398902 -960 399014 480 0 FreeSans 448 90 0 0 la_data_in[77]
port 245 nsew signal input
flabel metal2 s 402490 -960 402602 480 0 FreeSans 448 90 0 0 la_data_in[78]
port 246 nsew signal input
flabel metal2 s 405986 -960 406098 480 0 FreeSans 448 90 0 0 la_data_in[79]
port 247 nsew signal input
flabel metal2 s 150594 -960 150706 480 0 FreeSans 448 90 0 0 la_data_in[7]
port 248 nsew signal input
flabel metal2 s 409574 -960 409686 480 0 FreeSans 448 90 0 0 la_data_in[80]
port 249 nsew signal input
flabel metal2 s 413070 -960 413182 480 0 FreeSans 448 90 0 0 la_data_in[81]
port 250 nsew signal input
flabel metal2 s 416658 -960 416770 480 0 FreeSans 448 90 0 0 la_data_in[82]
port 251 nsew signal input
flabel metal2 s 420154 -960 420266 480 0 FreeSans 448 90 0 0 la_data_in[83]
port 252 nsew signal input
flabel metal2 s 423742 -960 423854 480 0 FreeSans 448 90 0 0 la_data_in[84]
port 253 nsew signal input
flabel metal2 s 427238 -960 427350 480 0 FreeSans 448 90 0 0 la_data_in[85]
port 254 nsew signal input
flabel metal2 s 430826 -960 430938 480 0 FreeSans 448 90 0 0 la_data_in[86]
port 255 nsew signal input
flabel metal2 s 434414 -960 434526 480 0 FreeSans 448 90 0 0 la_data_in[87]
port 256 nsew signal input
flabel metal2 s 437910 -960 438022 480 0 FreeSans 448 90 0 0 la_data_in[88]
port 257 nsew signal input
flabel metal2 s 441498 -960 441610 480 0 FreeSans 448 90 0 0 la_data_in[89]
port 258 nsew signal input
flabel metal2 s 154182 -960 154294 480 0 FreeSans 448 90 0 0 la_data_in[8]
port 259 nsew signal input
flabel metal2 s 444994 -960 445106 480 0 FreeSans 448 90 0 0 la_data_in[90]
port 260 nsew signal input
flabel metal2 s 448582 -960 448694 480 0 FreeSans 448 90 0 0 la_data_in[91]
port 261 nsew signal input
flabel metal2 s 452078 -960 452190 480 0 FreeSans 448 90 0 0 la_data_in[92]
port 262 nsew signal input
flabel metal2 s 455666 -960 455778 480 0 FreeSans 448 90 0 0 la_data_in[93]
port 263 nsew signal input
flabel metal2 s 459162 -960 459274 480 0 FreeSans 448 90 0 0 la_data_in[94]
port 264 nsew signal input
flabel metal2 s 462750 -960 462862 480 0 FreeSans 448 90 0 0 la_data_in[95]
port 265 nsew signal input
flabel metal2 s 466246 -960 466358 480 0 FreeSans 448 90 0 0 la_data_in[96]
port 266 nsew signal input
flabel metal2 s 469834 -960 469946 480 0 FreeSans 448 90 0 0 la_data_in[97]
port 267 nsew signal input
flabel metal2 s 473422 -960 473534 480 0 FreeSans 448 90 0 0 la_data_in[98]
port 268 nsew signal input
flabel metal2 s 476918 -960 477030 480 0 FreeSans 448 90 0 0 la_data_in[99]
port 269 nsew signal input
flabel metal2 s 157770 -960 157882 480 0 FreeSans 448 90 0 0 la_data_in[9]
port 270 nsew signal input
flabel metal2 s 126950 -960 127062 480 0 FreeSans 448 90 0 0 la_data_out[0]
port 271 nsew signal tristate
flabel metal2 s 481702 -960 481814 480 0 FreeSans 448 90 0 0 la_data_out[100]
port 272 nsew signal tristate
flabel metal2 s 485198 -960 485310 480 0 FreeSans 448 90 0 0 la_data_out[101]
port 273 nsew signal tristate
flabel metal2 s 488786 -960 488898 480 0 FreeSans 448 90 0 0 la_data_out[102]
port 274 nsew signal tristate
flabel metal2 s 492282 -960 492394 480 0 FreeSans 448 90 0 0 la_data_out[103]
port 275 nsew signal tristate
flabel metal2 s 495870 -960 495982 480 0 FreeSans 448 90 0 0 la_data_out[104]
port 276 nsew signal tristate
flabel metal2 s 499366 -960 499478 480 0 FreeSans 448 90 0 0 la_data_out[105]
port 277 nsew signal tristate
flabel metal2 s 502954 -960 503066 480 0 FreeSans 448 90 0 0 la_data_out[106]
port 278 nsew signal tristate
flabel metal2 s 506450 -960 506562 480 0 FreeSans 448 90 0 0 la_data_out[107]
port 279 nsew signal tristate
flabel metal2 s 510038 -960 510150 480 0 FreeSans 448 90 0 0 la_data_out[108]
port 280 nsew signal tristate
flabel metal2 s 513534 -960 513646 480 0 FreeSans 448 90 0 0 la_data_out[109]
port 281 nsew signal tristate
flabel metal2 s 162462 -960 162574 480 0 FreeSans 448 90 0 0 la_data_out[10]
port 282 nsew signal tristate
flabel metal2 s 517122 -960 517234 480 0 FreeSans 448 90 0 0 la_data_out[110]
port 283 nsew signal tristate
flabel metal2 s 520710 -960 520822 480 0 FreeSans 448 90 0 0 la_data_out[111]
port 284 nsew signal tristate
flabel metal2 s 524206 -960 524318 480 0 FreeSans 448 90 0 0 la_data_out[112]
port 285 nsew signal tristate
flabel metal2 s 527794 -960 527906 480 0 FreeSans 448 90 0 0 la_data_out[113]
port 286 nsew signal tristate
flabel metal2 s 531290 -960 531402 480 0 FreeSans 448 90 0 0 la_data_out[114]
port 287 nsew signal tristate
flabel metal2 s 534878 -960 534990 480 0 FreeSans 448 90 0 0 la_data_out[115]
port 288 nsew signal tristate
flabel metal2 s 538374 -960 538486 480 0 FreeSans 448 90 0 0 la_data_out[116]
port 289 nsew signal tristate
flabel metal2 s 541962 -960 542074 480 0 FreeSans 448 90 0 0 la_data_out[117]
port 290 nsew signal tristate
flabel metal2 s 545458 -960 545570 480 0 FreeSans 448 90 0 0 la_data_out[118]
port 291 nsew signal tristate
flabel metal2 s 549046 -960 549158 480 0 FreeSans 448 90 0 0 la_data_out[119]
port 292 nsew signal tristate
flabel metal2 s 166050 -960 166162 480 0 FreeSans 448 90 0 0 la_data_out[11]
port 293 nsew signal tristate
flabel metal2 s 552634 -960 552746 480 0 FreeSans 448 90 0 0 la_data_out[120]
port 294 nsew signal tristate
flabel metal2 s 556130 -960 556242 480 0 FreeSans 448 90 0 0 la_data_out[121]
port 295 nsew signal tristate
flabel metal2 s 559718 -960 559830 480 0 FreeSans 448 90 0 0 la_data_out[122]
port 296 nsew signal tristate
flabel metal2 s 563214 -960 563326 480 0 FreeSans 448 90 0 0 la_data_out[123]
port 297 nsew signal tristate
flabel metal2 s 566802 -960 566914 480 0 FreeSans 448 90 0 0 la_data_out[124]
port 298 nsew signal tristate
flabel metal2 s 570298 -960 570410 480 0 FreeSans 448 90 0 0 la_data_out[125]
port 299 nsew signal tristate
flabel metal2 s 573886 -960 573998 480 0 FreeSans 448 90 0 0 la_data_out[126]
port 300 nsew signal tristate
flabel metal2 s 577382 -960 577494 480 0 FreeSans 448 90 0 0 la_data_out[127]
port 301 nsew signal tristate
flabel metal2 s 169546 -960 169658 480 0 FreeSans 448 90 0 0 la_data_out[12]
port 302 nsew signal tristate
flabel metal2 s 173134 -960 173246 480 0 FreeSans 448 90 0 0 la_data_out[13]
port 303 nsew signal tristate
flabel metal2 s 176630 -960 176742 480 0 FreeSans 448 90 0 0 la_data_out[14]
port 304 nsew signal tristate
flabel metal2 s 180218 -960 180330 480 0 FreeSans 448 90 0 0 la_data_out[15]
port 305 nsew signal tristate
flabel metal2 s 183714 -960 183826 480 0 FreeSans 448 90 0 0 la_data_out[16]
port 306 nsew signal tristate
flabel metal2 s 187302 -960 187414 480 0 FreeSans 448 90 0 0 la_data_out[17]
port 307 nsew signal tristate
flabel metal2 s 190798 -960 190910 480 0 FreeSans 448 90 0 0 la_data_out[18]
port 308 nsew signal tristate
flabel metal2 s 194386 -960 194498 480 0 FreeSans 448 90 0 0 la_data_out[19]
port 309 nsew signal tristate
flabel metal2 s 130538 -960 130650 480 0 FreeSans 448 90 0 0 la_data_out[1]
port 310 nsew signal tristate
flabel metal2 s 197882 -960 197994 480 0 FreeSans 448 90 0 0 la_data_out[20]
port 311 nsew signal tristate
flabel metal2 s 201470 -960 201582 480 0 FreeSans 448 90 0 0 la_data_out[21]
port 312 nsew signal tristate
flabel metal2 s 205058 -960 205170 480 0 FreeSans 448 90 0 0 la_data_out[22]
port 313 nsew signal tristate
flabel metal2 s 208554 -960 208666 480 0 FreeSans 448 90 0 0 la_data_out[23]
port 314 nsew signal tristate
flabel metal2 s 212142 -960 212254 480 0 FreeSans 448 90 0 0 la_data_out[24]
port 315 nsew signal tristate
flabel metal2 s 215638 -960 215750 480 0 FreeSans 448 90 0 0 la_data_out[25]
port 316 nsew signal tristate
flabel metal2 s 219226 -960 219338 480 0 FreeSans 448 90 0 0 la_data_out[26]
port 317 nsew signal tristate
flabel metal2 s 222722 -960 222834 480 0 FreeSans 448 90 0 0 la_data_out[27]
port 318 nsew signal tristate
flabel metal2 s 226310 -960 226422 480 0 FreeSans 448 90 0 0 la_data_out[28]
port 319 nsew signal tristate
flabel metal2 s 229806 -960 229918 480 0 FreeSans 448 90 0 0 la_data_out[29]
port 320 nsew signal tristate
flabel metal2 s 134126 -960 134238 480 0 FreeSans 448 90 0 0 la_data_out[2]
port 321 nsew signal tristate
flabel metal2 s 233394 -960 233506 480 0 FreeSans 448 90 0 0 la_data_out[30]
port 322 nsew signal tristate
flabel metal2 s 236982 -960 237094 480 0 FreeSans 448 90 0 0 la_data_out[31]
port 323 nsew signal tristate
flabel metal2 s 240478 -960 240590 480 0 FreeSans 448 90 0 0 la_data_out[32]
port 324 nsew signal tristate
flabel metal2 s 244066 -960 244178 480 0 FreeSans 448 90 0 0 la_data_out[33]
port 325 nsew signal tristate
flabel metal2 s 247562 -960 247674 480 0 FreeSans 448 90 0 0 la_data_out[34]
port 326 nsew signal tristate
flabel metal2 s 251150 -960 251262 480 0 FreeSans 448 90 0 0 la_data_out[35]
port 327 nsew signal tristate
flabel metal2 s 254646 -960 254758 480 0 FreeSans 448 90 0 0 la_data_out[36]
port 328 nsew signal tristate
flabel metal2 s 258234 -960 258346 480 0 FreeSans 448 90 0 0 la_data_out[37]
port 329 nsew signal tristate
flabel metal2 s 261730 -960 261842 480 0 FreeSans 448 90 0 0 la_data_out[38]
port 330 nsew signal tristate
flabel metal2 s 265318 -960 265430 480 0 FreeSans 448 90 0 0 la_data_out[39]
port 331 nsew signal tristate
flabel metal2 s 137622 -960 137734 480 0 FreeSans 448 90 0 0 la_data_out[3]
port 332 nsew signal tristate
flabel metal2 s 268814 -960 268926 480 0 FreeSans 448 90 0 0 la_data_out[40]
port 333 nsew signal tristate
flabel metal2 s 272402 -960 272514 480 0 FreeSans 448 90 0 0 la_data_out[41]
port 334 nsew signal tristate
flabel metal2 s 275990 -960 276102 480 0 FreeSans 448 90 0 0 la_data_out[42]
port 335 nsew signal tristate
flabel metal2 s 279486 -960 279598 480 0 FreeSans 448 90 0 0 la_data_out[43]
port 336 nsew signal tristate
flabel metal2 s 283074 -960 283186 480 0 FreeSans 448 90 0 0 la_data_out[44]
port 337 nsew signal tristate
flabel metal2 s 286570 -960 286682 480 0 FreeSans 448 90 0 0 la_data_out[45]
port 338 nsew signal tristate
flabel metal2 s 290158 -960 290270 480 0 FreeSans 448 90 0 0 la_data_out[46]
port 339 nsew signal tristate
flabel metal2 s 293654 -960 293766 480 0 FreeSans 448 90 0 0 la_data_out[47]
port 340 nsew signal tristate
flabel metal2 s 297242 -960 297354 480 0 FreeSans 448 90 0 0 la_data_out[48]
port 341 nsew signal tristate
flabel metal2 s 300738 -960 300850 480 0 FreeSans 448 90 0 0 la_data_out[49]
port 342 nsew signal tristate
flabel metal2 s 141210 -960 141322 480 0 FreeSans 448 90 0 0 la_data_out[4]
port 343 nsew signal tristate
flabel metal2 s 304326 -960 304438 480 0 FreeSans 448 90 0 0 la_data_out[50]
port 344 nsew signal tristate
flabel metal2 s 307914 -960 308026 480 0 FreeSans 448 90 0 0 la_data_out[51]
port 345 nsew signal tristate
flabel metal2 s 311410 -960 311522 480 0 FreeSans 448 90 0 0 la_data_out[52]
port 346 nsew signal tristate
flabel metal2 s 314998 -960 315110 480 0 FreeSans 448 90 0 0 la_data_out[53]
port 347 nsew signal tristate
flabel metal2 s 318494 -960 318606 480 0 FreeSans 448 90 0 0 la_data_out[54]
port 348 nsew signal tristate
flabel metal2 s 322082 -960 322194 480 0 FreeSans 448 90 0 0 la_data_out[55]
port 349 nsew signal tristate
flabel metal2 s 325578 -960 325690 480 0 FreeSans 448 90 0 0 la_data_out[56]
port 350 nsew signal tristate
flabel metal2 s 329166 -960 329278 480 0 FreeSans 448 90 0 0 la_data_out[57]
port 351 nsew signal tristate
flabel metal2 s 332662 -960 332774 480 0 FreeSans 448 90 0 0 la_data_out[58]
port 352 nsew signal tristate
flabel metal2 s 336250 -960 336362 480 0 FreeSans 448 90 0 0 la_data_out[59]
port 353 nsew signal tristate
flabel metal2 s 144706 -960 144818 480 0 FreeSans 448 90 0 0 la_data_out[5]
port 354 nsew signal tristate
flabel metal2 s 339838 -960 339950 480 0 FreeSans 448 90 0 0 la_data_out[60]
port 355 nsew signal tristate
flabel metal2 s 343334 -960 343446 480 0 FreeSans 448 90 0 0 la_data_out[61]
port 356 nsew signal tristate
flabel metal2 s 346922 -960 347034 480 0 FreeSans 448 90 0 0 la_data_out[62]
port 357 nsew signal tristate
flabel metal2 s 350418 -960 350530 480 0 FreeSans 448 90 0 0 la_data_out[63]
port 358 nsew signal tristate
flabel metal2 s 354006 -960 354118 480 0 FreeSans 448 90 0 0 la_data_out[64]
port 359 nsew signal tristate
flabel metal2 s 357502 -960 357614 480 0 FreeSans 448 90 0 0 la_data_out[65]
port 360 nsew signal tristate
flabel metal2 s 361090 -960 361202 480 0 FreeSans 448 90 0 0 la_data_out[66]
port 361 nsew signal tristate
flabel metal2 s 364586 -960 364698 480 0 FreeSans 448 90 0 0 la_data_out[67]
port 362 nsew signal tristate
flabel metal2 s 368174 -960 368286 480 0 FreeSans 448 90 0 0 la_data_out[68]
port 363 nsew signal tristate
flabel metal2 s 371670 -960 371782 480 0 FreeSans 448 90 0 0 la_data_out[69]
port 364 nsew signal tristate
flabel metal2 s 148294 -960 148406 480 0 FreeSans 448 90 0 0 la_data_out[6]
port 365 nsew signal tristate
flabel metal2 s 375258 -960 375370 480 0 FreeSans 448 90 0 0 la_data_out[70]
port 366 nsew signal tristate
flabel metal2 s 378846 -960 378958 480 0 FreeSans 448 90 0 0 la_data_out[71]
port 367 nsew signal tristate
flabel metal2 s 382342 -960 382454 480 0 FreeSans 448 90 0 0 la_data_out[72]
port 368 nsew signal tristate
flabel metal2 s 385930 -960 386042 480 0 FreeSans 448 90 0 0 la_data_out[73]
port 369 nsew signal tristate
flabel metal2 s 389426 -960 389538 480 0 FreeSans 448 90 0 0 la_data_out[74]
port 370 nsew signal tristate
flabel metal2 s 393014 -960 393126 480 0 FreeSans 448 90 0 0 la_data_out[75]
port 371 nsew signal tristate
flabel metal2 s 396510 -960 396622 480 0 FreeSans 448 90 0 0 la_data_out[76]
port 372 nsew signal tristate
flabel metal2 s 400098 -960 400210 480 0 FreeSans 448 90 0 0 la_data_out[77]
port 373 nsew signal tristate
flabel metal2 s 403594 -960 403706 480 0 FreeSans 448 90 0 0 la_data_out[78]
port 374 nsew signal tristate
flabel metal2 s 407182 -960 407294 480 0 FreeSans 448 90 0 0 la_data_out[79]
port 375 nsew signal tristate
flabel metal2 s 151790 -960 151902 480 0 FreeSans 448 90 0 0 la_data_out[7]
port 376 nsew signal tristate
flabel metal2 s 410770 -960 410882 480 0 FreeSans 448 90 0 0 la_data_out[80]
port 377 nsew signal tristate
flabel metal2 s 414266 -960 414378 480 0 FreeSans 448 90 0 0 la_data_out[81]
port 378 nsew signal tristate
flabel metal2 s 417854 -960 417966 480 0 FreeSans 448 90 0 0 la_data_out[82]
port 379 nsew signal tristate
flabel metal2 s 421350 -960 421462 480 0 FreeSans 448 90 0 0 la_data_out[83]
port 380 nsew signal tristate
flabel metal2 s 424938 -960 425050 480 0 FreeSans 448 90 0 0 la_data_out[84]
port 381 nsew signal tristate
flabel metal2 s 428434 -960 428546 480 0 FreeSans 448 90 0 0 la_data_out[85]
port 382 nsew signal tristate
flabel metal2 s 432022 -960 432134 480 0 FreeSans 448 90 0 0 la_data_out[86]
port 383 nsew signal tristate
flabel metal2 s 435518 -960 435630 480 0 FreeSans 448 90 0 0 la_data_out[87]
port 384 nsew signal tristate
flabel metal2 s 439106 -960 439218 480 0 FreeSans 448 90 0 0 la_data_out[88]
port 385 nsew signal tristate
flabel metal2 s 442602 -960 442714 480 0 FreeSans 448 90 0 0 la_data_out[89]
port 386 nsew signal tristate
flabel metal2 s 155378 -960 155490 480 0 FreeSans 448 90 0 0 la_data_out[8]
port 387 nsew signal tristate
flabel metal2 s 446190 -960 446302 480 0 FreeSans 448 90 0 0 la_data_out[90]
port 388 nsew signal tristate
flabel metal2 s 449778 -960 449890 480 0 FreeSans 448 90 0 0 la_data_out[91]
port 389 nsew signal tristate
flabel metal2 s 453274 -960 453386 480 0 FreeSans 448 90 0 0 la_data_out[92]
port 390 nsew signal tristate
flabel metal2 s 456862 -960 456974 480 0 FreeSans 448 90 0 0 la_data_out[93]
port 391 nsew signal tristate
flabel metal2 s 460358 -960 460470 480 0 FreeSans 448 90 0 0 la_data_out[94]
port 392 nsew signal tristate
flabel metal2 s 463946 -960 464058 480 0 FreeSans 448 90 0 0 la_data_out[95]
port 393 nsew signal tristate
flabel metal2 s 467442 -960 467554 480 0 FreeSans 448 90 0 0 la_data_out[96]
port 394 nsew signal tristate
flabel metal2 s 471030 -960 471142 480 0 FreeSans 448 90 0 0 la_data_out[97]
port 395 nsew signal tristate
flabel metal2 s 474526 -960 474638 480 0 FreeSans 448 90 0 0 la_data_out[98]
port 396 nsew signal tristate
flabel metal2 s 478114 -960 478226 480 0 FreeSans 448 90 0 0 la_data_out[99]
port 397 nsew signal tristate
flabel metal2 s 158874 -960 158986 480 0 FreeSans 448 90 0 0 la_data_out[9]
port 398 nsew signal tristate
flabel metal2 s 128146 -960 128258 480 0 FreeSans 448 90 0 0 la_oenb[0]
port 399 nsew signal input
flabel metal2 s 482806 -960 482918 480 0 FreeSans 448 90 0 0 la_oenb[100]
port 400 nsew signal input
flabel metal2 s 486394 -960 486506 480 0 FreeSans 448 90 0 0 la_oenb[101]
port 401 nsew signal input
flabel metal2 s 489890 -960 490002 480 0 FreeSans 448 90 0 0 la_oenb[102]
port 402 nsew signal input
flabel metal2 s 493478 -960 493590 480 0 FreeSans 448 90 0 0 la_oenb[103]
port 403 nsew signal input
flabel metal2 s 497066 -960 497178 480 0 FreeSans 448 90 0 0 la_oenb[104]
port 404 nsew signal input
flabel metal2 s 500562 -960 500674 480 0 FreeSans 448 90 0 0 la_oenb[105]
port 405 nsew signal input
flabel metal2 s 504150 -960 504262 480 0 FreeSans 448 90 0 0 la_oenb[106]
port 406 nsew signal input
flabel metal2 s 507646 -960 507758 480 0 FreeSans 448 90 0 0 la_oenb[107]
port 407 nsew signal input
flabel metal2 s 511234 -960 511346 480 0 FreeSans 448 90 0 0 la_oenb[108]
port 408 nsew signal input
flabel metal2 s 514730 -960 514842 480 0 FreeSans 448 90 0 0 la_oenb[109]
port 409 nsew signal input
flabel metal2 s 163658 -960 163770 480 0 FreeSans 448 90 0 0 la_oenb[10]
port 410 nsew signal input
flabel metal2 s 518318 -960 518430 480 0 FreeSans 448 90 0 0 la_oenb[110]
port 411 nsew signal input
flabel metal2 s 521814 -960 521926 480 0 FreeSans 448 90 0 0 la_oenb[111]
port 412 nsew signal input
flabel metal2 s 525402 -960 525514 480 0 FreeSans 448 90 0 0 la_oenb[112]
port 413 nsew signal input
flabel metal2 s 528990 -960 529102 480 0 FreeSans 448 90 0 0 la_oenb[113]
port 414 nsew signal input
flabel metal2 s 532486 -960 532598 480 0 FreeSans 448 90 0 0 la_oenb[114]
port 415 nsew signal input
flabel metal2 s 536074 -960 536186 480 0 FreeSans 448 90 0 0 la_oenb[115]
port 416 nsew signal input
flabel metal2 s 539570 -960 539682 480 0 FreeSans 448 90 0 0 la_oenb[116]
port 417 nsew signal input
flabel metal2 s 543158 -960 543270 480 0 FreeSans 448 90 0 0 la_oenb[117]
port 418 nsew signal input
flabel metal2 s 546654 -960 546766 480 0 FreeSans 448 90 0 0 la_oenb[118]
port 419 nsew signal input
flabel metal2 s 550242 -960 550354 480 0 FreeSans 448 90 0 0 la_oenb[119]
port 420 nsew signal input
flabel metal2 s 167154 -960 167266 480 0 FreeSans 448 90 0 0 la_oenb[11]
port 421 nsew signal input
flabel metal2 s 553738 -960 553850 480 0 FreeSans 448 90 0 0 la_oenb[120]
port 422 nsew signal input
flabel metal2 s 557326 -960 557438 480 0 FreeSans 448 90 0 0 la_oenb[121]
port 423 nsew signal input
flabel metal2 s 560822 -960 560934 480 0 FreeSans 448 90 0 0 la_oenb[122]
port 424 nsew signal input
flabel metal2 s 564410 -960 564522 480 0 FreeSans 448 90 0 0 la_oenb[123]
port 425 nsew signal input
flabel metal2 s 567998 -960 568110 480 0 FreeSans 448 90 0 0 la_oenb[124]
port 426 nsew signal input
flabel metal2 s 571494 -960 571606 480 0 FreeSans 448 90 0 0 la_oenb[125]
port 427 nsew signal input
flabel metal2 s 575082 -960 575194 480 0 FreeSans 448 90 0 0 la_oenb[126]
port 428 nsew signal input
flabel metal2 s 578578 -960 578690 480 0 FreeSans 448 90 0 0 la_oenb[127]
port 429 nsew signal input
flabel metal2 s 170742 -960 170854 480 0 FreeSans 448 90 0 0 la_oenb[12]
port 430 nsew signal input
flabel metal2 s 174238 -960 174350 480 0 FreeSans 448 90 0 0 la_oenb[13]
port 431 nsew signal input
flabel metal2 s 177826 -960 177938 480 0 FreeSans 448 90 0 0 la_oenb[14]
port 432 nsew signal input
flabel metal2 s 181414 -960 181526 480 0 FreeSans 448 90 0 0 la_oenb[15]
port 433 nsew signal input
flabel metal2 s 184910 -960 185022 480 0 FreeSans 448 90 0 0 la_oenb[16]
port 434 nsew signal input
flabel metal2 s 188498 -960 188610 480 0 FreeSans 448 90 0 0 la_oenb[17]
port 435 nsew signal input
flabel metal2 s 191994 -960 192106 480 0 FreeSans 448 90 0 0 la_oenb[18]
port 436 nsew signal input
flabel metal2 s 195582 -960 195694 480 0 FreeSans 448 90 0 0 la_oenb[19]
port 437 nsew signal input
flabel metal2 s 131734 -960 131846 480 0 FreeSans 448 90 0 0 la_oenb[1]
port 438 nsew signal input
flabel metal2 s 199078 -960 199190 480 0 FreeSans 448 90 0 0 la_oenb[20]
port 439 nsew signal input
flabel metal2 s 202666 -960 202778 480 0 FreeSans 448 90 0 0 la_oenb[21]
port 440 nsew signal input
flabel metal2 s 206162 -960 206274 480 0 FreeSans 448 90 0 0 la_oenb[22]
port 441 nsew signal input
flabel metal2 s 209750 -960 209862 480 0 FreeSans 448 90 0 0 la_oenb[23]
port 442 nsew signal input
flabel metal2 s 213338 -960 213450 480 0 FreeSans 448 90 0 0 la_oenb[24]
port 443 nsew signal input
flabel metal2 s 216834 -960 216946 480 0 FreeSans 448 90 0 0 la_oenb[25]
port 444 nsew signal input
flabel metal2 s 220422 -960 220534 480 0 FreeSans 448 90 0 0 la_oenb[26]
port 445 nsew signal input
flabel metal2 s 223918 -960 224030 480 0 FreeSans 448 90 0 0 la_oenb[27]
port 446 nsew signal input
flabel metal2 s 227506 -960 227618 480 0 FreeSans 448 90 0 0 la_oenb[28]
port 447 nsew signal input
flabel metal2 s 231002 -960 231114 480 0 FreeSans 448 90 0 0 la_oenb[29]
port 448 nsew signal input
flabel metal2 s 135230 -960 135342 480 0 FreeSans 448 90 0 0 la_oenb[2]
port 449 nsew signal input
flabel metal2 s 234590 -960 234702 480 0 FreeSans 448 90 0 0 la_oenb[30]
port 450 nsew signal input
flabel metal2 s 238086 -960 238198 480 0 FreeSans 448 90 0 0 la_oenb[31]
port 451 nsew signal input
flabel metal2 s 241674 -960 241786 480 0 FreeSans 448 90 0 0 la_oenb[32]
port 452 nsew signal input
flabel metal2 s 245170 -960 245282 480 0 FreeSans 448 90 0 0 la_oenb[33]
port 453 nsew signal input
flabel metal2 s 248758 -960 248870 480 0 FreeSans 448 90 0 0 la_oenb[34]
port 454 nsew signal input
flabel metal2 s 252346 -960 252458 480 0 FreeSans 448 90 0 0 la_oenb[35]
port 455 nsew signal input
flabel metal2 s 255842 -960 255954 480 0 FreeSans 448 90 0 0 la_oenb[36]
port 456 nsew signal input
flabel metal2 s 259430 -960 259542 480 0 FreeSans 448 90 0 0 la_oenb[37]
port 457 nsew signal input
flabel metal2 s 262926 -960 263038 480 0 FreeSans 448 90 0 0 la_oenb[38]
port 458 nsew signal input
flabel metal2 s 266514 -960 266626 480 0 FreeSans 448 90 0 0 la_oenb[39]
port 459 nsew signal input
flabel metal2 s 138818 -960 138930 480 0 FreeSans 448 90 0 0 la_oenb[3]
port 460 nsew signal input
flabel metal2 s 270010 -960 270122 480 0 FreeSans 448 90 0 0 la_oenb[40]
port 461 nsew signal input
flabel metal2 s 273598 -960 273710 480 0 FreeSans 448 90 0 0 la_oenb[41]
port 462 nsew signal input
flabel metal2 s 277094 -960 277206 480 0 FreeSans 448 90 0 0 la_oenb[42]
port 463 nsew signal input
flabel metal2 s 280682 -960 280794 480 0 FreeSans 448 90 0 0 la_oenb[43]
port 464 nsew signal input
flabel metal2 s 284270 -960 284382 480 0 FreeSans 448 90 0 0 la_oenb[44]
port 465 nsew signal input
flabel metal2 s 287766 -960 287878 480 0 FreeSans 448 90 0 0 la_oenb[45]
port 466 nsew signal input
flabel metal2 s 291354 -960 291466 480 0 FreeSans 448 90 0 0 la_oenb[46]
port 467 nsew signal input
flabel metal2 s 294850 -960 294962 480 0 FreeSans 448 90 0 0 la_oenb[47]
port 468 nsew signal input
flabel metal2 s 298438 -960 298550 480 0 FreeSans 448 90 0 0 la_oenb[48]
port 469 nsew signal input
flabel metal2 s 301934 -960 302046 480 0 FreeSans 448 90 0 0 la_oenb[49]
port 470 nsew signal input
flabel metal2 s 142406 -960 142518 480 0 FreeSans 448 90 0 0 la_oenb[4]
port 471 nsew signal input
flabel metal2 s 305522 -960 305634 480 0 FreeSans 448 90 0 0 la_oenb[50]
port 472 nsew signal input
flabel metal2 s 309018 -960 309130 480 0 FreeSans 448 90 0 0 la_oenb[51]
port 473 nsew signal input
flabel metal2 s 312606 -960 312718 480 0 FreeSans 448 90 0 0 la_oenb[52]
port 474 nsew signal input
flabel metal2 s 316194 -960 316306 480 0 FreeSans 448 90 0 0 la_oenb[53]
port 475 nsew signal input
flabel metal2 s 319690 -960 319802 480 0 FreeSans 448 90 0 0 la_oenb[54]
port 476 nsew signal input
flabel metal2 s 323278 -960 323390 480 0 FreeSans 448 90 0 0 la_oenb[55]
port 477 nsew signal input
flabel metal2 s 326774 -960 326886 480 0 FreeSans 448 90 0 0 la_oenb[56]
port 478 nsew signal input
flabel metal2 s 330362 -960 330474 480 0 FreeSans 448 90 0 0 la_oenb[57]
port 479 nsew signal input
flabel metal2 s 333858 -960 333970 480 0 FreeSans 448 90 0 0 la_oenb[58]
port 480 nsew signal input
flabel metal2 s 337446 -960 337558 480 0 FreeSans 448 90 0 0 la_oenb[59]
port 481 nsew signal input
flabel metal2 s 145902 -960 146014 480 0 FreeSans 448 90 0 0 la_oenb[5]
port 482 nsew signal input
flabel metal2 s 340942 -960 341054 480 0 FreeSans 448 90 0 0 la_oenb[60]
port 483 nsew signal input
flabel metal2 s 344530 -960 344642 480 0 FreeSans 448 90 0 0 la_oenb[61]
port 484 nsew signal input
flabel metal2 s 348026 -960 348138 480 0 FreeSans 448 90 0 0 la_oenb[62]
port 485 nsew signal input
flabel metal2 s 351614 -960 351726 480 0 FreeSans 448 90 0 0 la_oenb[63]
port 486 nsew signal input
flabel metal2 s 355202 -960 355314 480 0 FreeSans 448 90 0 0 la_oenb[64]
port 487 nsew signal input
flabel metal2 s 358698 -960 358810 480 0 FreeSans 448 90 0 0 la_oenb[65]
port 488 nsew signal input
flabel metal2 s 362286 -960 362398 480 0 FreeSans 448 90 0 0 la_oenb[66]
port 489 nsew signal input
flabel metal2 s 365782 -960 365894 480 0 FreeSans 448 90 0 0 la_oenb[67]
port 490 nsew signal input
flabel metal2 s 369370 -960 369482 480 0 FreeSans 448 90 0 0 la_oenb[68]
port 491 nsew signal input
flabel metal2 s 372866 -960 372978 480 0 FreeSans 448 90 0 0 la_oenb[69]
port 492 nsew signal input
flabel metal2 s 149490 -960 149602 480 0 FreeSans 448 90 0 0 la_oenb[6]
port 493 nsew signal input
flabel metal2 s 376454 -960 376566 480 0 FreeSans 448 90 0 0 la_oenb[70]
port 494 nsew signal input
flabel metal2 s 379950 -960 380062 480 0 FreeSans 448 90 0 0 la_oenb[71]
port 495 nsew signal input
flabel metal2 s 383538 -960 383650 480 0 FreeSans 448 90 0 0 la_oenb[72]
port 496 nsew signal input
flabel metal2 s 387126 -960 387238 480 0 FreeSans 448 90 0 0 la_oenb[73]
port 497 nsew signal input
flabel metal2 s 390622 -960 390734 480 0 FreeSans 448 90 0 0 la_oenb[74]
port 498 nsew signal input
flabel metal2 s 394210 -960 394322 480 0 FreeSans 448 90 0 0 la_oenb[75]
port 499 nsew signal input
flabel metal2 s 397706 -960 397818 480 0 FreeSans 448 90 0 0 la_oenb[76]
port 500 nsew signal input
flabel metal2 s 401294 -960 401406 480 0 FreeSans 448 90 0 0 la_oenb[77]
port 501 nsew signal input
flabel metal2 s 404790 -960 404902 480 0 FreeSans 448 90 0 0 la_oenb[78]
port 502 nsew signal input
flabel metal2 s 408378 -960 408490 480 0 FreeSans 448 90 0 0 la_oenb[79]
port 503 nsew signal input
flabel metal2 s 152986 -960 153098 480 0 FreeSans 448 90 0 0 la_oenb[7]
port 504 nsew signal input
flabel metal2 s 411874 -960 411986 480 0 FreeSans 448 90 0 0 la_oenb[80]
port 505 nsew signal input
flabel metal2 s 415462 -960 415574 480 0 FreeSans 448 90 0 0 la_oenb[81]
port 506 nsew signal input
flabel metal2 s 418958 -960 419070 480 0 FreeSans 448 90 0 0 la_oenb[82]
port 507 nsew signal input
flabel metal2 s 422546 -960 422658 480 0 FreeSans 448 90 0 0 la_oenb[83]
port 508 nsew signal input
flabel metal2 s 426134 -960 426246 480 0 FreeSans 448 90 0 0 la_oenb[84]
port 509 nsew signal input
flabel metal2 s 429630 -960 429742 480 0 FreeSans 448 90 0 0 la_oenb[85]
port 510 nsew signal input
flabel metal2 s 433218 -960 433330 480 0 FreeSans 448 90 0 0 la_oenb[86]
port 511 nsew signal input
flabel metal2 s 436714 -960 436826 480 0 FreeSans 448 90 0 0 la_oenb[87]
port 512 nsew signal input
flabel metal2 s 440302 -960 440414 480 0 FreeSans 448 90 0 0 la_oenb[88]
port 513 nsew signal input
flabel metal2 s 443798 -960 443910 480 0 FreeSans 448 90 0 0 la_oenb[89]
port 514 nsew signal input
flabel metal2 s 156574 -960 156686 480 0 FreeSans 448 90 0 0 la_oenb[8]
port 515 nsew signal input
flabel metal2 s 447386 -960 447498 480 0 FreeSans 448 90 0 0 la_oenb[90]
port 516 nsew signal input
flabel metal2 s 450882 -960 450994 480 0 FreeSans 448 90 0 0 la_oenb[91]
port 517 nsew signal input
flabel metal2 s 454470 -960 454582 480 0 FreeSans 448 90 0 0 la_oenb[92]
port 518 nsew signal input
flabel metal2 s 458058 -960 458170 480 0 FreeSans 448 90 0 0 la_oenb[93]
port 519 nsew signal input
flabel metal2 s 461554 -960 461666 480 0 FreeSans 448 90 0 0 la_oenb[94]
port 520 nsew signal input
flabel metal2 s 465142 -960 465254 480 0 FreeSans 448 90 0 0 la_oenb[95]
port 521 nsew signal input
flabel metal2 s 468638 -960 468750 480 0 FreeSans 448 90 0 0 la_oenb[96]
port 522 nsew signal input
flabel metal2 s 472226 -960 472338 480 0 FreeSans 448 90 0 0 la_oenb[97]
port 523 nsew signal input
flabel metal2 s 475722 -960 475834 480 0 FreeSans 448 90 0 0 la_oenb[98]
port 524 nsew signal input
flabel metal2 s 479310 -960 479422 480 0 FreeSans 448 90 0 0 la_oenb[99]
port 525 nsew signal input
flabel metal2 s 160070 -960 160182 480 0 FreeSans 448 90 0 0 la_oenb[9]
port 526 nsew signal input
flabel metal2 s 579774 -960 579886 480 0 FreeSans 448 90 0 0 user_clock2
port 527 nsew signal input
flabel metal2 s 580970 -960 581082 480 0 FreeSans 448 90 0 0 user_irq[0]
port 528 nsew signal tristate
flabel metal2 s 582166 -960 582278 480 0 FreeSans 448 90 0 0 user_irq[1]
port 529 nsew signal tristate
flabel metal2 s 583362 -960 583474 480 0 FreeSans 448 90 0 0 user_irq[2]
port 530 nsew signal tristate
flabel metal4 s -2006 -934 -1386 704870 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -2006 -934 585930 -314 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -2006 704250 585930 704870 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 585310 -934 585930 704870 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 41714 -7654 42334 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 69714 -7654 70334 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 97714 -7654 98334 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 125714 53748 126334 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 153714 -7654 154334 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 181714 -7654 182334 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 209714 -7654 210334 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 237714 54481 238334 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 265714 53748 266334 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 293714 -7654 294334 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 321714 -7654 322334 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 349714 -7654 350334 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 377714 -7654 378334 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 405714 -7654 406334 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 433714 -7654 434334 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 461714 -7654 462334 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 489714 -7654 490334 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 517714 -7654 518334 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 545714 -7654 546334 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 573714 -7654 574334 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 31586 592650 32206 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 68586 592650 69206 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 105586 592650 106206 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 142586 592650 143206 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 179586 592650 180206 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 216586 592650 217206 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 253586 592650 254206 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 290586 592650 291206 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 327586 592650 328206 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 364586 592650 365206 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 401586 592650 402206 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 438586 592650 439206 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 475586 592650 476206 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 512586 592650 513206 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 549586 592650 550206 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 586586 592650 587206 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 623586 592650 624206 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 660586 592650 661206 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 697586 592650 698206 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s -3926 -2854 -3306 706790 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -3926 -2854 587850 -2234 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -3926 706170 587850 706790 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 587230 -2854 587850 706790 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s -5846 -4774 -5226 708710 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -5846 -4774 589770 -4154 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -5846 708090 589770 708710 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 589150 -4774 589770 708710 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s -7766 -6694 -7146 710630 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -7766 -6694 591690 -6074 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -7766 710010 591690 710630 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 591070 -6694 591690 710630 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s -6806 -5734 -6186 709670 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -6806 -5734 590730 -5114 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -6806 709050 590730 709670 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 590110 -5734 590730 709670 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s -8726 -7654 -8106 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 -7654 592650 -7034 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 710970 592650 711590 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 592030 -7654 592650 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s -2966 -1894 -2346 705830 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -2966 -1894 586890 -1274 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -2966 705210 586890 705830 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 586270 -1894 586890 705830 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 37994 -7654 38614 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 65994 -7654 66614 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 93994 43956 94614 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 121994 -7654 122614 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 149994 -7654 150614 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 177994 -7654 178614 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 205994 -7654 206614 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 233994 54481 234614 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 261994 53393 262614 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 289994 -7654 290614 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 317994 -7654 318614 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 345994 -7654 346614 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 373994 -7654 374614 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 401994 -7654 402614 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 429994 -7654 430614 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 457994 -7654 458614 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 485994 -7654 486614 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 513994 -7654 514614 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 541994 -7654 542614 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 569994 -7654 570614 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 27866 592650 28486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 64866 592650 65486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 101866 592650 102486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 138866 592650 139486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 175866 592650 176486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 212866 592650 213486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 249866 592650 250486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 286866 592650 287486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 323866 592650 324486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 360866 592650 361486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 397866 592650 398486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 434866 592650 435486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 471866 592650 472486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 508866 592650 509486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 545866 592650 546486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 582866 592650 583486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 619866 592650 620486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 656866 592650 657486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 693866 592650 694486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s -4886 -3814 -4266 707750 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -4886 -3814 588810 -3194 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -4886 707130 588810 707750 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 588190 -3814 588810 707750 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal2 s 542 -960 654 480 0 FreeSans 448 90 0 0 wb_clk_i
port 539 nsew signal input
flabel metal2 s 1646 -960 1758 480 0 FreeSans 448 90 0 0 wb_rst_i
port 540 nsew signal input
flabel metal2 s 2842 -960 2954 480 0 FreeSans 448 90 0 0 wbs_ack_o
port 541 nsew signal tristate
flabel metal2 s 7626 -960 7738 480 0 FreeSans 448 90 0 0 wbs_adr_i[0]
port 542 nsew signal input
flabel metal2 s 47830 -960 47942 480 0 FreeSans 448 90 0 0 wbs_adr_i[10]
port 543 nsew signal input
flabel metal2 s 51326 -960 51438 480 0 FreeSans 448 90 0 0 wbs_adr_i[11]
port 544 nsew signal input
flabel metal2 s 54914 -960 55026 480 0 FreeSans 448 90 0 0 wbs_adr_i[12]
port 545 nsew signal input
flabel metal2 s 58410 -960 58522 480 0 FreeSans 448 90 0 0 wbs_adr_i[13]
port 546 nsew signal input
flabel metal2 s 61998 -960 62110 480 0 FreeSans 448 90 0 0 wbs_adr_i[14]
port 547 nsew signal input
flabel metal2 s 65494 -960 65606 480 0 FreeSans 448 90 0 0 wbs_adr_i[15]
port 548 nsew signal input
flabel metal2 s 69082 -960 69194 480 0 FreeSans 448 90 0 0 wbs_adr_i[16]
port 549 nsew signal input
flabel metal2 s 72578 -960 72690 480 0 FreeSans 448 90 0 0 wbs_adr_i[17]
port 550 nsew signal input
flabel metal2 s 76166 -960 76278 480 0 FreeSans 448 90 0 0 wbs_adr_i[18]
port 551 nsew signal input
flabel metal2 s 79662 -960 79774 480 0 FreeSans 448 90 0 0 wbs_adr_i[19]
port 552 nsew signal input
flabel metal2 s 12318 -960 12430 480 0 FreeSans 448 90 0 0 wbs_adr_i[1]
port 553 nsew signal input
flabel metal2 s 83250 -960 83362 480 0 FreeSans 448 90 0 0 wbs_adr_i[20]
port 554 nsew signal input
flabel metal2 s 86838 -960 86950 480 0 FreeSans 448 90 0 0 wbs_adr_i[21]
port 555 nsew signal input
flabel metal2 s 90334 -960 90446 480 0 FreeSans 448 90 0 0 wbs_adr_i[22]
port 556 nsew signal input
flabel metal2 s 93922 -960 94034 480 0 FreeSans 448 90 0 0 wbs_adr_i[23]
port 557 nsew signal input
flabel metal2 s 97418 -960 97530 480 0 FreeSans 448 90 0 0 wbs_adr_i[24]
port 558 nsew signal input
flabel metal2 s 101006 -960 101118 480 0 FreeSans 448 90 0 0 wbs_adr_i[25]
port 559 nsew signal input
flabel metal2 s 104502 -960 104614 480 0 FreeSans 448 90 0 0 wbs_adr_i[26]
port 560 nsew signal input
flabel metal2 s 108090 -960 108202 480 0 FreeSans 448 90 0 0 wbs_adr_i[27]
port 561 nsew signal input
flabel metal2 s 111586 -960 111698 480 0 FreeSans 448 90 0 0 wbs_adr_i[28]
port 562 nsew signal input
flabel metal2 s 115174 -960 115286 480 0 FreeSans 448 90 0 0 wbs_adr_i[29]
port 563 nsew signal input
flabel metal2 s 17010 -960 17122 480 0 FreeSans 448 90 0 0 wbs_adr_i[2]
port 564 nsew signal input
flabel metal2 s 118762 -960 118874 480 0 FreeSans 448 90 0 0 wbs_adr_i[30]
port 565 nsew signal input
flabel metal2 s 122258 -960 122370 480 0 FreeSans 448 90 0 0 wbs_adr_i[31]
port 566 nsew signal input
flabel metal2 s 21794 -960 21906 480 0 FreeSans 448 90 0 0 wbs_adr_i[3]
port 567 nsew signal input
flabel metal2 s 26486 -960 26598 480 0 FreeSans 448 90 0 0 wbs_adr_i[4]
port 568 nsew signal input
flabel metal2 s 30074 -960 30186 480 0 FreeSans 448 90 0 0 wbs_adr_i[5]
port 569 nsew signal input
flabel metal2 s 33570 -960 33682 480 0 FreeSans 448 90 0 0 wbs_adr_i[6]
port 570 nsew signal input
flabel metal2 s 37158 -960 37270 480 0 FreeSans 448 90 0 0 wbs_adr_i[7]
port 571 nsew signal input
flabel metal2 s 40654 -960 40766 480 0 FreeSans 448 90 0 0 wbs_adr_i[8]
port 572 nsew signal input
flabel metal2 s 44242 -960 44354 480 0 FreeSans 448 90 0 0 wbs_adr_i[9]
port 573 nsew signal input
flabel metal2 s 4038 -960 4150 480 0 FreeSans 448 90 0 0 wbs_cyc_i
port 574 nsew signal input
flabel metal2 s 8730 -960 8842 480 0 FreeSans 448 90 0 0 wbs_dat_i[0]
port 575 nsew signal input
flabel metal2 s 48934 -960 49046 480 0 FreeSans 448 90 0 0 wbs_dat_i[10]
port 576 nsew signal input
flabel metal2 s 52522 -960 52634 480 0 FreeSans 448 90 0 0 wbs_dat_i[11]
port 577 nsew signal input
flabel metal2 s 56018 -960 56130 480 0 FreeSans 448 90 0 0 wbs_dat_i[12]
port 578 nsew signal input
flabel metal2 s 59606 -960 59718 480 0 FreeSans 448 90 0 0 wbs_dat_i[13]
port 579 nsew signal input
flabel metal2 s 63194 -960 63306 480 0 FreeSans 448 90 0 0 wbs_dat_i[14]
port 580 nsew signal input
flabel metal2 s 66690 -960 66802 480 0 FreeSans 448 90 0 0 wbs_dat_i[15]
port 581 nsew signal input
flabel metal2 s 70278 -960 70390 480 0 FreeSans 448 90 0 0 wbs_dat_i[16]
port 582 nsew signal input
flabel metal2 s 73774 -960 73886 480 0 FreeSans 448 90 0 0 wbs_dat_i[17]
port 583 nsew signal input
flabel metal2 s 77362 -960 77474 480 0 FreeSans 448 90 0 0 wbs_dat_i[18]
port 584 nsew signal input
flabel metal2 s 80858 -960 80970 480 0 FreeSans 448 90 0 0 wbs_dat_i[19]
port 585 nsew signal input
flabel metal2 s 13514 -960 13626 480 0 FreeSans 448 90 0 0 wbs_dat_i[1]
port 586 nsew signal input
flabel metal2 s 84446 -960 84558 480 0 FreeSans 448 90 0 0 wbs_dat_i[20]
port 587 nsew signal input
flabel metal2 s 87942 -960 88054 480 0 FreeSans 448 90 0 0 wbs_dat_i[21]
port 588 nsew signal input
flabel metal2 s 91530 -960 91642 480 0 FreeSans 448 90 0 0 wbs_dat_i[22]
port 589 nsew signal input
flabel metal2 s 95118 -960 95230 480 0 FreeSans 448 90 0 0 wbs_dat_i[23]
port 590 nsew signal input
flabel metal2 s 98614 -960 98726 480 0 FreeSans 448 90 0 0 wbs_dat_i[24]
port 591 nsew signal input
flabel metal2 s 102202 -960 102314 480 0 FreeSans 448 90 0 0 wbs_dat_i[25]
port 592 nsew signal input
flabel metal2 s 105698 -960 105810 480 0 FreeSans 448 90 0 0 wbs_dat_i[26]
port 593 nsew signal input
flabel metal2 s 109286 -960 109398 480 0 FreeSans 448 90 0 0 wbs_dat_i[27]
port 594 nsew signal input
flabel metal2 s 112782 -960 112894 480 0 FreeSans 448 90 0 0 wbs_dat_i[28]
port 595 nsew signal input
flabel metal2 s 116370 -960 116482 480 0 FreeSans 448 90 0 0 wbs_dat_i[29]
port 596 nsew signal input
flabel metal2 s 18206 -960 18318 480 0 FreeSans 448 90 0 0 wbs_dat_i[2]
port 597 nsew signal input
flabel metal2 s 119866 -960 119978 480 0 FreeSans 448 90 0 0 wbs_dat_i[30]
port 598 nsew signal input
flabel metal2 s 123454 -960 123566 480 0 FreeSans 448 90 0 0 wbs_dat_i[31]
port 599 nsew signal input
flabel metal2 s 22990 -960 23102 480 0 FreeSans 448 90 0 0 wbs_dat_i[3]
port 600 nsew signal input
flabel metal2 s 27682 -960 27794 480 0 FreeSans 448 90 0 0 wbs_dat_i[4]
port 601 nsew signal input
flabel metal2 s 31270 -960 31382 480 0 FreeSans 448 90 0 0 wbs_dat_i[5]
port 602 nsew signal input
flabel metal2 s 34766 -960 34878 480 0 FreeSans 448 90 0 0 wbs_dat_i[6]
port 603 nsew signal input
flabel metal2 s 38354 -960 38466 480 0 FreeSans 448 90 0 0 wbs_dat_i[7]
port 604 nsew signal input
flabel metal2 s 41850 -960 41962 480 0 FreeSans 448 90 0 0 wbs_dat_i[8]
port 605 nsew signal input
flabel metal2 s 45438 -960 45550 480 0 FreeSans 448 90 0 0 wbs_dat_i[9]
port 606 nsew signal input
flabel metal2 s 9926 -960 10038 480 0 FreeSans 448 90 0 0 wbs_dat_o[0]
port 607 nsew signal tristate
flabel metal2 s 50130 -960 50242 480 0 FreeSans 448 90 0 0 wbs_dat_o[10]
port 608 nsew signal tristate
flabel metal2 s 53718 -960 53830 480 0 FreeSans 448 90 0 0 wbs_dat_o[11]
port 609 nsew signal tristate
flabel metal2 s 57214 -960 57326 480 0 FreeSans 448 90 0 0 wbs_dat_o[12]
port 610 nsew signal tristate
flabel metal2 s 60802 -960 60914 480 0 FreeSans 448 90 0 0 wbs_dat_o[13]
port 611 nsew signal tristate
flabel metal2 s 64298 -960 64410 480 0 FreeSans 448 90 0 0 wbs_dat_o[14]
port 612 nsew signal tristate
flabel metal2 s 67886 -960 67998 480 0 FreeSans 448 90 0 0 wbs_dat_o[15]
port 613 nsew signal tristate
flabel metal2 s 71474 -960 71586 480 0 FreeSans 448 90 0 0 wbs_dat_o[16]
port 614 nsew signal tristate
flabel metal2 s 74970 -960 75082 480 0 FreeSans 448 90 0 0 wbs_dat_o[17]
port 615 nsew signal tristate
flabel metal2 s 78558 -960 78670 480 0 FreeSans 448 90 0 0 wbs_dat_o[18]
port 616 nsew signal tristate
flabel metal2 s 82054 -960 82166 480 0 FreeSans 448 90 0 0 wbs_dat_o[19]
port 617 nsew signal tristate
flabel metal2 s 14710 -960 14822 480 0 FreeSans 448 90 0 0 wbs_dat_o[1]
port 618 nsew signal tristate
flabel metal2 s 85642 -960 85754 480 0 FreeSans 448 90 0 0 wbs_dat_o[20]
port 619 nsew signal tristate
flabel metal2 s 89138 -960 89250 480 0 FreeSans 448 90 0 0 wbs_dat_o[21]
port 620 nsew signal tristate
flabel metal2 s 92726 -960 92838 480 0 FreeSans 448 90 0 0 wbs_dat_o[22]
port 621 nsew signal tristate
flabel metal2 s 96222 -960 96334 480 0 FreeSans 448 90 0 0 wbs_dat_o[23]
port 622 nsew signal tristate
flabel metal2 s 99810 -960 99922 480 0 FreeSans 448 90 0 0 wbs_dat_o[24]
port 623 nsew signal tristate
flabel metal2 s 103306 -960 103418 480 0 FreeSans 448 90 0 0 wbs_dat_o[25]
port 624 nsew signal tristate
flabel metal2 s 106894 -960 107006 480 0 FreeSans 448 90 0 0 wbs_dat_o[26]
port 625 nsew signal tristate
flabel metal2 s 110482 -960 110594 480 0 FreeSans 448 90 0 0 wbs_dat_o[27]
port 626 nsew signal tristate
flabel metal2 s 113978 -960 114090 480 0 FreeSans 448 90 0 0 wbs_dat_o[28]
port 627 nsew signal tristate
flabel metal2 s 117566 -960 117678 480 0 FreeSans 448 90 0 0 wbs_dat_o[29]
port 628 nsew signal tristate
flabel metal2 s 19402 -960 19514 480 0 FreeSans 448 90 0 0 wbs_dat_o[2]
port 629 nsew signal tristate
flabel metal2 s 121062 -960 121174 480 0 FreeSans 448 90 0 0 wbs_dat_o[30]
port 630 nsew signal tristate
flabel metal2 s 124650 -960 124762 480 0 FreeSans 448 90 0 0 wbs_dat_o[31]
port 631 nsew signal tristate
flabel metal2 s 24186 -960 24298 480 0 FreeSans 448 90 0 0 wbs_dat_o[3]
port 632 nsew signal tristate
flabel metal2 s 28878 -960 28990 480 0 FreeSans 448 90 0 0 wbs_dat_o[4]
port 633 nsew signal tristate
flabel metal2 s 32374 -960 32486 480 0 FreeSans 448 90 0 0 wbs_dat_o[5]
port 634 nsew signal tristate
flabel metal2 s 35962 -960 36074 480 0 FreeSans 448 90 0 0 wbs_dat_o[6]
port 635 nsew signal tristate
flabel metal2 s 39550 -960 39662 480 0 FreeSans 448 90 0 0 wbs_dat_o[7]
port 636 nsew signal tristate
flabel metal2 s 43046 -960 43158 480 0 FreeSans 448 90 0 0 wbs_dat_o[8]
port 637 nsew signal tristate
flabel metal2 s 46634 -960 46746 480 0 FreeSans 448 90 0 0 wbs_dat_o[9]
port 638 nsew signal tristate
flabel metal2 s 11122 -960 11234 480 0 FreeSans 448 90 0 0 wbs_sel_i[0]
port 639 nsew signal input
flabel metal2 s 15906 -960 16018 480 0 FreeSans 448 90 0 0 wbs_sel_i[1]
port 640 nsew signal input
flabel metal2 s 20598 -960 20710 480 0 FreeSans 448 90 0 0 wbs_sel_i[2]
port 641 nsew signal input
flabel metal2 s 25290 -960 25402 480 0 FreeSans 448 90 0 0 wbs_sel_i[3]
port 642 nsew signal input
flabel metal2 s 5234 -960 5346 480 0 FreeSans 448 90 0 0 wbs_stb_i
port 643 nsew signal input
flabel metal2 s 6430 -960 6542 480 0 FreeSans 448 90 0 0 wbs_we_i
port 644 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
